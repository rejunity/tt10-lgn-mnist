// Generated from: test_rnd_d16r1_8x1024_256i_1024o.npz
module net (
    input wire  [255:0] in,
    output wire [1023:0] out
);
    wire [1024:0] layer_0;
    wire [1024:0] layer_1;
    wire [1024:0] layer_2;
    wire [1024:0] layer_3;
    wire [1024:0] layer_4;
    wire [1024:0] layer_5;
    wire [1024:0] layer_6;

    // Layer 0 ============================================================
    assign layer_0[0] = in[6] | in[12]; 
    assign layer_0[1] = ~in[11] | (in[11] & in[1]); 
    assign layer_0[2] = ~in[0]; 
    assign layer_0[3] = ~(in[6] | in[11]); 
    assign layer_0[4] = in[1] | in[4]; 
    assign layer_0[5] = ~(in[4] ^ in[7]); 
    assign layer_0[6] = in[3] | in[13]; 
    assign layer_0[7] = ~in[4]; 
    assign layer_0[8] = in[9] & ~in[12]; 
    assign layer_0[9] = in[10] & ~in[5]; 
    assign layer_0[10] = in[13] & ~in[0]; 
    assign layer_0[11] = ~(in[14] | in[3]); 
    assign layer_0[12] = ~(in[11] ^ in[1]); 
    assign layer_0[13] = in[17] ^ in[9]; 
    assign layer_0[14] = in[11] ^ in[6]; 
    assign layer_0[15] = ~in[6]; 
    assign layer_0[16] = in[5] | in[17]; 
    assign layer_0[17] = ~(in[8] | in[5]); 
    assign layer_0[18] = in[17] & in[1]; 
    assign layer_0[19] = ~in[1] | (in[11] & in[1]); 
    assign layer_0[20] = ~in[5] | (in[5] & in[4]); 
    assign layer_0[21] = in[3] ^ in[4]; 
    assign layer_0[22] = in[6] ^ in[3]; 
    assign layer_0[23] = in[1] & ~in[6]; 
    assign layer_0[24] = in[3] & ~in[6]; 
    assign layer_0[25] = ~(in[7] ^ in[9]); 
    assign layer_0[26] = ~(in[2] | in[6]); 
    assign layer_0[27] = ~in[10] | (in[6] & in[10]); 
    assign layer_0[28] = in[3] & in[7]; 
    assign layer_0[29] = ~in[1]; 
    assign layer_0[30] = in[8] | in[1]; 
    assign layer_0[31] = in[15]; 
    assign layer_0[32] = ~(in[0] & in[4]); 
    assign layer_0[33] = in[6] & in[11]; 
    assign layer_0[34] = 1'b1; 
    assign layer_0[35] = ~in[19] | (in[17] & in[19]); 
    assign layer_0[36] = in[23]; 
    assign layer_0[37] = ~(in[3] ^ in[7]); 
    assign layer_0[38] = in[14]; 
    assign layer_0[39] = in[5] & ~in[15]; 
    assign layer_0[40] = ~(in[0] | in[1]); 
    assign layer_0[41] = ~(in[23] | in[21]); 
    assign layer_0[42] = ~in[14] | (in[14] & in[19]); 
    assign layer_0[43] = in[9] | in[14]; 
    assign layer_0[44] = ~in[7]; 
    assign layer_0[45] = ~in[3] | (in[4] & in[3]); 
    assign layer_0[46] = ~(in[5] ^ in[5]); 
    assign layer_0[47] = in[27] & ~in[24]; 
    assign layer_0[48] = 1'b1; 
    assign layer_0[49] = in[14] & in[22]; 
    assign layer_0[50] = ~in[16]; 
    assign layer_0[51] = in[17] ^ in[1]; 
    assign layer_0[52] = in[6] & ~in[11]; 
    assign layer_0[53] = in[25] & ~in[15]; 
    assign layer_0[54] = in[13] & ~in[29]; 
    assign layer_0[55] = in[27]; 
    assign layer_0[56] = ~(in[6] & in[9]); 
    assign layer_0[57] = in[7] | in[7]; 
    assign layer_0[58] = in[26] & ~in[4]; 
    assign layer_0[59] = in[18] & ~in[15]; 
    assign layer_0[60] = ~in[10]; 
    assign layer_0[61] = in[4]; 
    assign layer_0[62] = ~(in[18] ^ in[13]); 
    assign layer_0[63] = in[28] & ~in[1]; 
    assign layer_0[64] = ~in[0]; 
    assign layer_0[65] = in[25] & ~in[10]; 
    assign layer_0[66] = ~in[17] | (in[15] & in[17]); 
    assign layer_0[67] = ~(in[13] | in[31]); 
    assign layer_0[68] = ~(in[18] & in[16]); 
    assign layer_0[69] = in[13] ^ in[10]; 
    assign layer_0[70] = in[17]; 
    assign layer_0[71] = ~(in[5] | in[14]); 
    assign layer_0[72] = ~in[33] | (in[33] & in[19]); 
    assign layer_0[73] = ~(in[3] | in[1]); 
    assign layer_0[74] = 1'b1; 
    assign layer_0[75] = in[30] | in[19]; 
    assign layer_0[76] = in[5] & ~in[26]; 
    assign layer_0[77] = in[7]; 
    assign layer_0[78] = in[13] & ~in[34]; 
    assign layer_0[79] = ~in[21] | (in[21] & in[5]); 
    assign layer_0[80] = ~(in[16] ^ in[34]); 
    assign layer_0[81] = in[32] & in[33]; 
    assign layer_0[82] = ~in[4]; 
    assign layer_0[83] = ~in[12] | (in[12] & in[9]); 
    assign layer_0[84] = in[28] & ~in[23]; 
    assign layer_0[85] = ~in[13]; 
    assign layer_0[86] = 1'b0; 
    assign layer_0[87] = ~in[29] | (in[29] & in[23]); 
    assign layer_0[88] = in[21]; 
    assign layer_0[89] = ~(in[22] | in[37]); 
    assign layer_0[90] = in[33] & ~in[20]; 
    assign layer_0[91] = in[22] & in[25]; 
    assign layer_0[92] = ~in[7] | (in[7] & in[7]); 
    assign layer_0[93] = 1'b0; 
    assign layer_0[94] = in[13] & in[29]; 
    assign layer_0[95] = ~(in[20] ^ in[31]); 
    assign layer_0[96] = in[16] & ~in[25]; 
    assign layer_0[97] = 1'b1; 
    assign layer_0[98] = ~in[35] | (in[35] & in[25]); 
    assign layer_0[99] = in[33] & ~in[30]; 
    assign layer_0[100] = 1'b0; 
    assign layer_0[101] = 1'b0; 
    assign layer_0[102] = ~in[17] | (in[14] & in[17]); 
    assign layer_0[103] = ~in[35]; 
    assign layer_0[104] = in[15] | in[14]; 
    assign layer_0[105] = ~in[26] | (in[26] & in[19]); 
    assign layer_0[106] = in[28] & ~in[25]; 
    assign layer_0[107] = in[33] ^ in[36]; 
    assign layer_0[108] = in[38]; 
    assign layer_0[109] = in[28] ^ in[10]; 
    assign layer_0[110] = ~in[28]; 
    assign layer_0[111] = in[12]; 
    assign layer_0[112] = 1'b0; 
    assign layer_0[113] = 1'b0; 
    assign layer_0[114] = in[35] & ~in[35]; 
    assign layer_0[115] = in[21] & ~in[37]; 
    assign layer_0[116] = in[20]; 
    assign layer_0[117] = ~(in[24] ^ in[13]); 
    assign layer_0[118] = ~(in[29] ^ in[18]); 
    assign layer_0[119] = 1'b0; 
    assign layer_0[120] = in[17] & ~in[45]; 
    assign layer_0[121] = ~in[44] | (in[44] & in[16]); 
    assign layer_0[122] = in[46] & ~in[21]; 
    assign layer_0[123] = in[31] | in[26]; 
    assign layer_0[124] = in[27]; 
    assign layer_0[125] = in[41] ^ in[41]; 
    assign layer_0[126] = ~in[37]; 
    assign layer_0[127] = ~in[28] | (in[28] & in[24]); 
    assign layer_0[128] = ~in[30]; 
    assign layer_0[129] = ~in[29]; 
    assign layer_0[130] = in[40]; 
    assign layer_0[131] = ~in[29] | (in[29] & in[31]); 
    assign layer_0[132] = ~in[43]; 
    assign layer_0[133] = 1'b0; 
    assign layer_0[134] = ~in[27] | (in[36] & in[27]); 
    assign layer_0[135] = ~in[26] | (in[20] & in[26]); 
    assign layer_0[136] = in[44]; 
    assign layer_0[137] = ~(in[33] ^ in[17]); 
    assign layer_0[138] = ~in[43]; 
    assign layer_0[139] = ~in[22] | (in[22] & in[25]); 
    assign layer_0[140] = 1'b1; 
    assign layer_0[141] = 1'b0; 
    assign layer_0[142] = ~in[33]; 
    assign layer_0[143] = in[37] | in[44]; 
    assign layer_0[144] = in[20]; 
    assign layer_0[145] = ~in[26] | (in[20] & in[26]); 
    assign layer_0[146] = in[34] & in[31]; 
    assign layer_0[147] = in[51] ^ in[29]; 
    assign layer_0[148] = in[36] & in[45]; 
    assign layer_0[149] = ~(in[34] | in[20]); 
    assign layer_0[150] = in[21]; 
    assign layer_0[151] = ~in[53]; 
    assign layer_0[152] = ~in[23] | (in[23] & in[51]); 
    assign layer_0[153] = ~in[31]; 
    assign layer_0[154] = ~(in[44] ^ in[42]); 
    assign layer_0[155] = in[37] & ~in[39]; 
    assign layer_0[156] = in[41] | in[28]; 
    assign layer_0[157] = in[32] & in[50]; 
    assign layer_0[158] = in[34] ^ in[27]; 
    assign layer_0[159] = in[28] | in[28]; 
    assign layer_0[160] = 1'b1; 
    assign layer_0[161] = ~in[48]; 
    assign layer_0[162] = ~in[34]; 
    assign layer_0[163] = in[44] | in[27]; 
    assign layer_0[164] = in[26] ^ in[39]; 
    assign layer_0[165] = in[32]; 
    assign layer_0[166] = ~in[30] | (in[48] & in[30]); 
    assign layer_0[167] = ~in[33] | (in[53] & in[33]); 
    assign layer_0[168] = in[25]; 
    assign layer_0[169] = ~in[47]; 
    assign layer_0[170] = 1'b1; 
    assign layer_0[171] = ~(in[50] & in[55]); 
    assign layer_0[172] = ~(in[30] & in[29]); 
    assign layer_0[173] = ~(in[40] ^ in[57]); 
    assign layer_0[174] = in[50] & ~in[45]; 
    assign layer_0[175] = in[40] & in[48]; 
    assign layer_0[176] = 1'b0; 
    assign layer_0[177] = in[41] | in[47]; 
    assign layer_0[178] = in[36] | in[55]; 
    assign layer_0[179] = in[57] & ~in[29]; 
    assign layer_0[180] = in[52] & ~in[59]; 
    assign layer_0[181] = in[56] & ~in[54]; 
    assign layer_0[182] = ~(in[45] ^ in[42]); 
    assign layer_0[183] = in[45] ^ in[54]; 
    assign layer_0[184] = in[58] & in[52]; 
    assign layer_0[185] = in[49] ^ in[55]; 
    assign layer_0[186] = 1'b1; 
    assign layer_0[187] = ~in[57] | (in[57] & in[46]); 
    assign layer_0[188] = in[44] & ~in[45]; 
    assign layer_0[189] = ~in[42]; 
    assign layer_0[190] = ~(in[35] & in[56]); 
    assign layer_0[191] = ~in[39]; 
    assign layer_0[192] = in[61] | in[35]; 
    assign layer_0[193] = ~(in[53] ^ in[34]); 
    assign layer_0[194] = in[46]; 
    assign layer_0[195] = ~in[53]; 
    assign layer_0[196] = ~in[44]; 
    assign layer_0[197] = 1'b0; 
    assign layer_0[198] = in[38]; 
    assign layer_0[199] = in[64] & in[33]; 
    assign layer_0[200] = in[43] & ~in[41]; 
    assign layer_0[201] = ~in[47] | (in[47] & in[54]); 
    assign layer_0[202] = ~in[58] | (in[59] & in[58]); 
    assign layer_0[203] = in[41]; 
    assign layer_0[204] = in[37] & ~in[47]; 
    assign layer_0[205] = in[54] & in[54]; 
    assign layer_0[206] = ~in[46]; 
    assign layer_0[207] = ~(in[60] & in[58]); 
    assign layer_0[208] = in[41]; 
    assign layer_0[209] = ~in[39] | (in[54] & in[39]); 
    assign layer_0[210] = in[42] & in[63]; 
    assign layer_0[211] = ~(in[36] & in[37]); 
    assign layer_0[212] = in[52] & in[68]; 
    assign layer_0[213] = in[57]; 
    assign layer_0[214] = in[48] | in[53]; 
    assign layer_0[215] = in[65] & ~in[58]; 
    assign layer_0[216] = in[47] | in[40]; 
    assign layer_0[217] = in[60] | in[46]; 
    assign layer_0[218] = ~in[56] | (in[48] & in[56]); 
    assign layer_0[219] = ~in[40]; 
    assign layer_0[220] = in[46] ^ in[55]; 
    assign layer_0[221] = ~in[43]; 
    assign layer_0[222] = in[45] ^ in[44]; 
    assign layer_0[223] = ~in[52]; 
    assign layer_0[224] = ~(in[61] ^ in[56]); 
    assign layer_0[225] = ~in[63]; 
    assign layer_0[226] = ~(in[57] & in[59]); 
    assign layer_0[227] = in[45] & ~in[56]; 
    assign layer_0[228] = in[51] ^ in[57]; 
    assign layer_0[229] = in[44] & ~in[64]; 
    assign layer_0[230] = ~in[68]; 
    assign layer_0[231] = in[48] & ~in[41]; 
    assign layer_0[232] = 1'b1; 
    assign layer_0[233] = in[52] & ~in[44]; 
    assign layer_0[234] = in[53] ^ in[54]; 
    assign layer_0[235] = in[60] & in[72]; 
    assign layer_0[236] = ~(in[46] | in[61]); 
    assign layer_0[237] = ~in[70] | (in[70] & in[44]); 
    assign layer_0[238] = ~(in[61] & in[62]); 
    assign layer_0[239] = 1'b0; 
    assign layer_0[240] = ~in[57]; 
    assign layer_0[241] = ~(in[70] | in[53]); 
    assign layer_0[242] = 1'b0; 
    assign layer_0[243] = ~(in[63] | in[72]); 
    assign layer_0[244] = ~in[57] | (in[57] & in[59]); 
    assign layer_0[245] = in[72]; 
    assign layer_0[246] = ~in[46]; 
    assign layer_0[247] = ~in[50] | (in[50] & in[68]); 
    assign layer_0[248] = ~in[68] | (in[75] & in[68]); 
    assign layer_0[249] = in[54] ^ in[60]; 
    assign layer_0[250] = in[50] & ~in[64]; 
    assign layer_0[251] = in[70] & in[72]; 
    assign layer_0[252] = ~in[63] | (in[63] & in[74]); 
    assign layer_0[253] = in[76]; 
    assign layer_0[254] = in[57]; 
    assign layer_0[255] = in[48]; 
    assign layer_0[256] = ~(in[57] ^ in[73]); 
    assign layer_0[257] = in[56] & ~in[65]; 
    assign layer_0[258] = in[50] | in[50]; 
    assign layer_0[259] = ~in[72]; 
    assign layer_0[260] = 1'b1; 
    assign layer_0[261] = ~in[50]; 
    assign layer_0[262] = in[64] ^ in[54]; 
    assign layer_0[263] = in[77]; 
    assign layer_0[264] = 1'b1; 
    assign layer_0[265] = in[60] ^ in[56]; 
    assign layer_0[266] = in[56] & in[57]; 
    assign layer_0[267] = ~(in[55] & in[77]); 
    assign layer_0[268] = in[61] ^ in[76]; 
    assign layer_0[269] = ~(in[70] & in[64]); 
    assign layer_0[270] = in[78] & in[74]; 
    assign layer_0[271] = ~in[74] | (in[57] & in[74]); 
    assign layer_0[272] = in[62]; 
    assign layer_0[273] = 1'b1; 
    assign layer_0[274] = in[60] & ~in[79]; 
    assign layer_0[275] = ~in[66]; 
    assign layer_0[276] = 1'b0; 
    assign layer_0[277] = ~(in[70] & in[57]); 
    assign layer_0[278] = in[69] & in[60]; 
    assign layer_0[279] = in[64] & ~in[70]; 
    assign layer_0[280] = 1'b0; 
    assign layer_0[281] = in[80] & ~in[75]; 
    assign layer_0[282] = ~in[77] | (in[77] & in[70]); 
    assign layer_0[283] = ~(in[64] ^ in[68]); 
    assign layer_0[284] = in[84]; 
    assign layer_0[285] = in[79] & in[84]; 
    assign layer_0[286] = in[73] & in[59]; 
    assign layer_0[287] = 1'b1; 
    assign layer_0[288] = in[73] | in[57]; 
    assign layer_0[289] = 1'b1; 
    assign layer_0[290] = in[74]; 
    assign layer_0[291] = in[69] & ~in[75]; 
    assign layer_0[292] = in[62] & ~in[68]; 
    assign layer_0[293] = in[87] | in[64]; 
    assign layer_0[294] = in[84] ^ in[63]; 
    assign layer_0[295] = 1'b1; 
    assign layer_0[296] = ~(in[64] ^ in[61]); 
    assign layer_0[297] = ~(in[86] & in[83]); 
    assign layer_0[298] = 1'b0; 
    assign layer_0[299] = ~in[67]; 
    assign layer_0[300] = 1'b1; 
    assign layer_0[301] = ~(in[60] & in[73]); 
    assign layer_0[302] = in[69]; 
    assign layer_0[303] = ~in[88]; 
    assign layer_0[304] = ~in[90] | (in[82] & in[90]); 
    assign layer_0[305] = ~in[79] | (in[76] & in[79]); 
    assign layer_0[306] = in[74]; 
    assign layer_0[307] = ~(in[72] ^ in[85]); 
    assign layer_0[308] = in[92] & ~in[77]; 
    assign layer_0[309] = in[76] & ~in[85]; 
    assign layer_0[310] = in[80] & in[93]; 
    assign layer_0[311] = ~in[86] | (in[68] & in[86]); 
    assign layer_0[312] = ~(in[75] | in[78]); 
    assign layer_0[313] = ~in[92]; 
    assign layer_0[314] = ~in[88]; 
    assign layer_0[315] = ~in[94]; 
    assign layer_0[316] = in[81]; 
    assign layer_0[317] = 1'b0; 
    assign layer_0[318] = 1'b0; 
    assign layer_0[319] = ~in[95]; 
    assign layer_0[320] = ~(in[91] ^ in[81]); 
    assign layer_0[321] = in[81] ^ in[86]; 
    assign layer_0[322] = ~in[84]; 
    assign layer_0[323] = in[95] & ~in[66]; 
    assign layer_0[324] = ~in[85] | (in[85] & in[65]); 
    assign layer_0[325] = in[67] | in[68]; 
    assign layer_0[326] = ~in[84] | (in[84] & in[74]); 
    assign layer_0[327] = in[90] & ~in[65]; 
    assign layer_0[328] = in[96] | in[77]; 
    assign layer_0[329] = ~(in[78] ^ in[65]); 
    assign layer_0[330] = in[69]; 
    assign layer_0[331] = in[78]; 
    assign layer_0[332] = in[79] | in[66]; 
    assign layer_0[333] = in[91] & in[85]; 
    assign layer_0[334] = ~in[90] | (in[90] & in[79]); 
    assign layer_0[335] = in[72] | in[94]; 
    assign layer_0[336] = ~(in[81] ^ in[90]); 
    assign layer_0[337] = in[92] | in[77]; 
    assign layer_0[338] = in[96]; 
    assign layer_0[339] = ~(in[95] ^ in[88]); 
    assign layer_0[340] = ~in[100] | (in[97] & in[100]); 
    assign layer_0[341] = in[97] & ~in[68]; 
    assign layer_0[342] = ~(in[87] ^ in[96]); 
    assign layer_0[343] = in[101] | in[70]; 
    assign layer_0[344] = ~(in[84] | in[94]); 
    assign layer_0[345] = in[78]; 
    assign layer_0[346] = ~in[77]; 
    assign layer_0[347] = ~(in[92] | in[83]); 
    assign layer_0[348] = ~in[79] | (in[79] & in[72]); 
    assign layer_0[349] = ~in[76] | (in[76] & in[79]); 
    assign layer_0[350] = ~in[89] | (in[73] & in[89]); 
    assign layer_0[351] = ~in[98] | (in[102] & in[98]); 
    assign layer_0[352] = ~in[103]; 
    assign layer_0[353] = ~in[78]; 
    assign layer_0[354] = in[100] & ~in[88]; 
    assign layer_0[355] = ~(in[73] & in[92]); 
    assign layer_0[356] = in[99] | in[79]; 
    assign layer_0[357] = in[102] & ~in[86]; 
    assign layer_0[358] = in[74] | in[89]; 
    assign layer_0[359] = in[78] ^ in[73]; 
    assign layer_0[360] = ~(in[102] & in[94]); 
    assign layer_0[361] = ~in[95] | (in[95] & in[93]); 
    assign layer_0[362] = ~(in[91] | in[86]); 
    assign layer_0[363] = ~in[99]; 
    assign layer_0[364] = in[78] & ~in[78]; 
    assign layer_0[365] = ~in[106]; 
    assign layer_0[366] = 1'b0; 
    assign layer_0[367] = in[79]; 
    assign layer_0[368] = ~in[99]; 
    assign layer_0[369] = 1'b0; 
    assign layer_0[370] = ~in[83] | (in[102] & in[83]); 
    assign layer_0[371] = 1'b0; 
    assign layer_0[372] = ~(in[79] ^ in[84]); 
    assign layer_0[373] = in[101]; 
    assign layer_0[374] = ~in[90]; 
    assign layer_0[375] = in[81] ^ in[77]; 
    assign layer_0[376] = 1'b1; 
    assign layer_0[377] = ~in[89] | (in[89] & in[78]); 
    assign layer_0[378] = 1'b1; 
    assign layer_0[379] = in[91] | in[82]; 
    assign layer_0[380] = in[81] & in[81]; 
    assign layer_0[381] = in[87]; 
    assign layer_0[382] = in[99] & ~in[102]; 
    assign layer_0[383] = ~in[91]; 
    assign layer_0[384] = in[104] | in[104]; 
    assign layer_0[385] = in[84] | in[81]; 
    assign layer_0[386] = ~(in[97] ^ in[98]); 
    assign layer_0[387] = in[99] ^ in[108]; 
    assign layer_0[388] = in[93] & ~in[102]; 
    assign layer_0[389] = in[90]; 
    assign layer_0[390] = ~(in[108] | in[96]); 
    assign layer_0[391] = in[90]; 
    assign layer_0[392] = 1'b1; 
    assign layer_0[393] = ~(in[84] ^ in[87]); 
    assign layer_0[394] = ~in[83]; 
    assign layer_0[395] = in[93]; 
    assign layer_0[396] = ~(in[95] & in[86]); 
    assign layer_0[397] = 1'b0; 
    assign layer_0[398] = 1'b1; 
    assign layer_0[399] = in[83] & in[87]; 
    assign layer_0[400] = 1'b1; 
    assign layer_0[401] = in[114] ^ in[105]; 
    assign layer_0[402] = ~(in[90] ^ in[99]); 
    assign layer_0[403] = in[94]; 
    assign layer_0[404] = 1'b1; 
    assign layer_0[405] = ~(in[95] ^ in[107]); 
    assign layer_0[406] = in[112] & ~in[114]; 
    assign layer_0[407] = in[97] & ~in[103]; 
    assign layer_0[408] = in[111]; 
    assign layer_0[409] = in[108] & ~in[105]; 
    assign layer_0[410] = ~in[107] | (in[107] & in[88]); 
    assign layer_0[411] = ~in[89]; 
    assign layer_0[412] = ~in[112]; 
    assign layer_0[413] = in[112] & in[108]; 
    assign layer_0[414] = 1'b1; 
    assign layer_0[415] = ~(in[108] | in[88]); 
    assign layer_0[416] = in[112] & ~in[88]; 
    assign layer_0[417] = ~(in[90] | in[93]); 
    assign layer_0[418] = in[110]; 
    assign layer_0[419] = in[117]; 
    assign layer_0[420] = ~in[100]; 
    assign layer_0[421] = in[90]; 
    assign layer_0[422] = ~in[98] | (in[98] & in[120]); 
    assign layer_0[423] = ~in[93] | (in[111] & in[93]); 
    assign layer_0[424] = ~(in[91] ^ in[106]); 
    assign layer_0[425] = 1'b0; 
    assign layer_0[426] = in[94] & ~in[97]; 
    assign layer_0[427] = in[103]; 
    assign layer_0[428] = 1'b0; 
    assign layer_0[429] = ~in[105]; 
    assign layer_0[430] = ~(in[104] | in[102]); 
    assign layer_0[431] = ~(in[99] | in[118]); 
    assign layer_0[432] = 1'b0; 
    assign layer_0[433] = in[121] & ~in[113]; 
    assign layer_0[434] = in[92] & in[119]; 
    assign layer_0[435] = 1'b0; 
    assign layer_0[436] = in[106] | in[106]; 
    assign layer_0[437] = ~(in[100] | in[117]); 
    assign layer_0[438] = ~in[92]; 
    assign layer_0[439] = in[99] | in[104]; 
    assign layer_0[440] = ~in[110] | (in[110] & in[122]); 
    assign layer_0[441] = ~in[111]; 
    assign layer_0[442] = ~in[100]; 
    assign layer_0[443] = ~in[122]; 
    assign layer_0[444] = 1'b0; 
    assign layer_0[445] = 1'b0; 
    assign layer_0[446] = in[96] | in[94]; 
    assign layer_0[447] = in[105] & ~in[96]; 
    assign layer_0[448] = ~in[97]; 
    assign layer_0[449] = ~in[113] | (in[97] & in[113]); 
    assign layer_0[450] = in[122] & ~in[119]; 
    assign layer_0[451] = in[127]; 
    assign layer_0[452] = in[128] & ~in[121]; 
    assign layer_0[453] = ~in[122]; 
    assign layer_0[454] = ~in[116]; 
    assign layer_0[455] = ~(in[109] | in[122]); 
    assign layer_0[456] = ~in[107]; 
    assign layer_0[457] = in[127]; 
    assign layer_0[458] = ~(in[99] & in[124]); 
    assign layer_0[459] = ~in[124]; 
    assign layer_0[460] = ~(in[112] ^ in[119]); 
    assign layer_0[461] = in[130] & in[113]; 
    assign layer_0[462] = in[110] & ~in[110]; 
    assign layer_0[463] = ~in[108]; 
    assign layer_0[464] = in[105]; 
    assign layer_0[465] = 1'b1; 
    assign layer_0[466] = 1'b1; 
    assign layer_0[467] = ~in[102] | (in[102] & in[116]); 
    assign layer_0[468] = in[100]; 
    assign layer_0[469] = in[127] & ~in[108]; 
    assign layer_0[470] = in[104] & ~in[100]; 
    assign layer_0[471] = 1'b1; 
    assign layer_0[472] = ~in[115]; 
    assign layer_0[473] = in[105] | in[132]; 
    assign layer_0[474] = in[117] & in[104]; 
    assign layer_0[475] = in[116]; 
    assign layer_0[476] = ~in[132]; 
    assign layer_0[477] = ~(in[112] & in[127]); 
    assign layer_0[478] = in[122] & ~in[119]; 
    assign layer_0[479] = in[122]; 
    assign layer_0[480] = in[114] & in[117]; 
    assign layer_0[481] = ~in[103] | (in[103] & in[113]); 
    assign layer_0[482] = in[120] & ~in[133]; 
    assign layer_0[483] = in[119] & in[105]; 
    assign layer_0[484] = in[118] & ~in[113]; 
    assign layer_0[485] = ~(in[106] ^ in[127]); 
    assign layer_0[486] = 1'b0; 
    assign layer_0[487] = in[121] & in[120]; 
    assign layer_0[488] = ~(in[105] | in[111]); 
    assign layer_0[489] = 1'b1; 
    assign layer_0[490] = in[116] & ~in[137]; 
    assign layer_0[491] = 1'b0; 
    assign layer_0[492] = 1'b0; 
    assign layer_0[493] = in[112]; 
    assign layer_0[494] = 1'b0; 
    assign layer_0[495] = in[139] & in[118]; 
    assign layer_0[496] = ~(in[107] | in[137]); 
    assign layer_0[497] = ~in[110]; 
    assign layer_0[498] = in[140] ^ in[125]; 
    assign layer_0[499] = ~in[127]; 
    assign layer_0[500] = ~(in[123] | in[109]); 
    assign layer_0[501] = ~in[111]; 
    assign layer_0[502] = ~in[140] | (in[135] & in[140]); 
    assign layer_0[503] = in[136] & in[119]; 
    assign layer_0[504] = ~(in[119] ^ in[125]); 
    assign layer_0[505] = in[127] & ~in[130]; 
    assign layer_0[506] = in[124]; 
    assign layer_0[507] = ~in[138] | (in[137] & in[138]); 
    assign layer_0[508] = in[127] & ~in[137]; 
    assign layer_0[509] = in[131]; 
    assign layer_0[510] = ~in[125] | (in[126] & in[125]); 
    assign layer_0[511] = in[130] & ~in[129]; 
    assign layer_0[512] = 1'b1; 
    assign layer_0[513] = ~in[122]; 
    assign layer_0[514] = in[134] | in[142]; 
    assign layer_0[515] = in[118] ^ in[120]; 
    assign layer_0[516] = in[129]; 
    assign layer_0[517] = in[141] & ~in[127]; 
    assign layer_0[518] = in[138] | in[119]; 
    assign layer_0[519] = ~(in[120] ^ in[141]); 
    assign layer_0[520] = 1'b1; 
    assign layer_0[521] = ~in[145]; 
    assign layer_0[522] = in[115] & ~in[124]; 
    assign layer_0[523] = in[125] & in[125]; 
    assign layer_0[524] = in[128] & ~in[115]; 
    assign layer_0[525] = ~(in[122] | in[141]); 
    assign layer_0[526] = ~(in[124] ^ in[136]); 
    assign layer_0[527] = ~(in[147] & in[118]); 
    assign layer_0[528] = 1'b0; 
    assign layer_0[529] = ~(in[137] & in[126]); 
    assign layer_0[530] = in[122] | in[141]; 
    assign layer_0[531] = ~(in[137] ^ in[144]); 
    assign layer_0[532] = ~in[144] | (in[144] & in[140]); 
    assign layer_0[533] = ~(in[134] | in[133]); 
    assign layer_0[534] = in[128] & ~in[144]; 
    assign layer_0[535] = ~in[128]; 
    assign layer_0[536] = in[144]; 
    assign layer_0[537] = ~in[145] | (in[145] & in[141]); 
    assign layer_0[538] = in[145] & ~in[137]; 
    assign layer_0[539] = ~(in[124] | in[127]); 
    assign layer_0[540] = in[122] & ~in[127]; 
    assign layer_0[541] = ~in[142]; 
    assign layer_0[542] = in[125] & ~in[126]; 
    assign layer_0[543] = ~(in[142] & in[125]); 
    assign layer_0[544] = ~in[124] | (in[150] & in[124]); 
    assign layer_0[545] = ~in[129]; 
    assign layer_0[546] = ~in[141]; 
    assign layer_0[547] = in[134] & ~in[151]; 
    assign layer_0[548] = in[142] | in[138]; 
    assign layer_0[549] = in[126] | in[140]; 
    assign layer_0[550] = ~(in[147] & in[140]); 
    assign layer_0[551] = in[124] ^ in[141]; 
    assign layer_0[552] = ~in[140] | (in[140] & in[150]); 
    assign layer_0[553] = ~(in[126] & in[149]); 
    assign layer_0[554] = in[139] ^ in[146]; 
    assign layer_0[555] = in[142] & ~in[122]; 
    assign layer_0[556] = 1'b0; 
    assign layer_0[557] = 1'b1; 
    assign layer_0[558] = in[151] & ~in[149]; 
    assign layer_0[559] = ~in[150]; 
    assign layer_0[560] = in[137] | in[149]; 
    assign layer_0[561] = in[132] & in[144]; 
    assign layer_0[562] = in[148] ^ in[127]; 
    assign layer_0[563] = in[140]; 
    assign layer_0[564] = ~in[132]; 
    assign layer_0[565] = in[155] | in[127]; 
    assign layer_0[566] = in[129] & in[136]; 
    assign layer_0[567] = ~in[141]; 
    assign layer_0[568] = in[128] ^ in[154]; 
    assign layer_0[569] = in[149]; 
    assign layer_0[570] = in[136]; 
    assign layer_0[571] = in[146]; 
    assign layer_0[572] = ~in[130]; 
    assign layer_0[573] = in[138] & ~in[131]; 
    assign layer_0[574] = in[135] & ~in[151]; 
    assign layer_0[575] = ~(in[154] | in[155]); 
    assign layer_0[576] = in[130] & ~in[146]; 
    assign layer_0[577] = in[130] & ~in[156]; 
    assign layer_0[578] = ~(in[152] ^ in[128]); 
    assign layer_0[579] = in[158] ^ in[160]; 
    assign layer_0[580] = in[151] & ~in[158]; 
    assign layer_0[581] = in[150] | in[153]; 
    assign layer_0[582] = in[134] & ~in[145]; 
    assign layer_0[583] = in[144]; 
    assign layer_0[584] = in[146]; 
    assign layer_0[585] = in[135] ^ in[151]; 
    assign layer_0[586] = 1'b1; 
    assign layer_0[587] = ~in[146]; 
    assign layer_0[588] = in[134] & ~in[134]; 
    assign layer_0[589] = ~in[159]; 
    assign layer_0[590] = in[150] ^ in[130]; 
    assign layer_0[591] = 1'b1; 
    assign layer_0[592] = in[160] ^ in[146]; 
    assign layer_0[593] = ~in[152] | (in[131] & in[152]); 
    assign layer_0[594] = ~in[152] | (in[150] & in[152]); 
    assign layer_0[595] = ~in[138]; 
    assign layer_0[596] = ~(in[143] | in[151]); 
    assign layer_0[597] = ~in[163] | (in[155] & in[163]); 
    assign layer_0[598] = in[146]; 
    assign layer_0[599] = in[146]; 
    assign layer_0[600] = ~(in[134] & in[157]); 
    assign layer_0[601] = ~in[142]; 
    assign layer_0[602] = in[137] ^ in[151]; 
    assign layer_0[603] = in[162]; 
    assign layer_0[604] = ~in[149] | (in[149] & in[151]); 
    assign layer_0[605] = ~in[143]; 
    assign layer_0[606] = in[164]; 
    assign layer_0[607] = ~in[156]; 
    assign layer_0[608] = ~(in[163] | in[152]); 
    assign layer_0[609] = in[160]; 
    assign layer_0[610] = in[142] & ~in[157]; 
    assign layer_0[611] = 1'b0; 
    assign layer_0[612] = in[152] | in[167]; 
    assign layer_0[613] = ~(in[157] ^ in[155]); 
    assign layer_0[614] = ~in[162]; 
    assign layer_0[615] = ~in[143] | (in[143] & in[146]); 
    assign layer_0[616] = in[139]; 
    assign layer_0[617] = ~in[147]; 
    assign layer_0[618] = ~in[160]; 
    assign layer_0[619] = in[146] | in[154]; 
    assign layer_0[620] = in[158] ^ in[164]; 
    assign layer_0[621] = 1'b1; 
    assign layer_0[622] = 1'b0; 
    assign layer_0[623] = ~(in[162] | in[148]); 
    assign layer_0[624] = ~in[170]; 
    assign layer_0[625] = ~in[148]; 
    assign layer_0[626] = ~(in[161] & in[152]); 
    assign layer_0[627] = ~(in[155] & in[154]); 
    assign layer_0[628] = ~in[169] | (in[169] & in[160]); 
    assign layer_0[629] = in[147] ^ in[143]; 
    assign layer_0[630] = in[146] | in[165]; 
    assign layer_0[631] = ~in[144] | (in[144] & in[162]); 
    assign layer_0[632] = in[163] ^ in[144]; 
    assign layer_0[633] = in[156]; 
    assign layer_0[634] = ~(in[166] & in[154]); 
    assign layer_0[635] = 1'b1; 
    assign layer_0[636] = 1'b0; 
    assign layer_0[637] = in[152] & ~in[142]; 
    assign layer_0[638] = in[154] & ~in[165]; 
    assign layer_0[639] = in[164] & ~in[168]; 
    assign layer_0[640] = ~in[145]; 
    assign layer_0[641] = in[150] & in[164]; 
    assign layer_0[642] = in[147] & in[168]; 
    assign layer_0[643] = in[145] ^ in[164]; 
    assign layer_0[644] = in[158] & ~in[165]; 
    assign layer_0[645] = 1'b0; 
    assign layer_0[646] = in[154] & ~in[166]; 
    assign layer_0[647] = in[170] & in[161]; 
    assign layer_0[648] = in[158] | in[150]; 
    assign layer_0[649] = in[163] ^ in[157]; 
    assign layer_0[650] = in[151] & in[156]; 
    assign layer_0[651] = in[161] ^ in[148]; 
    assign layer_0[652] = in[155] & ~in[177]; 
    assign layer_0[653] = ~in[173]; 
    assign layer_0[654] = in[149]; 
    assign layer_0[655] = 1'b0; 
    assign layer_0[656] = ~in[170]; 
    assign layer_0[657] = in[167] & ~in[161]; 
    assign layer_0[658] = ~in[169]; 
    assign layer_0[659] = in[180] ^ in[167]; 
    assign layer_0[660] = ~in[159] | (in[159] & in[168]); 
    assign layer_0[661] = in[175] ^ in[166]; 
    assign layer_0[662] = ~(in[180] ^ in[151]); 
    assign layer_0[663] = in[159]; 
    assign layer_0[664] = ~in[151]; 
    assign layer_0[665] = ~(in[149] ^ in[162]); 
    assign layer_0[666] = in[150] | in[152]; 
    assign layer_0[667] = 1'b0; 
    assign layer_0[668] = ~(in[180] | in[153]); 
    assign layer_0[669] = ~(in[161] & in[170]); 
    assign layer_0[670] = ~in[175]; 
    assign layer_0[671] = ~in[167] | (in[176] & in[167]); 
    assign layer_0[672] = ~(in[181] ^ in[160]); 
    assign layer_0[673] = in[182]; 
    assign layer_0[674] = in[156] | in[175]; 
    assign layer_0[675] = in[156] | in[183]; 
    assign layer_0[676] = 1'b1; 
    assign layer_0[677] = in[156] & in[158]; 
    assign layer_0[678] = in[183]; 
    assign layer_0[679] = ~in[158] | (in[158] & in[175]); 
    assign layer_0[680] = ~in[164]; 
    assign layer_0[681] = in[185] & in[155]; 
    assign layer_0[682] = ~in[183]; 
    assign layer_0[683] = ~in[162] | (in[180] & in[162]); 
    assign layer_0[684] = ~(in[162] | in[174]); 
    assign layer_0[685] = ~(in[182] & in[161]); 
    assign layer_0[686] = 1'b1; 
    assign layer_0[687] = in[173]; 
    assign layer_0[688] = ~in[168]; 
    assign layer_0[689] = ~(in[175] & in[168]); 
    assign layer_0[690] = in[177] & ~in[165]; 
    assign layer_0[691] = in[183] & ~in[173]; 
    assign layer_0[692] = in[187] & in[160]; 
    assign layer_0[693] = in[182] ^ in[158]; 
    assign layer_0[694] = ~in[163] | (in[163] & in[179]); 
    assign layer_0[695] = ~in[165] | (in[165] & in[165]); 
    assign layer_0[696] = in[175]; 
    assign layer_0[697] = in[159] & ~in[165]; 
    assign layer_0[698] = ~in[163] | (in[158] & in[163]); 
    assign layer_0[699] = 1'b0; 
    assign layer_0[700] = 1'b0; 
    assign layer_0[701] = ~(in[172] | in[159]); 
    assign layer_0[702] = in[173] & in[175]; 
    assign layer_0[703] = in[183] & in[176]; 
    assign layer_0[704] = ~(in[183] ^ in[174]); 
    assign layer_0[705] = ~in[165]; 
    assign layer_0[706] = in[167] & ~in[191]; 
    assign layer_0[707] = 1'b1; 
    assign layer_0[708] = in[175] | in[163]; 
    assign layer_0[709] = in[167]; 
    assign layer_0[710] = 1'b1; 
    assign layer_0[711] = ~(in[167] | in[189]); 
    assign layer_0[712] = ~(in[185] | in[191]); 
    assign layer_0[713] = ~in[191]; 
    assign layer_0[714] = 1'b0; 
    assign layer_0[715] = ~(in[174] & in[172]); 
    assign layer_0[716] = ~in[191] | (in[191] & in[185]); 
    assign layer_0[717] = 1'b0; 
    assign layer_0[718] = in[168] & ~in[179]; 
    assign layer_0[719] = ~(in[176] | in[188]); 
    assign layer_0[720] = in[185] & in[176]; 
    assign layer_0[721] = in[187] ^ in[164]; 
    assign layer_0[722] = ~in[178] | (in[178] & in[168]); 
    assign layer_0[723] = in[169]; 
    assign layer_0[724] = in[169] ^ in[172]; 
    assign layer_0[725] = ~in[196]; 
    assign layer_0[726] = in[194] & ~in[174]; 
    assign layer_0[727] = 1'b1; 
    assign layer_0[728] = ~in[192] | (in[169] & in[192]); 
    assign layer_0[729] = in[181] | in[196]; 
    assign layer_0[730] = ~in[195] | (in[165] & in[195]); 
    assign layer_0[731] = in[181] ^ in[180]; 
    assign layer_0[732] = 1'b0; 
    assign layer_0[733] = ~in[167] | (in[194] & in[167]); 
    assign layer_0[734] = ~(in[169] & in[170]); 
    assign layer_0[735] = ~in[190] | (in[190] & in[197]); 
    assign layer_0[736] = in[167] ^ in[193]; 
    assign layer_0[737] = 1'b1; 
    assign layer_0[738] = ~in[195] | (in[183] & in[195]); 
    assign layer_0[739] = ~in[190] | (in[180] & in[190]); 
    assign layer_0[740] = ~(in[195] & in[173]); 
    assign layer_0[741] = in[195] | in[188]; 
    assign layer_0[742] = in[180]; 
    assign layer_0[743] = 1'b0; 
    assign layer_0[744] = ~in[169] | (in[193] & in[169]); 
    assign layer_0[745] = ~(in[181] ^ in[189]); 
    assign layer_0[746] = ~(in[188] ^ in[174]); 
    assign layer_0[747] = in[180] & ~in[199]; 
    assign layer_0[748] = in[187]; 
    assign layer_0[749] = in[179]; 
    assign layer_0[750] = ~(in[193] & in[180]); 
    assign layer_0[751] = ~in[200]; 
    assign layer_0[752] = in[193] & in[194]; 
    assign layer_0[753] = in[193] ^ in[197]; 
    assign layer_0[754] = ~in[178] | (in[178] & in[171]); 
    assign layer_0[755] = in[188] & ~in[176]; 
    assign layer_0[756] = ~(in[178] & in[203]); 
    assign layer_0[757] = in[190]; 
    assign layer_0[758] = in[193] ^ in[197]; 
    assign layer_0[759] = in[174] & ~in[177]; 
    assign layer_0[760] = ~(in[194] & in[201]); 
    assign layer_0[761] = ~(in[195] | in[188]); 
    assign layer_0[762] = 1'b1; 
    assign layer_0[763] = in[187] ^ in[179]; 
    assign layer_0[764] = in[176] & ~in[198]; 
    assign layer_0[765] = in[182] & in[196]; 
    assign layer_0[766] = ~(in[198] | in[192]); 
    assign layer_0[767] = in[181] | in[196]; 
    assign layer_0[768] = ~(in[192] & in[186]); 
    assign layer_0[769] = 1'b1; 
    assign layer_0[770] = ~(in[201] ^ in[182]); 
    assign layer_0[771] = ~(in[205] & in[200]); 
    assign layer_0[772] = ~in[194]; 
    assign layer_0[773] = ~(in[187] ^ in[196]); 
    assign layer_0[774] = in[180] | in[196]; 
    assign layer_0[775] = 1'b1; 
    assign layer_0[776] = ~(in[185] & in[188]); 
    assign layer_0[777] = in[203] & in[186]; 
    assign layer_0[778] = ~in[203]; 
    assign layer_0[779] = ~(in[180] & in[195]); 
    assign layer_0[780] = 1'b0; 
    assign layer_0[781] = 1'b1; 
    assign layer_0[782] = ~in[178]; 
    assign layer_0[783] = in[183] | in[199]; 
    assign layer_0[784] = in[206] & in[199]; 
    assign layer_0[785] = ~in[183]; 
    assign layer_0[786] = ~(in[197] | in[210]); 
    assign layer_0[787] = 1'b0; 
    assign layer_0[788] = in[209] & ~in[188]; 
    assign layer_0[789] = in[192] | in[199]; 
    assign layer_0[790] = ~(in[181] & in[196]); 
    assign layer_0[791] = ~(in[206] ^ in[193]); 
    assign layer_0[792] = ~in[207]; 
    assign layer_0[793] = 1'b0; 
    assign layer_0[794] = 1'b1; 
    assign layer_0[795] = ~(in[210] | in[212]); 
    assign layer_0[796] = ~in[208]; 
    assign layer_0[797] = ~in[194]; 
    assign layer_0[798] = in[211] ^ in[205]; 
    assign layer_0[799] = 1'b1; 
    assign layer_0[800] = in[183] ^ in[198]; 
    assign layer_0[801] = in[195] & ~in[184]; 
    assign layer_0[802] = in[188]; 
    assign layer_0[803] = ~in[206] | (in[206] & in[201]); 
    assign layer_0[804] = in[199]; 
    assign layer_0[805] = in[204] & ~in[184]; 
    assign layer_0[806] = in[200] & ~in[198]; 
    assign layer_0[807] = ~in[210]; 
    assign layer_0[808] = in[207]; 
    assign layer_0[809] = in[193] & ~in[195]; 
    assign layer_0[810] = in[200] | in[188]; 
    assign layer_0[811] = in[191] ^ in[188]; 
    assign layer_0[812] = ~(in[194] & in[200]); 
    assign layer_0[813] = in[198]; 
    assign layer_0[814] = ~(in[195] | in[216]); 
    assign layer_0[815] = in[206] & ~in[191]; 
    assign layer_0[816] = in[196]; 
    assign layer_0[817] = in[189] ^ in[188]; 
    assign layer_0[818] = in[208] & in[211]; 
    assign layer_0[819] = in[190] & in[202]; 
    assign layer_0[820] = ~in[201]; 
    assign layer_0[821] = in[216]; 
    assign layer_0[822] = ~in[209] | (in[209] & in[210]); 
    assign layer_0[823] = in[220] & ~in[188]; 
    assign layer_0[824] = ~in[204]; 
    assign layer_0[825] = ~in[199] | (in[199] & in[205]); 
    assign layer_0[826] = in[211]; 
    assign layer_0[827] = in[211] & ~in[197]; 
    assign layer_0[828] = ~in[219] | (in[219] & in[207]); 
    assign layer_0[829] = ~in[205]; 
    assign layer_0[830] = in[192] ^ in[191]; 
    assign layer_0[831] = ~(in[213] ^ in[217]); 
    assign layer_0[832] = in[194] ^ in[195]; 
    assign layer_0[833] = ~(in[206] & in[192]); 
    assign layer_0[834] = 1'b1; 
    assign layer_0[835] = ~in[214] | (in[214] & in[214]); 
    assign layer_0[836] = 1'b1; 
    assign layer_0[837] = 1'b1; 
    assign layer_0[838] = in[194]; 
    assign layer_0[839] = in[206] | in[200]; 
    assign layer_0[840] = ~in[212] | (in[212] & in[213]); 
    assign layer_0[841] = 1'b0; 
    assign layer_0[842] = in[212]; 
    assign layer_0[843] = ~in[218]; 
    assign layer_0[844] = ~(in[215] & in[206]); 
    assign layer_0[845] = ~(in[197] & in[204]); 
    assign layer_0[846] = 1'b0; 
    assign layer_0[847] = in[202]; 
    assign layer_0[848] = ~in[213] | (in[210] & in[213]); 
    assign layer_0[849] = ~in[217]; 
    assign layer_0[850] = in[220] & in[218]; 
    assign layer_0[851] = ~in[224] | (in[224] & in[212]); 
    assign layer_0[852] = in[199]; 
    assign layer_0[853] = ~(in[214] & in[223]); 
    assign layer_0[854] = ~in[203] | (in[202] & in[203]); 
    assign layer_0[855] = ~in[201] | (in[201] & in[198]); 
    assign layer_0[856] = 1'b0; 
    assign layer_0[857] = ~in[210]; 
    assign layer_0[858] = in[208]; 
    assign layer_0[859] = ~in[207] | (in[217] & in[207]); 
    assign layer_0[860] = in[217] | in[212]; 
    assign layer_0[861] = in[204]; 
    assign layer_0[862] = in[198] ^ in[208]; 
    assign layer_0[863] = 1'b0; 
    assign layer_0[864] = 1'b1; 
    assign layer_0[865] = 1'b1; 
    assign layer_0[866] = ~in[226] | (in[199] & in[226]); 
    assign layer_0[867] = ~in[232] | (in[232] & in[223]); 
    assign layer_0[868] = ~in[225]; 
    assign layer_0[869] = in[222]; 
    assign layer_0[870] = ~(in[203] & in[205]); 
    assign layer_0[871] = in[223] | in[224]; 
    assign layer_0[872] = ~in[218]; 
    assign layer_0[873] = in[226] & ~in[233]; 
    assign layer_0[874] = 1'b1; 
    assign layer_0[875] = ~(in[214] & in[207]); 
    assign layer_0[876] = in[227] & ~in[213]; 
    assign layer_0[877] = ~in[228]; 
    assign layer_0[878] = 1'b1; 
    assign layer_0[879] = ~in[223] | (in[223] & in[223]); 
    assign layer_0[880] = ~(in[214] | in[211]); 
    assign layer_0[881] = ~(in[229] | in[223]); 
    assign layer_0[882] = 1'b0; 
    assign layer_0[883] = in[220]; 
    assign layer_0[884] = in[236]; 
    assign layer_0[885] = in[228] ^ in[236]; 
    assign layer_0[886] = ~in[235] | (in[208] & in[235]); 
    assign layer_0[887] = in[215] & ~in[233]; 
    assign layer_0[888] = 1'b0; 
    assign layer_0[889] = ~(in[213] ^ in[206]); 
    assign layer_0[890] = in[229] & in[220]; 
    assign layer_0[891] = ~(in[233] & in[237]); 
    assign layer_0[892] = ~in[228] | (in[228] & in[206]); 
    assign layer_0[893] = 1'b0; 
    assign layer_0[894] = ~in[233] | (in[233] & in[208]); 
    assign layer_0[895] = in[235]; 
    assign layer_0[896] = ~in[225]; 
    assign layer_0[897] = ~(in[224] & in[209]); 
    assign layer_0[898] = in[215]; 
    assign layer_0[899] = in[230] & ~in[223]; 
    assign layer_0[900] = ~in[217]; 
    assign layer_0[901] = in[211] & in[208]; 
    assign layer_0[902] = in[216]; 
    assign layer_0[903] = in[225] | in[208]; 
    assign layer_0[904] = ~in[233]; 
    assign layer_0[905] = ~in[225] | (in[228] & in[225]); 
    assign layer_0[906] = in[234] & ~in[230]; 
    assign layer_0[907] = ~in[234] | (in[228] & in[234]); 
    assign layer_0[908] = in[235] & ~in[240]; 
    assign layer_0[909] = in[220] & ~in[228]; 
    assign layer_0[910] = in[242]; 
    assign layer_0[911] = ~(in[212] | in[233]); 
    assign layer_0[912] = in[224] & in[226]; 
    assign layer_0[913] = in[237] & in[213]; 
    assign layer_0[914] = in[237] & in[233]; 
    assign layer_0[915] = 1'b1; 
    assign layer_0[916] = ~in[244]; 
    assign layer_0[917] = in[230] & ~in[236]; 
    assign layer_0[918] = ~in[227] | (in[227] & in[212]); 
    assign layer_0[919] = ~in[223]; 
    assign layer_0[920] = in[236] & in[232]; 
    assign layer_0[921] = in[245] & in[228]; 
    assign layer_0[922] = ~in[226] | (in[238] & in[226]); 
    assign layer_0[923] = ~in[214]; 
    assign layer_0[924] = in[238] & ~in[237]; 
    assign layer_0[925] = ~(in[216] ^ in[214]); 
    assign layer_0[926] = in[225] ^ in[222]; 
    assign layer_0[927] = in[238] | in[240]; 
    assign layer_0[928] = in[237]; 
    assign layer_0[929] = in[239] | in[225]; 
    assign layer_0[930] = ~in[227] | (in[226] & in[227]); 
    assign layer_0[931] = in[232] ^ in[229]; 
    assign layer_0[932] = ~(in[217] ^ in[224]); 
    assign layer_0[933] = in[240] ^ in[219]; 
    assign layer_0[934] = ~in[229] | (in[229] & in[240]); 
    assign layer_0[935] = in[246]; 
    assign layer_0[936] = 1'b1; 
    assign layer_0[937] = in[224]; 
    assign layer_0[938] = ~(in[234] ^ in[224]); 
    assign layer_0[939] = in[221] & ~in[231]; 
    assign layer_0[940] = in[238] & ~in[247]; 
    assign layer_0[941] = in[219] ^ in[238]; 
    assign layer_0[942] = ~in[225]; 
    assign layer_0[943] = ~(in[232] & in[228]); 
    assign layer_0[944] = ~in[223] | (in[241] & in[223]); 
    assign layer_0[945] = ~in[236]; 
    assign layer_0[946] = ~(in[237] ^ in[238]); 
    assign layer_0[947] = in[244] | in[235]; 
    assign layer_0[948] = ~in[246] | (in[250] & in[246]); 
    assign layer_0[949] = in[241] & ~in[233]; 
    assign layer_0[950] = in[247] & ~in[239]; 
    assign layer_0[951] = 1'b0; 
    assign layer_0[952] = ~(in[234] | in[237]); 
    assign layer_0[953] = ~(in[230] | in[234]); 
    assign layer_0[954] = ~in[221] | (in[240] & in[221]); 
    assign layer_0[955] = in[227] & in[228]; 
    assign layer_0[956] = in[244]; 
    assign layer_0[957] = ~in[253] | (in[230] & in[253]); 
    assign layer_0[958] = 1'b0; 
    assign layer_0[959] = 1'b0; 
    assign layer_0[960] = ~in[230]; 
    assign layer_0[961] = in[248] | in[230]; 
    assign layer_0[962] = ~(in[249] | in[235]); 
    assign layer_0[963] = 1'b1; 
    assign layer_0[964] = ~in[224]; 
    assign layer_0[965] = 1'b0; 
    assign layer_0[966] = in[237] & in[235]; 
    assign layer_0[967] = ~in[227] | (in[227] & in[244]); 
    assign layer_0[968] = in[225]; 
    assign layer_0[969] = ~in[240] | (in[242] & in[240]); 
    assign layer_0[970] = in[255] & ~in[237]; 
    assign layer_0[971] = 1'b1; 
    assign layer_0[972] = 1'b0; 
    assign layer_0[973] = in[244] & ~in[251]; 
    assign layer_0[974] = in[255] | in[253]; 
    assign layer_0[975] = in[241] & in[237]; 
    assign layer_0[976] = ~in[247]; 
    assign layer_0[977] = in[252]; 
    assign layer_0[978] = in[239] | in[245]; 
    assign layer_0[979] = ~in[231]; 
    assign layer_0[980] = 1'b0; 
    assign layer_0[981] = in[231] | in[249]; 
    assign layer_0[982] = ~(in[230] | in[237]); 
    assign layer_0[983] = ~(in[234] & in[248]); 
    assign layer_0[984] = ~in[238]; 
    assign layer_0[985] = in[245] | in[253]; 
    assign layer_0[986] = ~(in[243] | in[244]); 
    assign layer_0[987] = in[255] | in[247]; 
    assign layer_0[988] = ~in[247] | (in[247] & in[250]); 
    assign layer_0[989] = in[248]; 
    assign layer_0[990] = ~(in[237] | in[233]); 
    assign layer_0[991] = ~in[247]; 
    assign layer_0[992] = ~(in[255] & in[235]); 
    assign layer_0[993] = ~in[246]; 
    assign layer_0[994] = 1'b1; 
    assign layer_0[995] = ~in[250]; 
    assign layer_0[996] = ~(in[240] & in[248]); 
    assign layer_0[997] = ~(in[249] ^ in[233]); 
    assign layer_0[998] = ~(in[243] ^ in[247]); 
    assign layer_0[999] = ~in[241]; 
    assign layer_0[1000] = ~in[252]; 
    assign layer_0[1001] = ~(in[238] | in[237]); 
    assign layer_0[1002] = in[245]; 
    assign layer_0[1003] = in[234] & ~in[252]; 
    assign layer_0[1004] = ~(in[237] & in[245]); 
    assign layer_0[1005] = 1'b0; 
    assign layer_0[1006] = in[255] | in[241]; 
    assign layer_0[1007] = in[252] ^ in[249]; 
    assign layer_0[1008] = in[246]; 
    assign layer_0[1009] = in[254] & ~in[239]; 
    assign layer_0[1010] = ~(in[251] & in[240]); 
    assign layer_0[1011] = ~in[251]; 
    assign layer_0[1012] = in[248]; 
    assign layer_0[1013] = in[238] & in[251]; 
    assign layer_0[1014] = in[242]; 
    assign layer_0[1015] = in[246] ^ in[240]; 
    assign layer_0[1016] = 1'b0; 
    assign layer_0[1017] = in[254] & in[248]; 
    assign layer_0[1018] = in[237] ^ in[247]; 
    assign layer_0[1019] = 1'b0; 
    assign layer_0[1020] = ~(in[253] & in[240]); 
    assign layer_0[1021] = 1'b1; 
    assign layer_0[1022] = ~in[243] | (in[253] & in[243]); 
    assign layer_0[1023] = ~in[246]; 
    // Layer 1 ============================================================
    assign layer_1[0] = layer_0[4] | layer_0[5]; 
    assign layer_1[1] = layer_0[12] & layer_0[15]; 
    assign layer_1[2] = ~(layer_0[9] ^ layer_0[9]); 
    assign layer_1[3] = layer_0[9] & ~layer_0[8]; 
    assign layer_1[4] = 1'b0; 
    assign layer_1[5] = layer_0[18]; 
    assign layer_1[6] = ~(layer_0[9] | layer_0[0]); 
    assign layer_1[7] = ~(layer_0[22] & layer_0[9]); 
    assign layer_1[8] = layer_0[23] & ~layer_0[20]; 
    assign layer_1[9] = layer_0[7] & layer_0[20]; 
    assign layer_1[10] = ~layer_0[14]; 
    assign layer_1[11] = ~(layer_0[27] | layer_0[5]); 
    assign layer_1[12] = layer_0[12]; 
    assign layer_1[13] = layer_0[0] & ~layer_0[23]; 
    assign layer_1[14] = layer_0[30]; 
    assign layer_1[15] = 1'b0; 
    assign layer_1[16] = layer_0[3] & layer_0[20]; 
    assign layer_1[17] = layer_0[25] & layer_0[2]; 
    assign layer_1[18] = 1'b0; 
    assign layer_1[19] = ~(layer_0[25] ^ layer_0[25]); 
    assign layer_1[20] = ~layer_0[18]; 
    assign layer_1[21] = ~layer_0[8] | (layer_0[8] & layer_0[27]); 
    assign layer_1[22] = ~layer_0[23]; 
    assign layer_1[23] = layer_0[9]; 
    assign layer_1[24] = layer_0[23] ^ layer_0[11]; 
    assign layer_1[25] = layer_0[33]; 
    assign layer_1[26] = ~(layer_0[42] | layer_0[25]); 
    assign layer_1[27] = ~layer_0[37] | (layer_0[37] & layer_0[31]); 
    assign layer_1[28] = layer_0[43] ^ layer_0[30]; 
    assign layer_1[29] = layer_0[19] ^ layer_0[19]; 
    assign layer_1[30] = ~(layer_0[39] | layer_0[14]); 
    assign layer_1[31] = layer_0[33] | layer_0[29]; 
    assign layer_1[32] = layer_0[27]; 
    assign layer_1[33] = layer_0[33]; 
    assign layer_1[34] = 1'b1; 
    assign layer_1[35] = layer_0[37] & ~layer_0[27]; 
    assign layer_1[36] = ~layer_0[37]; 
    assign layer_1[37] = 1'b1; 
    assign layer_1[38] = layer_0[32] & ~layer_0[29]; 
    assign layer_1[39] = ~layer_0[30]; 
    assign layer_1[40] = layer_0[33] ^ layer_0[40]; 
    assign layer_1[41] = layer_0[26] & layer_0[37]; 
    assign layer_1[42] = ~(layer_0[35] | layer_0[29]); 
    assign layer_1[43] = ~(layer_0[31] & layer_0[30]); 
    assign layer_1[44] = ~(layer_0[60] & layer_0[43]); 
    assign layer_1[45] = ~layer_0[55]; 
    assign layer_1[46] = ~layer_0[59] | (layer_0[59] & layer_0[44]); 
    assign layer_1[47] = layer_0[34] | layer_0[59]; 
    assign layer_1[48] = layer_0[41]; 
    assign layer_1[49] = layer_0[49] & layer_0[33]; 
    assign layer_1[50] = layer_0[42]; 
    assign layer_1[51] = layer_0[65] & ~layer_0[58]; 
    assign layer_1[52] = ~layer_0[39]; 
    assign layer_1[53] = layer_0[52] & ~layer_0[47]; 
    assign layer_1[54] = layer_0[56] & ~layer_0[49]; 
    assign layer_1[55] = ~(layer_0[71] & layer_0[56]); 
    assign layer_1[56] = ~(layer_0[70] ^ layer_0[67]); 
    assign layer_1[57] = 1'b1; 
    assign layer_1[58] = ~layer_0[56] | (layer_0[72] & layer_0[56]); 
    assign layer_1[59] = layer_0[44]; 
    assign layer_1[60] = layer_0[60] & ~layer_0[45]; 
    assign layer_1[61] = layer_0[77] & layer_0[57]; 
    assign layer_1[62] = layer_0[54] | layer_0[54]; 
    assign layer_1[63] = ~layer_0[51] | (layer_0[51] & layer_0[51]); 
    assign layer_1[64] = layer_0[74] | layer_0[54]; 
    assign layer_1[65] = layer_0[70]; 
    assign layer_1[66] = ~layer_0[64] | (layer_0[73] & layer_0[64]); 
    assign layer_1[67] = layer_0[52]; 
    assign layer_1[68] = layer_0[80] & layer_0[80]; 
    assign layer_1[69] = layer_0[80] & layer_0[56]; 
    assign layer_1[70] = ~layer_0[77]; 
    assign layer_1[71] = ~(layer_0[80] | layer_0[64]); 
    assign layer_1[72] = 1'b0; 
    assign layer_1[73] = layer_0[61]; 
    assign layer_1[74] = 1'b0; 
    assign layer_1[75] = layer_0[87] & layer_0[87]; 
    assign layer_1[76] = layer_0[74] | layer_0[66]; 
    assign layer_1[77] = ~(layer_0[69] & layer_0[73]); 
    assign layer_1[78] = ~(layer_0[84] & layer_0[62]); 
    assign layer_1[79] = ~layer_0[78]; 
    assign layer_1[80] = 1'b0; 
    assign layer_1[81] = ~(layer_0[96] ^ layer_0[89]); 
    assign layer_1[82] = ~(layer_0[95] & layer_0[81]); 
    assign layer_1[83] = ~(layer_0[85] & layer_0[70]); 
    assign layer_1[84] = ~layer_0[94] | (layer_0[88] & layer_0[94]); 
    assign layer_1[85] = 1'b1; 
    assign layer_1[86] = layer_0[70] | layer_0[101]; 
    assign layer_1[87] = ~(layer_0[99] ^ layer_0[90]); 
    assign layer_1[88] = layer_0[76] & layer_0[101]; 
    assign layer_1[89] = layer_0[84]; 
    assign layer_1[90] = ~(layer_0[84] & layer_0[73]); 
    assign layer_1[91] = layer_0[86] & ~layer_0[104]; 
    assign layer_1[92] = layer_0[100]; 
    assign layer_1[93] = layer_0[104]; 
    assign layer_1[94] = 1'b0; 
    assign layer_1[95] = layer_0[89]; 
    assign layer_1[96] = 1'b1; 
    assign layer_1[97] = layer_0[102] & ~layer_0[102]; 
    assign layer_1[98] = layer_0[108] | layer_0[100]; 
    assign layer_1[99] = ~layer_0[82] | (layer_0[106] & layer_0[82]); 
    assign layer_1[100] = ~(layer_0[94] ^ layer_0[88]); 
    assign layer_1[101] = ~layer_0[107]; 
    assign layer_1[102] = ~layer_0[98] | (layer_0[104] & layer_0[98]); 
    assign layer_1[103] = layer_0[97] & ~layer_0[87]; 
    assign layer_1[104] = layer_0[115]; 
    assign layer_1[105] = layer_0[115] & ~layer_0[102]; 
    assign layer_1[106] = ~layer_0[92]; 
    assign layer_1[107] = layer_0[105] & ~layer_0[118]; 
    assign layer_1[108] = ~layer_0[119] | (layer_0[119] & layer_0[102]); 
    assign layer_1[109] = ~(layer_0[102] | layer_0[104]); 
    assign layer_1[110] = 1'b1; 
    assign layer_1[111] = ~layer_0[118] | (layer_0[118] & layer_0[123]); 
    assign layer_1[112] = layer_0[102] | layer_0[101]; 
    assign layer_1[113] = ~layer_0[103] | (layer_0[126] & layer_0[103]); 
    assign layer_1[114] = 1'b0; 
    assign layer_1[115] = layer_0[113] & layer_0[113]; 
    assign layer_1[116] = layer_0[130] & ~layer_0[129]; 
    assign layer_1[117] = layer_0[121] | layer_0[110]; 
    assign layer_1[118] = layer_0[108] & ~layer_0[102]; 
    assign layer_1[119] = 1'b0; 
    assign layer_1[120] = layer_0[116] & ~layer_0[120]; 
    assign layer_1[121] = 1'b0; 
    assign layer_1[122] = ~layer_0[125] | (layer_0[122] & layer_0[125]); 
    assign layer_1[123] = ~layer_0[118]; 
    assign layer_1[124] = ~layer_0[132]; 
    assign layer_1[125] = layer_0[140] | layer_0[121]; 
    assign layer_1[126] = ~layer_0[116]; 
    assign layer_1[127] = ~layer_0[122] | (layer_0[122] & layer_0[115]); 
    assign layer_1[128] = ~layer_0[112]; 
    assign layer_1[129] = layer_0[145] ^ layer_0[144]; 
    assign layer_1[130] = 1'b0; 
    assign layer_1[131] = layer_0[140] ^ layer_0[116]; 
    assign layer_1[132] = 1'b1; 
    assign layer_1[133] = ~layer_0[148]; 
    assign layer_1[134] = 1'b0; 
    assign layer_1[135] = layer_0[128]; 
    assign layer_1[136] = ~(layer_0[124] ^ layer_0[130]); 
    assign layer_1[137] = layer_0[123]; 
    assign layer_1[138] = layer_0[151] & layer_0[129]; 
    assign layer_1[139] = ~layer_0[150] | (layer_0[150] & layer_0[148]); 
    assign layer_1[140] = layer_0[152]; 
    assign layer_1[141] = layer_0[126] & ~layer_0[125]; 
    assign layer_1[142] = layer_0[137] & layer_0[152]; 
    assign layer_1[143] = layer_0[133]; 
    assign layer_1[144] = ~layer_0[153] | (layer_0[153] & layer_0[128]); 
    assign layer_1[145] = ~layer_0[142] | (layer_0[149] & layer_0[142]); 
    assign layer_1[146] = layer_0[141] & ~layer_0[147]; 
    assign layer_1[147] = ~(layer_0[135] ^ layer_0[161]); 
    assign layer_1[148] = ~(layer_0[161] ^ layer_0[159]); 
    assign layer_1[149] = ~layer_0[150]; 
    assign layer_1[150] = ~layer_0[165] | (layer_0[165] & layer_0[165]); 
    assign layer_1[151] = layer_0[155] & ~layer_0[142]; 
    assign layer_1[152] = ~layer_0[151]; 
    assign layer_1[153] = layer_0[141] ^ layer_0[150]; 
    assign layer_1[154] = layer_0[166]; 
    assign layer_1[155] = layer_0[156] & layer_0[146]; 
    assign layer_1[156] = ~layer_0[164] | (layer_0[146] & layer_0[164]); 
    assign layer_1[157] = ~layer_0[150]; 
    assign layer_1[158] = 1'b0; 
    assign layer_1[159] = layer_0[154] & ~layer_0[173]; 
    assign layer_1[160] = ~layer_0[176] | (layer_0[176] & layer_0[172]); 
    assign layer_1[161] = 1'b1; 
    assign layer_1[162] = ~layer_0[151]; 
    assign layer_1[163] = ~layer_0[154]; 
    assign layer_1[164] = layer_0[157] & layer_0[167]; 
    assign layer_1[165] = layer_0[156] & layer_0[153]; 
    assign layer_1[166] = layer_0[168] & ~layer_0[171]; 
    assign layer_1[167] = layer_0[169]; 
    assign layer_1[168] = layer_0[160] & ~layer_0[179]; 
    assign layer_1[169] = layer_0[159]; 
    assign layer_1[170] = layer_0[177]; 
    assign layer_1[171] = layer_0[180] & layer_0[175]; 
    assign layer_1[172] = layer_0[161]; 
    assign layer_1[173] = ~layer_0[175] | (layer_0[175] & layer_0[168]); 
    assign layer_1[174] = 1'b0; 
    assign layer_1[175] = layer_0[183] & layer_0[187]; 
    assign layer_1[176] = layer_0[189] & layer_0[181]; 
    assign layer_1[177] = layer_0[190] & layer_0[175]; 
    assign layer_1[178] = layer_0[189]; 
    assign layer_1[179] = layer_0[173]; 
    assign layer_1[180] = layer_0[179] & ~layer_0[165]; 
    assign layer_1[181] = ~layer_0[184]; 
    assign layer_1[182] = ~layer_0[167]; 
    assign layer_1[183] = ~(layer_0[194] & layer_0[186]); 
    assign layer_1[184] = layer_0[174] & ~layer_0[191]; 
    assign layer_1[185] = ~(layer_0[185] ^ layer_0[183]); 
    assign layer_1[186] = 1'b0; 
    assign layer_1[187] = layer_0[185] & layer_0[172]; 
    assign layer_1[188] = layer_0[181]; 
    assign layer_1[189] = ~(layer_0[175] | layer_0[181]); 
    assign layer_1[190] = layer_0[174] & ~layer_0[203]; 
    assign layer_1[191] = ~(layer_0[175] | layer_0[191]); 
    assign layer_1[192] = layer_0[180] & ~layer_0[196]; 
    assign layer_1[193] = ~layer_0[195]; 
    assign layer_1[194] = layer_0[201]; 
    assign layer_1[195] = 1'b1; 
    assign layer_1[196] = ~layer_0[204]; 
    assign layer_1[197] = layer_0[203] | layer_0[187]; 
    assign layer_1[198] = layer_0[212] & ~layer_0[182]; 
    assign layer_1[199] = ~layer_0[198]; 
    assign layer_1[200] = layer_0[198] ^ layer_0[214]; 
    assign layer_1[201] = 1'b0; 
    assign layer_1[202] = layer_0[207] & ~layer_0[198]; 
    assign layer_1[203] = ~layer_0[197] | (layer_0[197] & layer_0[213]); 
    assign layer_1[204] = layer_0[217] ^ layer_0[201]; 
    assign layer_1[205] = ~(layer_0[217] | layer_0[210]); 
    assign layer_1[206] = 1'b1; 
    assign layer_1[207] = layer_0[194] & ~layer_0[210]; 
    assign layer_1[208] = ~layer_0[199] | (layer_0[211] & layer_0[199]); 
    assign layer_1[209] = layer_0[223] | layer_0[208]; 
    assign layer_1[210] = ~(layer_0[222] ^ layer_0[214]); 
    assign layer_1[211] = layer_0[195] & ~layer_0[207]; 
    assign layer_1[212] = 1'b0; 
    assign layer_1[213] = layer_0[213]; 
    assign layer_1[214] = layer_0[229] | layer_0[203]; 
    assign layer_1[215] = layer_0[209]; 
    assign layer_1[216] = 1'b1; 
    assign layer_1[217] = layer_0[232] | layer_0[208]; 
    assign layer_1[218] = ~(layer_0[222] & layer_0[220]); 
    assign layer_1[219] = ~(layer_0[209] & layer_0[207]); 
    assign layer_1[220] = ~layer_0[213] | (layer_0[213] & layer_0[226]); 
    assign layer_1[221] = ~layer_0[231]; 
    assign layer_1[222] = ~(layer_0[213] ^ layer_0[237]); 
    assign layer_1[223] = ~(layer_0[215] ^ layer_0[208]); 
    assign layer_1[224] = ~layer_0[209] | (layer_0[237] & layer_0[209]); 
    assign layer_1[225] = layer_0[237] ^ layer_0[216]; 
    assign layer_1[226] = layer_0[210] | layer_0[232]; 
    assign layer_1[227] = ~layer_0[242] | (layer_0[242] & layer_0[228]); 
    assign layer_1[228] = ~layer_0[243] | (layer_0[217] & layer_0[243]); 
    assign layer_1[229] = ~(layer_0[229] & layer_0[241]); 
    assign layer_1[230] = ~layer_0[228]; 
    assign layer_1[231] = layer_0[233]; 
    assign layer_1[232] = ~layer_0[219] | (layer_0[248] & layer_0[219]); 
    assign layer_1[233] = layer_0[229] & layer_0[230]; 
    assign layer_1[234] = 1'b1; 
    assign layer_1[235] = ~(layer_0[227] & layer_0[229]); 
    assign layer_1[236] = ~layer_0[243] | (layer_0[243] & layer_0[242]); 
    assign layer_1[237] = layer_0[231] & layer_0[242]; 
    assign layer_1[238] = 1'b0; 
    assign layer_1[239] = ~(layer_0[228] | layer_0[230]); 
    assign layer_1[240] = ~layer_0[230] | (layer_0[225] & layer_0[230]); 
    assign layer_1[241] = layer_0[227] & ~layer_0[229]; 
    assign layer_1[242] = layer_0[241] & layer_0[254]; 
    assign layer_1[243] = layer_0[247] ^ layer_0[240]; 
    assign layer_1[244] = layer_0[258]; 
    assign layer_1[245] = 1'b0; 
    assign layer_1[246] = layer_0[259] & layer_0[253]; 
    assign layer_1[247] = layer_0[245] | layer_0[241]; 
    assign layer_1[248] = layer_0[258] & ~layer_0[252]; 
    assign layer_1[249] = ~(layer_0[246] ^ layer_0[244]); 
    assign layer_1[250] = ~layer_0[252] | (layer_0[252] & layer_0[265]); 
    assign layer_1[251] = 1'b0; 
    assign layer_1[252] = layer_0[251] | layer_0[261]; 
    assign layer_1[253] = ~layer_0[251]; 
    assign layer_1[254] = layer_0[263]; 
    assign layer_1[255] = 1'b0; 
    assign layer_1[256] = layer_0[268]; 
    assign layer_1[257] = layer_0[261] & ~layer_0[256]; 
    assign layer_1[258] = layer_0[273] & ~layer_0[244]; 
    assign layer_1[259] = ~(layer_0[264] | layer_0[268]); 
    assign layer_1[260] = ~layer_0[267]; 
    assign layer_1[261] = ~layer_0[271] | (layer_0[271] & layer_0[258]); 
    assign layer_1[262] = ~layer_0[273]; 
    assign layer_1[263] = ~(layer_0[256] | layer_0[275]); 
    assign layer_1[264] = layer_0[264]; 
    assign layer_1[265] = 1'b0; 
    assign layer_1[266] = ~(layer_0[259] ^ layer_0[258]); 
    assign layer_1[267] = layer_0[270] & layer_0[264]; 
    assign layer_1[268] = layer_0[260] ^ layer_0[276]; 
    assign layer_1[269] = layer_0[265] ^ layer_0[268]; 
    assign layer_1[270] = 1'b1; 
    assign layer_1[271] = layer_0[259] ^ layer_0[257]; 
    assign layer_1[272] = layer_0[283] & ~layer_0[267]; 
    assign layer_1[273] = layer_0[285] & ~layer_0[280]; 
    assign layer_1[274] = ~layer_0[268]; 
    assign layer_1[275] = layer_0[278] & ~layer_0[273]; 
    assign layer_1[276] = ~layer_0[262]; 
    assign layer_1[277] = layer_0[264] & layer_0[264]; 
    assign layer_1[278] = ~layer_0[277]; 
    assign layer_1[279] = ~layer_0[282] | (layer_0[283] & layer_0[282]); 
    assign layer_1[280] = layer_0[282]; 
    assign layer_1[281] = ~(layer_0[294] ^ layer_0[282]); 
    assign layer_1[282] = ~(layer_0[267] ^ layer_0[289]); 
    assign layer_1[283] = ~(layer_0[293] | layer_0[288]); 
    assign layer_1[284] = layer_0[296] & ~layer_0[284]; 
    assign layer_1[285] = layer_0[294] & ~layer_0[299]; 
    assign layer_1[286] = layer_0[300] & ~layer_0[270]; 
    assign layer_1[287] = layer_0[286] ^ layer_0[296]; 
    assign layer_1[288] = layer_0[284] | layer_0[292]; 
    assign layer_1[289] = layer_0[304] & layer_0[291]; 
    assign layer_1[290] = ~(layer_0[292] | layer_0[290]); 
    assign layer_1[291] = ~layer_0[301] | (layer_0[301] & layer_0[299]); 
    assign layer_1[292] = layer_0[282] & ~layer_0[278]; 
    assign layer_1[293] = 1'b0; 
    assign layer_1[294] = 1'b1; 
    assign layer_1[295] = 1'b1; 
    assign layer_1[296] = layer_0[288] & ~layer_0[294]; 
    assign layer_1[297] = ~layer_0[292] | (layer_0[312] & layer_0[292]); 
    assign layer_1[298] = 1'b0; 
    assign layer_1[299] = ~layer_0[298] | (layer_0[298] & layer_0[284]); 
    assign layer_1[300] = layer_0[298] ^ layer_0[303]; 
    assign layer_1[301] = 1'b0; 
    assign layer_1[302] = ~(layer_0[293] & layer_0[314]); 
    assign layer_1[303] = layer_0[299] & layer_0[315]; 
    assign layer_1[304] = layer_0[312] | layer_0[318]; 
    assign layer_1[305] = layer_0[297] ^ layer_0[316]; 
    assign layer_1[306] = 1'b1; 
    assign layer_1[307] = ~layer_0[304]; 
    assign layer_1[308] = ~(layer_0[317] ^ layer_0[304]); 
    assign layer_1[309] = ~layer_0[304] | (layer_0[322] & layer_0[304]); 
    assign layer_1[310] = layer_0[300]; 
    assign layer_1[311] = ~(layer_0[317] | layer_0[321]); 
    assign layer_1[312] = ~(layer_0[325] & layer_0[321]); 
    assign layer_1[313] = layer_0[315] | layer_0[305]; 
    assign layer_1[314] = ~(layer_0[302] | layer_0[308]); 
    assign layer_1[315] = ~layer_0[315]; 
    assign layer_1[316] = 1'b1; 
    assign layer_1[317] = layer_0[306] & layer_0[325]; 
    assign layer_1[318] = ~(layer_0[320] ^ layer_0[319]); 
    assign layer_1[319] = layer_0[325] & ~layer_0[331]; 
    assign layer_1[320] = layer_0[322]; 
    assign layer_1[321] = ~(layer_0[305] & layer_0[336]); 
    assign layer_1[322] = layer_0[316] | layer_0[311]; 
    assign layer_1[323] = ~(layer_0[324] & layer_0[319]); 
    assign layer_1[324] = ~layer_0[327] | (layer_0[327] & layer_0[314]); 
    assign layer_1[325] = ~layer_0[339] | (layer_0[339] & layer_0[337]); 
    assign layer_1[326] = ~layer_0[323]; 
    assign layer_1[327] = layer_0[341] | layer_0[312]; 
    assign layer_1[328] = ~layer_0[342] | (layer_0[342] & layer_0[334]); 
    assign layer_1[329] = layer_0[315] & ~layer_0[323]; 
    assign layer_1[330] = layer_0[341] | layer_0[328]; 
    assign layer_1[331] = ~(layer_0[334] | layer_0[343]); 
    assign layer_1[332] = ~(layer_0[319] ^ layer_0[324]); 
    assign layer_1[333] = ~layer_0[327] | (layer_0[349] & layer_0[327]); 
    assign layer_1[334] = ~(layer_0[319] ^ layer_0[320]); 
    assign layer_1[335] = ~layer_0[323] | (layer_0[323] & layer_0[349]); 
    assign layer_1[336] = layer_0[340] & layer_0[325]; 
    assign layer_1[337] = ~layer_0[322] | (layer_0[349] & layer_0[322]); 
    assign layer_1[338] = ~(layer_0[344] | layer_0[339]); 
    assign layer_1[339] = layer_0[344]; 
    assign layer_1[340] = ~layer_0[345]; 
    assign layer_1[341] = layer_0[325] ^ layer_0[332]; 
    assign layer_1[342] = layer_0[348] & ~layer_0[346]; 
    assign layer_1[343] = 1'b0; 
    assign layer_1[344] = layer_0[334]; 
    assign layer_1[345] = ~(layer_0[330] & layer_0[335]); 
    assign layer_1[346] = ~layer_0[361] | (layer_0[359] & layer_0[361]); 
    assign layer_1[347] = ~(layer_0[362] & layer_0[351]); 
    assign layer_1[348] = layer_0[338] & layer_0[347]; 
    assign layer_1[349] = layer_0[349]; 
    assign layer_1[350] = layer_0[363] & ~layer_0[355]; 
    assign layer_1[351] = ~(layer_0[344] ^ layer_0[341]); 
    assign layer_1[352] = ~layer_0[339]; 
    assign layer_1[353] = ~(layer_0[344] | layer_0[351]); 
    assign layer_1[354] = ~(layer_0[368] ^ layer_0[356]); 
    assign layer_1[355] = ~layer_0[368]; 
    assign layer_1[356] = ~(layer_0[372] & layer_0[343]); 
    assign layer_1[357] = layer_0[342] | layer_0[370]; 
    assign layer_1[358] = ~layer_0[342] | (layer_0[359] & layer_0[342]); 
    assign layer_1[359] = ~(layer_0[366] ^ layer_0[342]); 
    assign layer_1[360] = layer_0[348]; 
    assign layer_1[361] = layer_0[377] & layer_0[355]; 
    assign layer_1[362] = 1'b0; 
    assign layer_1[363] = 1'b1; 
    assign layer_1[364] = ~layer_0[375]; 
    assign layer_1[365] = layer_0[349]; 
    assign layer_1[366] = ~layer_0[358]; 
    assign layer_1[367] = ~layer_0[358]; 
    assign layer_1[368] = ~(layer_0[382] | layer_0[352]); 
    assign layer_1[369] = ~layer_0[361]; 
    assign layer_1[370] = 1'b1; 
    assign layer_1[371] = ~layer_0[387]; 
    assign layer_1[372] = ~(layer_0[363] & layer_0[357]); 
    assign layer_1[373] = ~(layer_0[375] | layer_0[374]); 
    assign layer_1[374] = ~layer_0[374] | (layer_0[374] & layer_0[388]); 
    assign layer_1[375] = 1'b0; 
    assign layer_1[376] = ~layer_0[381]; 
    assign layer_1[377] = layer_0[364] | layer_0[369]; 
    assign layer_1[378] = ~layer_0[386] | (layer_0[386] & layer_0[386]); 
    assign layer_1[379] = 1'b1; 
    assign layer_1[380] = ~layer_0[380] | (layer_0[380] & layer_0[384]); 
    assign layer_1[381] = layer_0[390] & ~layer_0[383]; 
    assign layer_1[382] = layer_0[370] & layer_0[393]; 
    assign layer_1[383] = ~layer_0[381]; 
    assign layer_1[384] = layer_0[368] & ~layer_0[396]; 
    assign layer_1[385] = layer_0[382]; 
    assign layer_1[386] = ~layer_0[389] | (layer_0[375] & layer_0[389]); 
    assign layer_1[387] = layer_0[399]; 
    assign layer_1[388] = layer_0[391] & ~layer_0[373]; 
    assign layer_1[389] = layer_0[390]; 
    assign layer_1[390] = 1'b1; 
    assign layer_1[391] = layer_0[400] | layer_0[396]; 
    assign layer_1[392] = ~layer_0[386] | (layer_0[407] & layer_0[386]); 
    assign layer_1[393] = ~(layer_0[403] | layer_0[405]); 
    assign layer_1[394] = ~(layer_0[404] ^ layer_0[381]); 
    assign layer_1[395] = ~layer_0[401]; 
    assign layer_1[396] = ~layer_0[401] | (layer_0[408] & layer_0[401]); 
    assign layer_1[397] = ~(layer_0[394] ^ layer_0[410]); 
    assign layer_1[398] = layer_0[412] & layer_0[407]; 
    assign layer_1[399] = ~layer_0[399] | (layer_0[399] & layer_0[405]); 
    assign layer_1[400] = layer_0[408] ^ layer_0[405]; 
    assign layer_1[401] = layer_0[410]; 
    assign layer_1[402] = 1'b1; 
    assign layer_1[403] = layer_0[406] & ~layer_0[403]; 
    assign layer_1[404] = layer_0[393]; 
    assign layer_1[405] = layer_0[401] & ~layer_0[397]; 
    assign layer_1[406] = layer_0[420]; 
    assign layer_1[407] = layer_0[391] | layer_0[414]; 
    assign layer_1[408] = layer_0[393]; 
    assign layer_1[409] = ~layer_0[394]; 
    assign layer_1[410] = ~(layer_0[399] | layer_0[409]); 
    assign layer_1[411] = layer_0[410] & layer_0[408]; 
    assign layer_1[412] = layer_0[417]; 
    assign layer_1[413] = ~(layer_0[399] & layer_0[423]); 
    assign layer_1[414] = ~(layer_0[420] | layer_0[424]); 
    assign layer_1[415] = 1'b1; 
    assign layer_1[416] = layer_0[417] & ~layer_0[422]; 
    assign layer_1[417] = layer_0[424] ^ layer_0[408]; 
    assign layer_1[418] = layer_0[413] | layer_0[417]; 
    assign layer_1[419] = ~(layer_0[404] & layer_0[406]); 
    assign layer_1[420] = layer_0[428] & ~layer_0[435]; 
    assign layer_1[421] = ~layer_0[407]; 
    assign layer_1[422] = 1'b1; 
    assign layer_1[423] = ~layer_0[426] | (layer_0[437] & layer_0[426]); 
    assign layer_1[424] = layer_0[439]; 
    assign layer_1[425] = ~layer_0[427] | (layer_0[424] & layer_0[427]); 
    assign layer_1[426] = layer_0[416] & layer_0[430]; 
    assign layer_1[427] = ~layer_0[436]; 
    assign layer_1[428] = layer_0[428]; 
    assign layer_1[429] = ~layer_0[430]; 
    assign layer_1[430] = ~layer_0[422] | (layer_0[422] & layer_0[417]); 
    assign layer_1[431] = layer_0[438] & ~layer_0[433]; 
    assign layer_1[432] = ~layer_0[447]; 
    assign layer_1[433] = ~(layer_0[417] ^ layer_0[435]); 
    assign layer_1[434] = 1'b1; 
    assign layer_1[435] = layer_0[448] & ~layer_0[446]; 
    assign layer_1[436] = ~layer_0[423]; 
    assign layer_1[437] = layer_0[431] | layer_0[422]; 
    assign layer_1[438] = layer_0[438] & ~layer_0[441]; 
    assign layer_1[439] = ~(layer_0[445] & layer_0[452]); 
    assign layer_1[440] = ~layer_0[438] | (layer_0[438] & layer_0[442]); 
    assign layer_1[441] = 1'b1; 
    assign layer_1[442] = layer_0[448] ^ layer_0[426]; 
    assign layer_1[443] = ~layer_0[452]; 
    assign layer_1[444] = ~(layer_0[450] | layer_0[459]); 
    assign layer_1[445] = layer_0[446]; 
    assign layer_1[446] = layer_0[446] & ~layer_0[440]; 
    assign layer_1[447] = ~(layer_0[457] ^ layer_0[444]); 
    assign layer_1[448] = 1'b1; 
    assign layer_1[449] = ~(layer_0[450] | layer_0[449]); 
    assign layer_1[450] = ~layer_0[443] | (layer_0[451] & layer_0[443]); 
    assign layer_1[451] = ~(layer_0[442] & layer_0[466]); 
    assign layer_1[452] = ~layer_0[452]; 
    assign layer_1[453] = ~(layer_0[458] | layer_0[458]); 
    assign layer_1[454] = ~(layer_0[440] | layer_0[456]); 
    assign layer_1[455] = layer_0[469] ^ layer_0[455]; 
    assign layer_1[456] = layer_0[463] & ~layer_0[445]; 
    assign layer_1[457] = ~layer_0[453]; 
    assign layer_1[458] = layer_0[459] & ~layer_0[446]; 
    assign layer_1[459] = layer_0[467] ^ layer_0[449]; 
    assign layer_1[460] = 1'b1; 
    assign layer_1[461] = ~(layer_0[447] ^ layer_0[455]); 
    assign layer_1[462] = layer_0[454] & ~layer_0[457]; 
    assign layer_1[463] = layer_0[470] | layer_0[458]; 
    assign layer_1[464] = layer_0[462]; 
    assign layer_1[465] = 1'b1; 
    assign layer_1[466] = 1'b1; 
    assign layer_1[467] = ~layer_0[472] | (layer_0[472] & layer_0[473]); 
    assign layer_1[468] = layer_0[454] | layer_0[474]; 
    assign layer_1[469] = ~layer_0[482]; 
    assign layer_1[470] = ~(layer_0[455] & layer_0[460]); 
    assign layer_1[471] = layer_0[482]; 
    assign layer_1[472] = ~layer_0[457] | (layer_0[471] & layer_0[457]); 
    assign layer_1[473] = layer_0[464] | layer_0[458]; 
    assign layer_1[474] = 1'b1; 
    assign layer_1[475] = layer_0[482] & layer_0[460]; 
    assign layer_1[476] = ~(layer_0[475] ^ layer_0[487]); 
    assign layer_1[477] = ~(layer_0[462] | layer_0[463]); 
    assign layer_1[478] = layer_0[493]; 
    assign layer_1[479] = layer_0[494] & ~layer_0[486]; 
    assign layer_1[480] = ~layer_0[490] | (layer_0[470] & layer_0[490]); 
    assign layer_1[481] = 1'b1; 
    assign layer_1[482] = layer_0[484] ^ layer_0[495]; 
    assign layer_1[483] = layer_0[491] | layer_0[498]; 
    assign layer_1[484] = layer_0[483]; 
    assign layer_1[485] = layer_0[473] & ~layer_0[473]; 
    assign layer_1[486] = ~layer_0[476] | (layer_0[481] & layer_0[476]); 
    assign layer_1[487] = layer_0[488] & layer_0[494]; 
    assign layer_1[488] = ~(layer_0[494] & layer_0[503]); 
    assign layer_1[489] = ~(layer_0[490] ^ layer_0[499]); 
    assign layer_1[490] = layer_0[500] ^ layer_0[495]; 
    assign layer_1[491] = layer_0[484] ^ layer_0[488]; 
    assign layer_1[492] = ~(layer_0[495] & layer_0[506]); 
    assign layer_1[493] = layer_0[485] & layer_0[484]; 
    assign layer_1[494] = layer_0[494] & ~layer_0[501]; 
    assign layer_1[495] = layer_0[508] & ~layer_0[487]; 
    assign layer_1[496] = ~layer_0[499]; 
    assign layer_1[497] = ~layer_0[499]; 
    assign layer_1[498] = layer_0[488] ^ layer_0[508]; 
    assign layer_1[499] = layer_0[506] & ~layer_0[491]; 
    assign layer_1[500] = ~(layer_0[497] & layer_0[495]); 
    assign layer_1[501] = layer_0[496]; 
    assign layer_1[502] = layer_0[498]; 
    assign layer_1[503] = layer_0[498] & layer_0[512]; 
    assign layer_1[504] = layer_0[490] & ~layer_0[507]; 
    assign layer_1[505] = layer_0[502] & ~layer_0[515]; 
    assign layer_1[506] = layer_0[518] | layer_0[495]; 
    assign layer_1[507] = ~(layer_0[491] ^ layer_0[500]); 
    assign layer_1[508] = ~(layer_0[514] | layer_0[510]); 
    assign layer_1[509] = layer_0[507] & ~layer_0[516]; 
    assign layer_1[510] = layer_0[508] | layer_0[505]; 
    assign layer_1[511] = layer_0[513]; 
    assign layer_1[512] = layer_0[527] & ~layer_0[501]; 
    assign layer_1[513] = 1'b1; 
    assign layer_1[514] = ~layer_0[529] | (layer_0[504] & layer_0[529]); 
    assign layer_1[515] = ~layer_0[506]; 
    assign layer_1[516] = ~(layer_0[526] | layer_0[506]); 
    assign layer_1[517] = ~layer_0[519]; 
    assign layer_1[518] = ~(layer_0[502] ^ layer_0[505]); 
    assign layer_1[519] = ~layer_0[524]; 
    assign layer_1[520] = ~layer_0[505]; 
    assign layer_1[521] = layer_0[537] & ~layer_0[516]; 
    assign layer_1[522] = ~(layer_0[529] & layer_0[514]); 
    assign layer_1[523] = ~layer_0[536]; 
    assign layer_1[524] = ~layer_0[528]; 
    assign layer_1[525] = ~layer_0[513]; 
    assign layer_1[526] = ~layer_0[522] | (layer_0[525] & layer_0[522]); 
    assign layer_1[527] = ~(layer_0[514] & layer_0[524]); 
    assign layer_1[528] = ~layer_0[531]; 
    assign layer_1[529] = ~layer_0[520]; 
    assign layer_1[530] = layer_0[521] ^ layer_0[527]; 
    assign layer_1[531] = layer_0[533] ^ layer_0[514]; 
    assign layer_1[532] = layer_0[538] & ~layer_0[520]; 
    assign layer_1[533] = ~layer_0[537] | (layer_0[537] & layer_0[532]); 
    assign layer_1[534] = layer_0[534] ^ layer_0[543]; 
    assign layer_1[535] = ~layer_0[529]; 
    assign layer_1[536] = layer_0[538] & layer_0[534]; 
    assign layer_1[537] = layer_0[551]; 
    assign layer_1[538] = ~(layer_0[551] & layer_0[539]); 
    assign layer_1[539] = 1'b1; 
    assign layer_1[540] = ~(layer_0[543] | layer_0[547]); 
    assign layer_1[541] = layer_0[545] & ~layer_0[555]; 
    assign layer_1[542] = ~layer_0[543] | (layer_0[543] & layer_0[535]); 
    assign layer_1[543] = 1'b0; 
    assign layer_1[544] = ~(layer_0[550] | layer_0[554]); 
    assign layer_1[545] = layer_0[545] ^ layer_0[534]; 
    assign layer_1[546] = ~layer_0[554]; 
    assign layer_1[547] = layer_0[541] | layer_0[556]; 
    assign layer_1[548] = ~(layer_0[554] & layer_0[554]); 
    assign layer_1[549] = ~(layer_0[553] | layer_0[562]); 
    assign layer_1[550] = 1'b1; 
    assign layer_1[551] = layer_0[547]; 
    assign layer_1[552] = layer_0[546] & ~layer_0[563]; 
    assign layer_1[553] = ~layer_0[561]; 
    assign layer_1[554] = layer_0[539] & ~layer_0[558]; 
    assign layer_1[555] = ~layer_0[564] | (layer_0[569] & layer_0[564]); 
    assign layer_1[556] = layer_0[557] | layer_0[546]; 
    assign layer_1[557] = layer_0[561]; 
    assign layer_1[558] = ~layer_0[541]; 
    assign layer_1[559] = ~layer_0[547]; 
    assign layer_1[560] = layer_0[576] | layer_0[556]; 
    assign layer_1[561] = layer_0[546]; 
    assign layer_1[562] = ~layer_0[553]; 
    assign layer_1[563] = layer_0[567]; 
    assign layer_1[564] = ~layer_0[560] | (layer_0[578] & layer_0[560]); 
    assign layer_1[565] = layer_0[550] & ~layer_0[571]; 
    assign layer_1[566] = 1'b0; 
    assign layer_1[567] = layer_0[566] & ~layer_0[556]; 
    assign layer_1[568] = layer_0[574] & layer_0[567]; 
    assign layer_1[569] = ~(layer_0[579] & layer_0[552]); 
    assign layer_1[570] = ~layer_0[575]; 
    assign layer_1[571] = layer_0[569] | layer_0[579]; 
    assign layer_1[572] = ~(layer_0[562] | layer_0[578]); 
    assign layer_1[573] = ~layer_0[575]; 
    assign layer_1[574] = ~(layer_0[570] & layer_0[579]); 
    assign layer_1[575] = ~layer_0[564] | (layer_0[564] & layer_0[584]); 
    assign layer_1[576] = 1'b1; 
    assign layer_1[577] = ~(layer_0[580] | layer_0[562]); 
    assign layer_1[578] = 1'b0; 
    assign layer_1[579] = layer_0[581] | layer_0[568]; 
    assign layer_1[580] = layer_0[584] | layer_0[591]; 
    assign layer_1[581] = layer_0[580] & layer_0[580]; 
    assign layer_1[582] = ~layer_0[565] | (layer_0[597] & layer_0[565]); 
    assign layer_1[583] = ~layer_0[589]; 
    assign layer_1[584] = layer_0[595]; 
    assign layer_1[585] = ~(layer_0[572] ^ layer_0[588]); 
    assign layer_1[586] = layer_0[599] | layer_0[569]; 
    assign layer_1[587] = ~(layer_0[591] | layer_0[578]); 
    assign layer_1[588] = ~(layer_0[595] | layer_0[581]); 
    assign layer_1[589] = layer_0[587] | layer_0[589]; 
    assign layer_1[590] = ~layer_0[597] | (layer_0[578] & layer_0[597]); 
    assign layer_1[591] = ~layer_0[579]; 
    assign layer_1[592] = 1'b0; 
    assign layer_1[593] = layer_0[581]; 
    assign layer_1[594] = layer_0[595] | layer_0[580]; 
    assign layer_1[595] = layer_0[605] | layer_0[580]; 
    assign layer_1[596] = layer_0[586] ^ layer_0[606]; 
    assign layer_1[597] = ~(layer_0[591] & layer_0[584]); 
    assign layer_1[598] = ~(layer_0[594] ^ layer_0[595]); 
    assign layer_1[599] = ~layer_0[601]; 
    assign layer_1[600] = layer_0[610]; 
    assign layer_1[601] = layer_0[610] & layer_0[587]; 
    assign layer_1[602] = ~(layer_0[589] & layer_0[597]); 
    assign layer_1[603] = layer_0[619] & ~layer_0[586]; 
    assign layer_1[604] = ~(layer_0[618] | layer_0[609]); 
    assign layer_1[605] = ~layer_0[608] | (layer_0[607] & layer_0[608]); 
    assign layer_1[606] = ~layer_0[589]; 
    assign layer_1[607] = layer_0[602] | layer_0[616]; 
    assign layer_1[608] = ~(layer_0[619] | layer_0[607]); 
    assign layer_1[609] = ~(layer_0[605] | layer_0[607]); 
    assign layer_1[610] = ~layer_0[622] | (layer_0[622] & layer_0[611]); 
    assign layer_1[611] = 1'b0; 
    assign layer_1[612] = 1'b0; 
    assign layer_1[613] = 1'b1; 
    assign layer_1[614] = layer_0[598] & ~layer_0[612]; 
    assign layer_1[615] = layer_0[601]; 
    assign layer_1[616] = ~layer_0[624] | (layer_0[622] & layer_0[624]); 
    assign layer_1[617] = layer_0[632]; 
    assign layer_1[618] = layer_0[621] & ~layer_0[617]; 
    assign layer_1[619] = ~layer_0[605] | (layer_0[625] & layer_0[605]); 
    assign layer_1[620] = ~(layer_0[630] | layer_0[622]); 
    assign layer_1[621] = ~layer_0[617] | (layer_0[619] & layer_0[617]); 
    assign layer_1[622] = ~(layer_0[607] & layer_0[622]); 
    assign layer_1[623] = ~layer_0[619]; 
    assign layer_1[624] = layer_0[618]; 
    assign layer_1[625] = ~layer_0[611] | (layer_0[617] & layer_0[611]); 
    assign layer_1[626] = layer_0[638] & layer_0[638]; 
    assign layer_1[627] = layer_0[623]; 
    assign layer_1[628] = ~(layer_0[623] | layer_0[627]); 
    assign layer_1[629] = layer_0[618] | layer_0[618]; 
    assign layer_1[630] = 1'b0; 
    assign layer_1[631] = ~layer_0[643] | (layer_0[643] & layer_0[644]); 
    assign layer_1[632] = ~(layer_0[616] | layer_0[641]); 
    assign layer_1[633] = layer_0[639] | layer_0[621]; 
    assign layer_1[634] = layer_0[632] ^ layer_0[618]; 
    assign layer_1[635] = layer_0[624] & ~layer_0[630]; 
    assign layer_1[636] = ~(layer_0[628] | layer_0[640]); 
    assign layer_1[637] = layer_0[648]; 
    assign layer_1[638] = layer_0[638]; 
    assign layer_1[639] = ~layer_0[636]; 
    assign layer_1[640] = ~layer_0[626]; 
    assign layer_1[641] = layer_0[650] & ~layer_0[653]; 
    assign layer_1[642] = ~(layer_0[644] & layer_0[646]); 
    assign layer_1[643] = layer_0[643]; 
    assign layer_1[644] = ~layer_0[651]; 
    assign layer_1[645] = ~layer_0[645] | (layer_0[657] & layer_0[645]); 
    assign layer_1[646] = layer_0[647] & ~layer_0[633]; 
    assign layer_1[647] = layer_0[635] & layer_0[653]; 
    assign layer_1[648] = layer_0[649] & layer_0[663]; 
    assign layer_1[649] = layer_0[646]; 
    assign layer_1[650] = 1'b0; 
    assign layer_1[651] = ~(layer_0[636] ^ layer_0[640]); 
    assign layer_1[652] = ~layer_0[640] | (layer_0[640] & layer_0[640]); 
    assign layer_1[653] = layer_0[653] | layer_0[649]; 
    assign layer_1[654] = ~layer_0[663] | (layer_0[663] & layer_0[638]); 
    assign layer_1[655] = layer_0[671]; 
    assign layer_1[656] = layer_0[668] | layer_0[663]; 
    assign layer_1[657] = 1'b1; 
    assign layer_1[658] = ~(layer_0[658] | layer_0[659]); 
    assign layer_1[659] = 1'b0; 
    assign layer_1[660] = layer_0[662]; 
    assign layer_1[661] = ~(layer_0[647] & layer_0[676]); 
    assign layer_1[662] = ~(layer_0[649] & layer_0[660]); 
    assign layer_1[663] = layer_0[676] ^ layer_0[665]; 
    assign layer_1[664] = ~(layer_0[673] | layer_0[670]); 
    assign layer_1[665] = layer_0[659]; 
    assign layer_1[666] = layer_0[679] | layer_0[680]; 
    assign layer_1[667] = 1'b1; 
    assign layer_1[668] = layer_0[673] & layer_0[654]; 
    assign layer_1[669] = layer_0[664] ^ layer_0[657]; 
    assign layer_1[670] = ~layer_0[685]; 
    assign layer_1[671] = 1'b1; 
    assign layer_1[672] = 1'b0; 
    assign layer_1[673] = ~layer_0[689] | (layer_0[689] & layer_0[680]); 
    assign layer_1[674] = ~layer_0[684] | (layer_0[684] & layer_0[676]); 
    assign layer_1[675] = ~(layer_0[671] | layer_0[667]); 
    assign layer_1[676] = ~layer_0[671] | (layer_0[671] & layer_0[677]); 
    assign layer_1[677] = ~layer_0[682]; 
    assign layer_1[678] = ~(layer_0[682] | layer_0[667]); 
    assign layer_1[679] = ~(layer_0[679] & layer_0[691]); 
    assign layer_1[680] = layer_0[685] ^ layer_0[692]; 
    assign layer_1[681] = layer_0[666] & ~layer_0[690]; 
    assign layer_1[682] = ~(layer_0[673] ^ layer_0[694]); 
    assign layer_1[683] = 1'b0; 
    assign layer_1[684] = layer_0[691]; 
    assign layer_1[685] = ~layer_0[677] | (layer_0[677] & layer_0[671]); 
    assign layer_1[686] = ~(layer_0[702] | layer_0[676]); 
    assign layer_1[687] = ~(layer_0[698] & layer_0[692]); 
    assign layer_1[688] = ~layer_0[685] | (layer_0[700] & layer_0[685]); 
    assign layer_1[689] = ~(layer_0[688] | layer_0[687]); 
    assign layer_1[690] = ~layer_0[697]; 
    assign layer_1[691] = layer_0[701] & ~layer_0[688]; 
    assign layer_1[692] = ~layer_0[706]; 
    assign layer_1[693] = ~layer_0[695] | (layer_0[695] & layer_0[683]); 
    assign layer_1[694] = layer_0[681] ^ layer_0[686]; 
    assign layer_1[695] = ~(layer_0[702] | layer_0[700]); 
    assign layer_1[696] = 1'b1; 
    assign layer_1[697] = layer_0[680] & ~layer_0[700]; 
    assign layer_1[698] = layer_0[701] ^ layer_0[689]; 
    assign layer_1[699] = ~layer_0[692] | (layer_0[692] & layer_0[700]); 
    assign layer_1[700] = layer_0[699]; 
    assign layer_1[701] = ~layer_0[704]; 
    assign layer_1[702] = ~layer_0[707]; 
    assign layer_1[703] = layer_0[701] ^ layer_0[709]; 
    assign layer_1[704] = layer_0[702] & layer_0[702]; 
    assign layer_1[705] = 1'b1; 
    assign layer_1[706] = layer_0[692]; 
    assign layer_1[707] = 1'b1; 
    assign layer_1[708] = layer_0[717] & layer_0[716]; 
    assign layer_1[709] = ~layer_0[695] | (layer_0[695] & layer_0[705]); 
    assign layer_1[710] = ~(layer_0[712] ^ layer_0[718]); 
    assign layer_1[711] = ~(layer_0[708] | layer_0[703]); 
    assign layer_1[712] = 1'b1; 
    assign layer_1[713] = ~layer_0[706] | (layer_0[706] & layer_0[696]); 
    assign layer_1[714] = ~(layer_0[700] & layer_0[699]); 
    assign layer_1[715] = layer_0[704] & layer_0[699]; 
    assign layer_1[716] = layer_0[706]; 
    assign layer_1[717] = 1'b0; 
    assign layer_1[718] = layer_0[728] & ~layer_0[729]; 
    assign layer_1[719] = layer_0[728] & layer_0[733]; 
    assign layer_1[720] = ~layer_0[724] | (layer_0[715] & layer_0[724]); 
    assign layer_1[721] = layer_0[726] & ~layer_0[707]; 
    assign layer_1[722] = layer_0[715]; 
    assign layer_1[723] = layer_0[707] & ~layer_0[723]; 
    assign layer_1[724] = 1'b1; 
    assign layer_1[725] = layer_0[731] | layer_0[722]; 
    assign layer_1[726] = ~layer_0[719]; 
    assign layer_1[727] = 1'b0; 
    assign layer_1[728] = layer_0[718]; 
    assign layer_1[729] = layer_0[741] & ~layer_0[741]; 
    assign layer_1[730] = layer_0[716] ^ layer_0[732]; 
    assign layer_1[731] = 1'b1; 
    assign layer_1[732] = 1'b0; 
    assign layer_1[733] = 1'b1; 
    assign layer_1[734] = ~layer_0[719] | (layer_0[722] & layer_0[719]); 
    assign layer_1[735] = ~layer_0[728]; 
    assign layer_1[736] = layer_0[724] & layer_0[749]; 
    assign layer_1[737] = ~layer_0[734] | (layer_0[744] & layer_0[734]); 
    assign layer_1[738] = ~(layer_0[732] ^ layer_0[723]); 
    assign layer_1[739] = 1'b1; 
    assign layer_1[740] = ~(layer_0[750] | layer_0[734]); 
    assign layer_1[741] = layer_0[754] & layer_0[739]; 
    assign layer_1[742] = layer_0[738]; 
    assign layer_1[743] = ~(layer_0[727] ^ layer_0[739]); 
    assign layer_1[744] = ~(layer_0[731] | layer_0[740]); 
    assign layer_1[745] = ~layer_0[753]; 
    assign layer_1[746] = ~layer_0[758] | (layer_0[755] & layer_0[758]); 
    assign layer_1[747] = layer_0[743] & ~layer_0[742]; 
    assign layer_1[748] = layer_0[743] & ~layer_0[741]; 
    assign layer_1[749] = ~(layer_0[743] & layer_0[749]); 
    assign layer_1[750] = ~layer_0[734]; 
    assign layer_1[751] = ~layer_0[741] | (layer_0[741] & layer_0[749]); 
    assign layer_1[752] = layer_0[760] & layer_0[748]; 
    assign layer_1[753] = layer_0[745] ^ layer_0[736]; 
    assign layer_1[754] = layer_0[751] & ~layer_0[758]; 
    assign layer_1[755] = layer_0[747]; 
    assign layer_1[756] = 1'b0; 
    assign layer_1[757] = 1'b0; 
    assign layer_1[758] = layer_0[742] ^ layer_0[743]; 
    assign layer_1[759] = ~(layer_0[764] ^ layer_0[760]); 
    assign layer_1[760] = ~(layer_0[759] | layer_0[770]); 
    assign layer_1[761] = ~layer_0[750]; 
    assign layer_1[762] = layer_0[756] ^ layer_0[763]; 
    assign layer_1[763] = layer_0[760]; 
    assign layer_1[764] = ~layer_0[753] | (layer_0[764] & layer_0[753]); 
    assign layer_1[765] = ~layer_0[767] | (layer_0[766] & layer_0[767]); 
    assign layer_1[766] = layer_0[759] & ~layer_0[769]; 
    assign layer_1[767] = layer_0[779] & ~layer_0[758]; 
    assign layer_1[768] = layer_0[764] & ~layer_0[759]; 
    assign layer_1[769] = ~layer_0[761] | (layer_0[773] & layer_0[761]); 
    assign layer_1[770] = ~layer_0[771]; 
    assign layer_1[771] = 1'b1; 
    assign layer_1[772] = layer_0[766] & layer_0[785]; 
    assign layer_1[773] = layer_0[776] | layer_0[757]; 
    assign layer_1[774] = 1'b1; 
    assign layer_1[775] = ~(layer_0[778] ^ layer_0[786]); 
    assign layer_1[776] = layer_0[765] | layer_0[759]; 
    assign layer_1[777] = ~(layer_0[776] | layer_0[764]); 
    assign layer_1[778] = ~layer_0[791]; 
    assign layer_1[779] = layer_0[770] & ~layer_0[777]; 
    assign layer_1[780] = 1'b1; 
    assign layer_1[781] = layer_0[788] | layer_0[790]; 
    assign layer_1[782] = ~(layer_0[792] | layer_0[792]); 
    assign layer_1[783] = ~layer_0[794] | (layer_0[794] & layer_0[775]); 
    assign layer_1[784] = 1'b0; 
    assign layer_1[785] = ~layer_0[788] | (layer_0[770] & layer_0[788]); 
    assign layer_1[786] = layer_0[792] & layer_0[794]; 
    assign layer_1[787] = layer_0[775] & layer_0[792]; 
    assign layer_1[788] = ~layer_0[772] | (layer_0[773] & layer_0[772]); 
    assign layer_1[789] = layer_0[792] | layer_0[797]; 
    assign layer_1[790] = 1'b1; 
    assign layer_1[791] = layer_0[806] & ~layer_0[790]; 
    assign layer_1[792] = layer_0[807] ^ layer_0[799]; 
    assign layer_1[793] = ~layer_0[796]; 
    assign layer_1[794] = layer_0[801] ^ layer_0[778]; 
    assign layer_1[795] = ~(layer_0[779] & layer_0[809]); 
    assign layer_1[796] = ~layer_0[789]; 
    assign layer_1[797] = ~(layer_0[788] & layer_0[801]); 
    assign layer_1[798] = ~layer_0[785]; 
    assign layer_1[799] = layer_0[787] ^ layer_0[802]; 
    assign layer_1[800] = ~layer_0[788] | (layer_0[792] & layer_0[788]); 
    assign layer_1[801] = layer_0[811] & layer_0[784]; 
    assign layer_1[802] = layer_0[796] ^ layer_0[799]; 
    assign layer_1[803] = layer_0[791] | layer_0[811]; 
    assign layer_1[804] = layer_0[817] & ~layer_0[798]; 
    assign layer_1[805] = layer_0[819] | layer_0[806]; 
    assign layer_1[806] = layer_0[807] & ~layer_0[796]; 
    assign layer_1[807] = 1'b1; 
    assign layer_1[808] = layer_0[811] | layer_0[817]; 
    assign layer_1[809] = layer_0[808] & ~layer_0[814]; 
    assign layer_1[810] = ~layer_0[794]; 
    assign layer_1[811] = layer_0[819] & layer_0[819]; 
    assign layer_1[812] = layer_0[798] | layer_0[823]; 
    assign layer_1[813] = layer_0[814]; 
    assign layer_1[814] = layer_0[812] & ~layer_0[816]; 
    assign layer_1[815] = layer_0[800]; 
    assign layer_1[816] = layer_0[831] & ~layer_0[819]; 
    assign layer_1[817] = ~layer_0[804] | (layer_0[804] & layer_0[829]); 
    assign layer_1[818] = ~(layer_0[833] & layer_0[833]); 
    assign layer_1[819] = ~(layer_0[808] | layer_0[824]); 
    assign layer_1[820] = 1'b1; 
    assign layer_1[821] = 1'b0; 
    assign layer_1[822] = layer_0[806] | layer_0[811]; 
    assign layer_1[823] = ~(layer_0[807] ^ layer_0[828]); 
    assign layer_1[824] = layer_0[832] & ~layer_0[822]; 
    assign layer_1[825] = ~layer_0[813] | (layer_0[835] & layer_0[813]); 
    assign layer_1[826] = layer_0[831] ^ layer_0[827]; 
    assign layer_1[827] = ~(layer_0[823] & layer_0[842]); 
    assign layer_1[828] = layer_0[825] | layer_0[840]; 
    assign layer_1[829] = layer_0[821] & layer_0[816]; 
    assign layer_1[830] = layer_0[827]; 
    assign layer_1[831] = layer_0[826] & ~layer_0[837]; 
    assign layer_1[832] = ~layer_0[842]; 
    assign layer_1[833] = layer_0[819] | layer_0[833]; 
    assign layer_1[834] = layer_0[835] & ~layer_0[819]; 
    assign layer_1[835] = ~(layer_0[847] & layer_0[821]); 
    assign layer_1[836] = layer_0[844]; 
    assign layer_1[837] = ~layer_0[842] | (layer_0[853] & layer_0[842]); 
    assign layer_1[838] = 1'b1; 
    assign layer_1[839] = 1'b1; 
    assign layer_1[840] = ~(layer_0[829] & layer_0[854]); 
    assign layer_1[841] = layer_0[844] & ~layer_0[843]; 
    assign layer_1[842] = ~layer_0[856] | (layer_0[856] & layer_0[825]); 
    assign layer_1[843] = ~layer_0[841] | (layer_0[841] & layer_0[856]); 
    assign layer_1[844] = ~(layer_0[829] ^ layer_0[833]); 
    assign layer_1[845] = 1'b1; 
    assign layer_1[846] = 1'b0; 
    assign layer_1[847] = layer_0[849]; 
    assign layer_1[848] = layer_0[852]; 
    assign layer_1[849] = layer_0[852] ^ layer_0[832]; 
    assign layer_1[850] = layer_0[848]; 
    assign layer_1[851] = 1'b0; 
    assign layer_1[852] = ~(layer_0[856] | layer_0[865]); 
    assign layer_1[853] = layer_0[862]; 
    assign layer_1[854] = layer_0[846]; 
    assign layer_1[855] = layer_0[840] ^ layer_0[866]; 
    assign layer_1[856] = 1'b1; 
    assign layer_1[857] = ~(layer_0[861] | layer_0[857]); 
    assign layer_1[858] = layer_0[855]; 
    assign layer_1[859] = layer_0[861]; 
    assign layer_1[860] = ~(layer_0[872] & layer_0[866]); 
    assign layer_1[861] = ~layer_0[876]; 
    assign layer_1[862] = layer_0[855] & ~layer_0[869]; 
    assign layer_1[863] = ~layer_0[878] | (layer_0[869] & layer_0[878]); 
    assign layer_1[864] = layer_0[853] & ~layer_0[864]; 
    assign layer_1[865] = ~layer_0[855]; 
    assign layer_1[866] = ~layer_0[873] | (layer_0[873] & layer_0[858]); 
    assign layer_1[867] = layer_0[871] ^ layer_0[863]; 
    assign layer_1[868] = ~layer_0[855] | (layer_0[878] & layer_0[855]); 
    assign layer_1[869] = layer_0[879]; 
    assign layer_1[870] = layer_0[878]; 
    assign layer_1[871] = layer_0[862] & layer_0[886]; 
    assign layer_1[872] = ~layer_0[862] | (layer_0[877] & layer_0[862]); 
    assign layer_1[873] = ~(layer_0[867] & layer_0[875]); 
    assign layer_1[874] = layer_0[876] | layer_0[870]; 
    assign layer_1[875] = 1'b0; 
    assign layer_1[876] = layer_0[873] & layer_0[870]; 
    assign layer_1[877] = layer_0[889] & ~layer_0[860]; 
    assign layer_1[878] = ~layer_0[892] | (layer_0[892] & layer_0[891]); 
    assign layer_1[879] = 1'b1; 
    assign layer_1[880] = layer_0[896] ^ layer_0[887]; 
    assign layer_1[881] = layer_0[897] & ~layer_0[893]; 
    assign layer_1[882] = layer_0[888] & ~layer_0[895]; 
    assign layer_1[883] = ~(layer_0[873] & layer_0[881]); 
    assign layer_1[884] = layer_0[898] & ~layer_0[888]; 
    assign layer_1[885] = ~layer_0[887] | (layer_0[887] & layer_0[870]); 
    assign layer_1[886] = layer_0[870] & ~layer_0[878]; 
    assign layer_1[887] = ~(layer_0[875] ^ layer_0[871]); 
    assign layer_1[888] = ~(layer_0[886] | layer_0[889]); 
    assign layer_1[889] = layer_0[874] & ~layer_0[877]; 
    assign layer_1[890] = ~layer_0[878]; 
    assign layer_1[891] = layer_0[887]; 
    assign layer_1[892] = layer_0[878]; 
    assign layer_1[893] = layer_0[882] & ~layer_0[881]; 
    assign layer_1[894] = layer_0[909] & layer_0[894]; 
    assign layer_1[895] = 1'b1; 
    assign layer_1[896] = ~layer_0[882]; 
    assign layer_1[897] = ~layer_0[893]; 
    assign layer_1[898] = layer_0[887] & layer_0[894]; 
    assign layer_1[899] = layer_0[897] & ~layer_0[893]; 
    assign layer_1[900] = layer_0[888] | layer_0[897]; 
    assign layer_1[901] = ~layer_0[896] | (layer_0[890] & layer_0[896]); 
    assign layer_1[902] = layer_0[909] & layer_0[887]; 
    assign layer_1[903] = ~layer_0[918] | (layer_0[901] & layer_0[918]); 
    assign layer_1[904] = layer_0[915] & ~layer_0[919]; 
    assign layer_1[905] = layer_0[919] & ~layer_0[897]; 
    assign layer_1[906] = layer_0[911] & layer_0[912]; 
    assign layer_1[907] = ~layer_0[891] | (layer_0[910] & layer_0[891]); 
    assign layer_1[908] = ~(layer_0[910] & layer_0[919]); 
    assign layer_1[909] = layer_0[910] & ~layer_0[903]; 
    assign layer_1[910] = ~(layer_0[897] | layer_0[914]); 
    assign layer_1[911] = layer_0[913]; 
    assign layer_1[912] = ~(layer_0[926] | layer_0[897]); 
    assign layer_1[913] = layer_0[929] & layer_0[914]; 
    assign layer_1[914] = layer_0[922]; 
    assign layer_1[915] = ~layer_0[920]; 
    assign layer_1[916] = ~layer_0[910] | (layer_0[910] & layer_0[919]); 
    assign layer_1[917] = ~layer_0[926]; 
    assign layer_1[918] = layer_0[929]; 
    assign layer_1[919] = layer_0[905] & layer_0[905]; 
    assign layer_1[920] = layer_0[917] ^ layer_0[927]; 
    assign layer_1[921] = layer_0[920] | layer_0[912]; 
    assign layer_1[922] = layer_0[925] & layer_0[933]; 
    assign layer_1[923] = layer_0[928] & ~layer_0[923]; 
    assign layer_1[924] = ~layer_0[939] | (layer_0[915] & layer_0[939]); 
    assign layer_1[925] = layer_0[933]; 
    assign layer_1[926] = ~layer_0[918]; 
    assign layer_1[927] = layer_0[937] | layer_0[938]; 
    assign layer_1[928] = ~layer_0[932] | (layer_0[932] & layer_0[942]); 
    assign layer_1[929] = layer_0[930] & ~layer_0[924]; 
    assign layer_1[930] = layer_0[916] | layer_0[927]; 
    assign layer_1[931] = layer_0[947] & layer_0[935]; 
    assign layer_1[932] = ~(layer_0[916] | layer_0[934]); 
    assign layer_1[933] = ~(layer_0[933] | layer_0[945]); 
    assign layer_1[934] = ~layer_0[921]; 
    assign layer_1[935] = layer_0[949] | layer_0[945]; 
    assign layer_1[936] = ~layer_0[924] | (layer_0[924] & layer_0[929]); 
    assign layer_1[937] = layer_0[937]; 
    assign layer_1[938] = ~(layer_0[923] ^ layer_0[940]); 
    assign layer_1[939] = ~(layer_0[929] | layer_0[927]); 
    assign layer_1[940] = 1'b1; 
    assign layer_1[941] = ~(layer_0[930] ^ layer_0[934]); 
    assign layer_1[942] = ~(layer_0[939] ^ layer_0[934]); 
    assign layer_1[943] = layer_0[939] & ~layer_0[941]; 
    assign layer_1[944] = 1'b0; 
    assign layer_1[945] = layer_0[934] ^ layer_0[939]; 
    assign layer_1[946] = 1'b0; 
    assign layer_1[947] = ~layer_0[933] | (layer_0[933] & layer_0[937]); 
    assign layer_1[948] = ~(layer_0[940] | layer_0[955]); 
    assign layer_1[949] = layer_0[964]; 
    assign layer_1[950] = layer_0[964] & ~layer_0[955]; 
    assign layer_1[951] = layer_0[950] & ~layer_0[943]; 
    assign layer_1[952] = ~(layer_0[952] & layer_0[962]); 
    assign layer_1[953] = ~layer_0[940]; 
    assign layer_1[954] = ~layer_0[940]; 
    assign layer_1[955] = layer_0[970] ^ layer_0[966]; 
    assign layer_1[956] = ~(layer_0[943] & layer_0[947]); 
    assign layer_1[957] = layer_0[972] & ~layer_0[963]; 
    assign layer_1[958] = ~layer_0[946] | (layer_0[946] & layer_0[941]); 
    assign layer_1[959] = layer_0[961] & layer_0[971]; 
    assign layer_1[960] = layer_0[950] ^ layer_0[971]; 
    assign layer_1[961] = ~layer_0[947] | (layer_0[960] & layer_0[947]); 
    assign layer_1[962] = layer_0[970]; 
    assign layer_1[963] = 1'b0; 
    assign layer_1[964] = layer_0[958] ^ layer_0[953]; 
    assign layer_1[965] = 1'b0; 
    assign layer_1[966] = layer_0[965] & ~layer_0[954]; 
    assign layer_1[967] = layer_0[977] & layer_0[954]; 
    assign layer_1[968] = ~layer_0[965]; 
    assign layer_1[969] = layer_0[955] ^ layer_0[975]; 
    assign layer_1[970] = layer_0[973]; 
    assign layer_1[971] = layer_0[984] & ~layer_0[956]; 
    assign layer_1[972] = ~(layer_0[970] ^ layer_0[969]); 
    assign layer_1[973] = layer_0[971] & layer_0[975]; 
    assign layer_1[974] = layer_0[975] ^ layer_0[983]; 
    assign layer_1[975] = ~(layer_0[971] | layer_0[971]); 
    assign layer_1[976] = layer_0[970] ^ layer_0[973]; 
    assign layer_1[977] = ~layer_0[972]; 
    assign layer_1[978] = ~(layer_0[970] ^ layer_0[988]); 
    assign layer_1[979] = ~layer_0[967] | (layer_0[984] & layer_0[967]); 
    assign layer_1[980] = layer_0[980] & ~layer_0[975]; 
    assign layer_1[981] = layer_0[992]; 
    assign layer_1[982] = layer_0[966] & layer_0[977]; 
    assign layer_1[983] = 1'b0; 
    assign layer_1[984] = layer_0[992] & layer_0[998]; 
    assign layer_1[985] = ~(layer_0[986] & layer_0[993]); 
    assign layer_1[986] = layer_0[989] & ~layer_0[992]; 
    assign layer_1[987] = ~layer_0[978] | (layer_0[978] & layer_0[987]); 
    assign layer_1[988] = layer_0[991] | layer_0[985]; 
    assign layer_1[989] = ~layer_0[1002]; 
    assign layer_1[990] = layer_0[978]; 
    assign layer_1[991] = ~layer_0[987]; 
    assign layer_1[992] = 1'b1; 
    assign layer_1[993] = layer_0[1005] & layer_0[993]; 
    assign layer_1[994] = 1'b1; 
    assign layer_1[995] = ~layer_0[990]; 
    assign layer_1[996] = 1'b1; 
    assign layer_1[997] = ~(layer_0[996] | layer_0[981]); 
    assign layer_1[998] = 1'b0; 
    assign layer_1[999] = 1'b1; 
    assign layer_1[1000] = layer_0[1014] & ~layer_0[1015]; 
    assign layer_1[1001] = layer_0[1015]; 
    assign layer_1[1002] = layer_0[997] & ~layer_0[997]; 
    assign layer_1[1003] = ~(layer_0[1013] | layer_0[997]); 
    assign layer_1[1004] = layer_0[998] & ~layer_0[993]; 
    assign layer_1[1005] = layer_0[1010] & ~layer_0[1005]; 
    assign layer_1[1006] = ~(layer_0[990] | layer_0[1008]); 
    assign layer_1[1007] = layer_0[1007] ^ layer_0[1016]; 
    assign layer_1[1008] = layer_0[992] & layer_0[999]; 
    assign layer_1[1009] = layer_0[1002] & layer_0[1011]; 
    assign layer_1[1010] = 1'b0; 
    assign layer_1[1011] = layer_0[1014] & ~layer_0[1014]; 
    assign layer_1[1012] = ~layer_0[1014]; 
    assign layer_1[1013] = layer_0[1018] & ~layer_0[1013]; 
    assign layer_1[1014] = layer_0[1000]; 
    assign layer_1[1015] = layer_0[1005] & ~layer_0[1019]; 
    assign layer_1[1016] = ~layer_0[999] | (layer_0[1019] & layer_0[999]); 
    assign layer_1[1017] = layer_0[1019]; 
    assign layer_1[1018] = 1'b1; 
    assign layer_1[1019] = layer_0[1013] & ~layer_0[1017]; 
    assign layer_1[1020] = ~layer_0[1018]; 
    assign layer_1[1021] = ~(layer_0[1014] & layer_0[1011]); 
    assign layer_1[1022] = layer_0[1021]; 
    assign layer_1[1023] = ~(layer_0[1013] | layer_0[1023]); 
    // Layer 2 ============================================================
    assign layer_2[0] = ~(layer_1[12] ^ layer_1[1]); 
    assign layer_2[1] = 1'b1; 
    assign layer_2[2] = ~layer_1[4]; 
    assign layer_2[3] = layer_1[13] & ~layer_1[12]; 
    assign layer_2[4] = layer_1[11]; 
    assign layer_2[5] = 1'b1; 
    assign layer_2[6] = ~layer_1[4] | (layer_1[4] & layer_1[3]); 
    assign layer_2[7] = layer_1[12] | layer_1[5]; 
    assign layer_2[8] = layer_1[3] & ~layer_1[22]; 
    assign layer_2[9] = ~(layer_1[2] & layer_1[0]); 
    assign layer_2[10] = ~(layer_1[10] | layer_1[7]); 
    assign layer_2[11] = layer_1[18] | layer_1[20]; 
    assign layer_2[12] = ~layer_1[16] | (layer_1[16] & layer_1[5]); 
    assign layer_2[13] = layer_1[3]; 
    assign layer_2[14] = layer_1[15]; 
    assign layer_2[15] = layer_1[11] ^ layer_1[21]; 
    assign layer_2[16] = ~(layer_1[6] ^ layer_1[22]); 
    assign layer_2[17] = ~layer_1[27] | (layer_1[23] & layer_1[27]); 
    assign layer_2[18] = layer_1[11] | layer_1[28]; 
    assign layer_2[19] = layer_1[14]; 
    assign layer_2[20] = ~layer_1[17] | (layer_1[17] & layer_1[12]); 
    assign layer_2[21] = layer_1[17] ^ layer_1[19]; 
    assign layer_2[22] = ~layer_1[36]; 
    assign layer_2[23] = layer_1[10] | layer_1[14]; 
    assign layer_2[24] = ~layer_1[11] | (layer_1[11] & layer_1[36]); 
    assign layer_2[25] = ~layer_1[37]; 
    assign layer_2[26] = layer_1[37] ^ layer_1[22]; 
    assign layer_2[27] = layer_1[20] & ~layer_1[14]; 
    assign layer_2[28] = layer_1[14] ^ layer_1[24]; 
    assign layer_2[29] = layer_1[19] | layer_1[32]; 
    assign layer_2[30] = layer_1[24] & ~layer_1[17]; 
    assign layer_2[31] = ~(layer_1[31] | layer_1[37]); 
    assign layer_2[32] = layer_1[46] & ~layer_1[18]; 
    assign layer_2[33] = ~(layer_1[37] | layer_1[41]); 
    assign layer_2[34] = ~(layer_1[41] & layer_1[48]); 
    assign layer_2[35] = 1'b1; 
    assign layer_2[36] = ~layer_1[52] | (layer_1[52] & layer_1[26]); 
    assign layer_2[37] = ~layer_1[52]; 
    assign layer_2[38] = layer_1[43] & layer_1[31]; 
    assign layer_2[39] = ~(layer_1[55] & layer_1[46]); 
    assign layer_2[40] = layer_1[47] & ~layer_1[31]; 
    assign layer_2[41] = ~(layer_1[30] & layer_1[48]); 
    assign layer_2[42] = ~layer_1[33] | (layer_1[33] & layer_1[49]); 
    assign layer_2[43] = ~(layer_1[43] & layer_1[35]); 
    assign layer_2[44] = 1'b1; 
    assign layer_2[45] = layer_1[52]; 
    assign layer_2[46] = ~layer_1[51]; 
    assign layer_2[47] = layer_1[53] & ~layer_1[37]; 
    assign layer_2[48] = ~layer_1[41]; 
    assign layer_2[49] = layer_1[58] ^ layer_1[56]; 
    assign layer_2[50] = 1'b1; 
    assign layer_2[51] = 1'b0; 
    assign layer_2[52] = ~(layer_1[50] ^ layer_1[42]); 
    assign layer_2[53] = ~(layer_1[46] ^ layer_1[38]); 
    assign layer_2[54] = ~(layer_1[70] & layer_1[43]); 
    assign layer_2[55] = ~(layer_1[58] & layer_1[61]); 
    assign layer_2[56] = ~layer_1[65]; 
    assign layer_2[57] = ~layer_1[72] | (layer_1[72] & layer_1[63]); 
    assign layer_2[58] = layer_1[43] | layer_1[70]; 
    assign layer_2[59] = ~layer_1[63]; 
    assign layer_2[60] = layer_1[71] ^ layer_1[74]; 
    assign layer_2[61] = layer_1[72]; 
    assign layer_2[62] = ~(layer_1[63] | layer_1[58]); 
    assign layer_2[63] = layer_1[73] & ~layer_1[63]; 
    assign layer_2[64] = layer_1[49] ^ layer_1[50]; 
    assign layer_2[65] = ~layer_1[70] | (layer_1[70] & layer_1[56]); 
    assign layer_2[66] = layer_1[75] & ~layer_1[71]; 
    assign layer_2[67] = ~layer_1[59] | (layer_1[68] & layer_1[59]); 
    assign layer_2[68] = layer_1[56] ^ layer_1[59]; 
    assign layer_2[69] = layer_1[59] ^ layer_1[71]; 
    assign layer_2[70] = 1'b0; 
    assign layer_2[71] = ~layer_1[73]; 
    assign layer_2[72] = ~(layer_1[61] & layer_1[85]); 
    assign layer_2[73] = ~(layer_1[65] | layer_1[56]); 
    assign layer_2[74] = ~(layer_1[90] & layer_1[80]); 
    assign layer_2[75] = ~(layer_1[73] & layer_1[75]); 
    assign layer_2[76] = ~layer_1[72] | (layer_1[82] & layer_1[72]); 
    assign layer_2[77] = ~layer_1[69]; 
    assign layer_2[78] = ~layer_1[62] | (layer_1[76] & layer_1[62]); 
    assign layer_2[79] = ~(layer_1[66] ^ layer_1[91]); 
    assign layer_2[80] = layer_1[92] & ~layer_1[91]; 
    assign layer_2[81] = ~layer_1[81] | (layer_1[88] & layer_1[81]); 
    assign layer_2[82] = ~layer_1[69] | (layer_1[69] & layer_1[84]); 
    assign layer_2[83] = ~layer_1[95]; 
    assign layer_2[84] = layer_1[100] ^ layer_1[71]; 
    assign layer_2[85] = 1'b1; 
    assign layer_2[86] = ~layer_1[75] | (layer_1[75] & layer_1[101]); 
    assign layer_2[87] = layer_1[103] ^ layer_1[77]; 
    assign layer_2[88] = ~layer_1[86]; 
    assign layer_2[89] = ~layer_1[94]; 
    assign layer_2[90] = layer_1[79] | layer_1[102]; 
    assign layer_2[91] = ~layer_1[97]; 
    assign layer_2[92] = ~layer_1[80] | (layer_1[80] & layer_1[101]); 
    assign layer_2[93] = 1'b0; 
    assign layer_2[94] = layer_1[102] & ~layer_1[101]; 
    assign layer_2[95] = layer_1[103]; 
    assign layer_2[96] = ~(layer_1[101] ^ layer_1[107]); 
    assign layer_2[97] = ~layer_1[89] | (layer_1[107] & layer_1[89]); 
    assign layer_2[98] = ~layer_1[89] | (layer_1[92] & layer_1[89]); 
    assign layer_2[99] = ~layer_1[86] | (layer_1[86] & layer_1[90]); 
    assign layer_2[100] = 1'b0; 
    assign layer_2[101] = layer_1[110]; 
    assign layer_2[102] = ~layer_1[103] | (layer_1[92] & layer_1[103]); 
    assign layer_2[103] = layer_1[98] | layer_1[104]; 
    assign layer_2[104] = 1'b0; 
    assign layer_2[105] = 1'b1; 
    assign layer_2[106] = ~layer_1[122]; 
    assign layer_2[107] = ~(layer_1[107] | layer_1[94]); 
    assign layer_2[108] = layer_1[97] & ~layer_1[122]; 
    assign layer_2[109] = ~(layer_1[120] ^ layer_1[117]); 
    assign layer_2[110] = layer_1[116] ^ layer_1[117]; 
    assign layer_2[111] = 1'b0; 
    assign layer_2[112] = ~layer_1[118]; 
    assign layer_2[113] = layer_1[129] | layer_1[110]; 
    assign layer_2[114] = layer_1[122]; 
    assign layer_2[115] = layer_1[128] ^ layer_1[115]; 
    assign layer_2[116] = ~layer_1[114]; 
    assign layer_2[117] = 1'b1; 
    assign layer_2[118] = layer_1[104]; 
    assign layer_2[119] = ~layer_1[127] | (layer_1[127] & layer_1[134]); 
    assign layer_2[120] = layer_1[107] & layer_1[135]; 
    assign layer_2[121] = layer_1[111] & layer_1[133]; 
    assign layer_2[122] = 1'b1; 
    assign layer_2[123] = ~(layer_1[138] | layer_1[109]); 
    assign layer_2[124] = layer_1[132] & layer_1[138]; 
    assign layer_2[125] = ~layer_1[130] | (layer_1[130] & layer_1[137]); 
    assign layer_2[126] = ~(layer_1[128] ^ layer_1[124]); 
    assign layer_2[127] = ~layer_1[132] | (layer_1[113] & layer_1[132]); 
    assign layer_2[128] = ~layer_1[122] | (layer_1[122] & layer_1[131]); 
    assign layer_2[129] = ~(layer_1[141] & layer_1[126]); 
    assign layer_2[130] = ~(layer_1[136] | layer_1[125]); 
    assign layer_2[131] = layer_1[120] & ~layer_1[116]; 
    assign layer_2[132] = layer_1[140] & ~layer_1[132]; 
    assign layer_2[133] = layer_1[118] & layer_1[123]; 
    assign layer_2[134] = layer_1[122] & ~layer_1[147]; 
    assign layer_2[135] = ~layer_1[126] | (layer_1[128] & layer_1[126]); 
    assign layer_2[136] = ~layer_1[142]; 
    assign layer_2[137] = layer_1[132] & layer_1[125]; 
    assign layer_2[138] = ~layer_1[134] | (layer_1[125] & layer_1[134]); 
    assign layer_2[139] = layer_1[127]; 
    assign layer_2[140] = layer_1[148]; 
    assign layer_2[141] = ~layer_1[144] | (layer_1[131] & layer_1[144]); 
    assign layer_2[142] = layer_1[140] ^ layer_1[141]; 
    assign layer_2[143] = layer_1[131]; 
    assign layer_2[144] = ~(layer_1[143] | layer_1[152]); 
    assign layer_2[145] = layer_1[142]; 
    assign layer_2[146] = ~layer_1[135]; 
    assign layer_2[147] = layer_1[137] & ~layer_1[130]; 
    assign layer_2[148] = layer_1[159] & layer_1[149]; 
    assign layer_2[149] = 1'b0; 
    assign layer_2[150] = 1'b1; 
    assign layer_2[151] = layer_1[154]; 
    assign layer_2[152] = 1'b0; 
    assign layer_2[153] = ~layer_1[147]; 
    assign layer_2[154] = ~(layer_1[166] ^ layer_1[139]); 
    assign layer_2[155] = layer_1[155]; 
    assign layer_2[156] = layer_1[140] & ~layer_1[164]; 
    assign layer_2[157] = ~(layer_1[154] ^ layer_1[172]); 
    assign layer_2[158] = layer_1[148] | layer_1[147]; 
    assign layer_2[159] = 1'b0; 
    assign layer_2[160] = ~(layer_1[163] | layer_1[150]); 
    assign layer_2[161] = 1'b1; 
    assign layer_2[162] = layer_1[152] ^ layer_1[160]; 
    assign layer_2[163] = layer_1[173] ^ layer_1[149]; 
    assign layer_2[164] = ~layer_1[164] | (layer_1[164] & layer_1[165]); 
    assign layer_2[165] = layer_1[180] ^ layer_1[174]; 
    assign layer_2[166] = ~layer_1[162]; 
    assign layer_2[167] = 1'b1; 
    assign layer_2[168] = layer_1[156]; 
    assign layer_2[169] = ~layer_1[169] | (layer_1[169] & layer_1[181]); 
    assign layer_2[170] = ~(layer_1[162] ^ layer_1[156]); 
    assign layer_2[171] = ~layer_1[155]; 
    assign layer_2[172] = 1'b0; 
    assign layer_2[173] = layer_1[161] | layer_1[172]; 
    assign layer_2[174] = ~layer_1[164] | (layer_1[164] & layer_1[189]); 
    assign layer_2[175] = ~layer_1[176] | (layer_1[181] & layer_1[176]); 
    assign layer_2[176] = ~layer_1[176] | (layer_1[176] & layer_1[175]); 
    assign layer_2[177] = layer_1[184] & ~layer_1[166]; 
    assign layer_2[178] = ~layer_1[177] | (layer_1[165] & layer_1[177]); 
    assign layer_2[179] = 1'b1; 
    assign layer_2[180] = ~(layer_1[196] ^ layer_1[180]); 
    assign layer_2[181] = 1'b0; 
    assign layer_2[182] = ~layer_1[166]; 
    assign layer_2[183] = 1'b1; 
    assign layer_2[184] = ~layer_1[181]; 
    assign layer_2[185] = layer_1[187] ^ layer_1[178]; 
    assign layer_2[186] = ~layer_1[183]; 
    assign layer_2[187] = ~(layer_1[178] & layer_1[179]); 
    assign layer_2[188] = layer_1[180]; 
    assign layer_2[189] = ~(layer_1[198] | layer_1[176]); 
    assign layer_2[190] = layer_1[174] | layer_1[193]; 
    assign layer_2[191] = layer_1[182] ^ layer_1[205]; 
    assign layer_2[192] = layer_1[196] ^ layer_1[191]; 
    assign layer_2[193] = ~(layer_1[193] ^ layer_1[199]); 
    assign layer_2[194] = ~layer_1[197]; 
    assign layer_2[195] = ~(layer_1[182] | layer_1[198]); 
    assign layer_2[196] = layer_1[204]; 
    assign layer_2[197] = layer_1[202] | layer_1[210]; 
    assign layer_2[198] = ~layer_1[201] | (layer_1[204] & layer_1[201]); 
    assign layer_2[199] = layer_1[214] ^ layer_1[207]; 
    assign layer_2[200] = layer_1[207]; 
    assign layer_2[201] = layer_1[205] & ~layer_1[185]; 
    assign layer_2[202] = ~layer_1[199] | (layer_1[199] & layer_1[203]); 
    assign layer_2[203] = ~layer_1[192] | (layer_1[192] & layer_1[212]); 
    assign layer_2[204] = ~layer_1[188] | (layer_1[188] & layer_1[204]); 
    assign layer_2[205] = ~(layer_1[219] ^ layer_1[216]); 
    assign layer_2[206] = ~layer_1[208] | (layer_1[208] & layer_1[212]); 
    assign layer_2[207] = layer_1[203] ^ layer_1[222]; 
    assign layer_2[208] = layer_1[208]; 
    assign layer_2[209] = 1'b0; 
    assign layer_2[210] = layer_1[215]; 
    assign layer_2[211] = layer_1[217] ^ layer_1[223]; 
    assign layer_2[212] = ~(layer_1[204] & layer_1[221]); 
    assign layer_2[213] = ~layer_1[198] | (layer_1[198] & layer_1[211]); 
    assign layer_2[214] = layer_1[208] & ~layer_1[204]; 
    assign layer_2[215] = ~(layer_1[215] ^ layer_1[219]); 
    assign layer_2[216] = ~layer_1[203]; 
    assign layer_2[217] = layer_1[231]; 
    assign layer_2[218] = layer_1[226] & ~layer_1[219]; 
    assign layer_2[219] = layer_1[227] ^ layer_1[227]; 
    assign layer_2[220] = layer_1[232] ^ layer_1[232]; 
    assign layer_2[221] = layer_1[237] | layer_1[204]; 
    assign layer_2[222] = layer_1[226] ^ layer_1[213]; 
    assign layer_2[223] = layer_1[231] | layer_1[223]; 
    assign layer_2[224] = ~layer_1[229] | (layer_1[229] & layer_1[235]); 
    assign layer_2[225] = layer_1[232] & ~layer_1[228]; 
    assign layer_2[226] = layer_1[238] & ~layer_1[221]; 
    assign layer_2[227] = layer_1[228] & ~layer_1[211]; 
    assign layer_2[228] = 1'b1; 
    assign layer_2[229] = layer_1[242] & ~layer_1[242]; 
    assign layer_2[230] = layer_1[230] & ~layer_1[246]; 
    assign layer_2[231] = layer_1[242] | layer_1[215]; 
    assign layer_2[232] = 1'b1; 
    assign layer_2[233] = ~(layer_1[221] & layer_1[235]); 
    assign layer_2[234] = ~(layer_1[242] & layer_1[236]); 
    assign layer_2[235] = layer_1[241] ^ layer_1[224]; 
    assign layer_2[236] = ~(layer_1[233] & layer_1[230]); 
    assign layer_2[237] = layer_1[239] & layer_1[252]; 
    assign layer_2[238] = layer_1[240] & ~layer_1[232]; 
    assign layer_2[239] = 1'b1; 
    assign layer_2[240] = 1'b1; 
    assign layer_2[241] = 1'b0; 
    assign layer_2[242] = ~(layer_1[229] & layer_1[225]); 
    assign layer_2[243] = layer_1[232] | layer_1[241]; 
    assign layer_2[244] = layer_1[234] & ~layer_1[245]; 
    assign layer_2[245] = layer_1[240] & ~layer_1[245]; 
    assign layer_2[246] = ~layer_1[250] | (layer_1[250] & layer_1[243]); 
    assign layer_2[247] = ~(layer_1[261] & layer_1[238]); 
    assign layer_2[248] = ~layer_1[255] | (layer_1[255] & layer_1[250]); 
    assign layer_2[249] = layer_1[254]; 
    assign layer_2[250] = layer_1[241] & layer_1[253]; 
    assign layer_2[251] = layer_1[263] | layer_1[243]; 
    assign layer_2[252] = layer_1[236]; 
    assign layer_2[253] = 1'b1; 
    assign layer_2[254] = ~layer_1[263] | (layer_1[239] & layer_1[263]); 
    assign layer_2[255] = layer_1[251] & ~layer_1[248]; 
    assign layer_2[256] = layer_1[240] ^ layer_1[252]; 
    assign layer_2[257] = layer_1[247] ^ layer_1[248]; 
    assign layer_2[258] = ~layer_1[241]; 
    assign layer_2[259] = ~(layer_1[248] ^ layer_1[243]); 
    assign layer_2[260] = layer_1[272] & ~layer_1[250]; 
    assign layer_2[261] = ~layer_1[252]; 
    assign layer_2[262] = ~layer_1[270]; 
    assign layer_2[263] = ~(layer_1[261] & layer_1[259]); 
    assign layer_2[264] = ~(layer_1[278] ^ layer_1[272]); 
    assign layer_2[265] = layer_1[268] ^ layer_1[248]; 
    assign layer_2[266] = ~(layer_1[264] | layer_1[252]); 
    assign layer_2[267] = ~layer_1[268]; 
    assign layer_2[268] = layer_1[262]; 
    assign layer_2[269] = layer_1[262] & layer_1[253]; 
    assign layer_2[270] = ~layer_1[285]; 
    assign layer_2[271] = 1'b1; 
    assign layer_2[272] = layer_1[258]; 
    assign layer_2[273] = ~(layer_1[289] ^ layer_1[264]); 
    assign layer_2[274] = layer_1[264] & layer_1[284]; 
    assign layer_2[275] = ~layer_1[270]; 
    assign layer_2[276] = 1'b0; 
    assign layer_2[277] = layer_1[271] & ~layer_1[292]; 
    assign layer_2[278] = ~layer_1[276] | (layer_1[278] & layer_1[276]); 
    assign layer_2[279] = ~layer_1[264]; 
    assign layer_2[280] = ~(layer_1[277] | layer_1[272]); 
    assign layer_2[281] = 1'b1; 
    assign layer_2[282] = layer_1[278] & layer_1[297]; 
    assign layer_2[283] = layer_1[271] ^ layer_1[273]; 
    assign layer_2[284] = layer_1[291] & layer_1[286]; 
    assign layer_2[285] = ~layer_1[273]; 
    assign layer_2[286] = ~layer_1[273]; 
    assign layer_2[287] = layer_1[282]; 
    assign layer_2[288] = ~(layer_1[278] & layer_1[283]); 
    assign layer_2[289] = layer_1[295]; 
    assign layer_2[290] = layer_1[304] ^ layer_1[297]; 
    assign layer_2[291] = layer_1[299]; 
    assign layer_2[292] = layer_1[282] ^ layer_1[299]; 
    assign layer_2[293] = layer_1[278]; 
    assign layer_2[294] = ~layer_1[281] | (layer_1[281] & layer_1[279]); 
    assign layer_2[295] = layer_1[283] ^ layer_1[291]; 
    assign layer_2[296] = ~layer_1[285] | (layer_1[285] & layer_1[288]); 
    assign layer_2[297] = layer_1[304]; 
    assign layer_2[298] = layer_1[298] | layer_1[283]; 
    assign layer_2[299] = ~(layer_1[314] | layer_1[314]); 
    assign layer_2[300] = ~(layer_1[312] & layer_1[296]); 
    assign layer_2[301] = layer_1[296] ^ layer_1[285]; 
    assign layer_2[302] = ~(layer_1[310] | layer_1[313]); 
    assign layer_2[303] = layer_1[311] | layer_1[298]; 
    assign layer_2[304] = layer_1[312] | layer_1[317]; 
    assign layer_2[305] = layer_1[302] & ~layer_1[320]; 
    assign layer_2[306] = 1'b0; 
    assign layer_2[307] = layer_1[296] & layer_1[290]; 
    assign layer_2[308] = ~layer_1[322]; 
    assign layer_2[309] = layer_1[308]; 
    assign layer_2[310] = ~layer_1[312]; 
    assign layer_2[311] = layer_1[326]; 
    assign layer_2[312] = layer_1[325] & ~layer_1[311]; 
    assign layer_2[313] = ~(layer_1[315] & layer_1[318]); 
    assign layer_2[314] = 1'b1; 
    assign layer_2[315] = layer_1[317] ^ layer_1[303]; 
    assign layer_2[316] = ~layer_1[331]; 
    assign layer_2[317] = ~layer_1[332]; 
    assign layer_2[318] = ~layer_1[304]; 
    assign layer_2[319] = ~layer_1[323] | (layer_1[310] & layer_1[323]); 
    assign layer_2[320] = ~(layer_1[318] | layer_1[322]); 
    assign layer_2[321] = 1'b0; 
    assign layer_2[322] = ~(layer_1[322] & layer_1[327]); 
    assign layer_2[323] = layer_1[329]; 
    assign layer_2[324] = ~layer_1[315] | (layer_1[315] & layer_1[319]); 
    assign layer_2[325] = ~(layer_1[318] | layer_1[326]); 
    assign layer_2[326] = layer_1[322] ^ layer_1[321]; 
    assign layer_2[327] = ~(layer_1[313] & layer_1[314]); 
    assign layer_2[328] = layer_1[314] ^ layer_1[339]; 
    assign layer_2[329] = ~layer_1[316] | (layer_1[344] & layer_1[316]); 
    assign layer_2[330] = ~layer_1[344] | (layer_1[343] & layer_1[344]); 
    assign layer_2[331] = ~layer_1[335]; 
    assign layer_2[332] = layer_1[331] & ~layer_1[323]; 
    assign layer_2[333] = 1'b0; 
    assign layer_2[334] = layer_1[329] & layer_1[344]; 
    assign layer_2[335] = ~(layer_1[335] ^ layer_1[341]); 
    assign layer_2[336] = layer_1[325] & ~layer_1[335]; 
    assign layer_2[337] = ~layer_1[322]; 
    assign layer_2[338] = 1'b0; 
    assign layer_2[339] = layer_1[325]; 
    assign layer_2[340] = layer_1[331] & ~layer_1[348]; 
    assign layer_2[341] = ~layer_1[331] | (layer_1[331] & layer_1[332]); 
    assign layer_2[342] = ~(layer_1[338] ^ layer_1[346]); 
    assign layer_2[343] = layer_1[340] | layer_1[326]; 
    assign layer_2[344] = 1'b0; 
    assign layer_2[345] = layer_1[348] & ~layer_1[336]; 
    assign layer_2[346] = ~(layer_1[361] & layer_1[341]); 
    assign layer_2[347] = layer_1[347]; 
    assign layer_2[348] = ~(layer_1[333] & layer_1[354]); 
    assign layer_2[349] = ~(layer_1[339] & layer_1[364]); 
    assign layer_2[350] = ~(layer_1[338] ^ layer_1[357]); 
    assign layer_2[351] = ~layer_1[342]; 
    assign layer_2[352] = ~(layer_1[340] ^ layer_1[336]); 
    assign layer_2[353] = layer_1[337]; 
    assign layer_2[354] = layer_1[347] & ~layer_1[356]; 
    assign layer_2[355] = 1'b1; 
    assign layer_2[356] = ~layer_1[368] | (layer_1[368] & layer_1[366]); 
    assign layer_2[357] = 1'b0; 
    assign layer_2[358] = layer_1[356] & ~layer_1[368]; 
    assign layer_2[359] = layer_1[349] & ~layer_1[359]; 
    assign layer_2[360] = ~(layer_1[372] | layer_1[348]); 
    assign layer_2[361] = ~(layer_1[372] & layer_1[344]); 
    assign layer_2[362] = layer_1[376] ^ layer_1[377]; 
    assign layer_2[363] = layer_1[369] ^ layer_1[373]; 
    assign layer_2[364] = ~(layer_1[366] ^ layer_1[379]); 
    assign layer_2[365] = 1'b0; 
    assign layer_2[366] = layer_1[364] | layer_1[354]; 
    assign layer_2[367] = ~(layer_1[378] | layer_1[362]); 
    assign layer_2[368] = ~layer_1[355] | (layer_1[372] & layer_1[355]); 
    assign layer_2[369] = ~layer_1[354] | (layer_1[354] & layer_1[362]); 
    assign layer_2[370] = layer_1[354]; 
    assign layer_2[371] = ~layer_1[357]; 
    assign layer_2[372] = layer_1[365]; 
    assign layer_2[373] = layer_1[372] & ~layer_1[375]; 
    assign layer_2[374] = ~(layer_1[381] & layer_1[357]); 
    assign layer_2[375] = layer_1[384]; 
    assign layer_2[376] = 1'b0; 
    assign layer_2[377] = layer_1[377] & ~layer_1[367]; 
    assign layer_2[378] = layer_1[371] & ~layer_1[373]; 
    assign layer_2[379] = ~(layer_1[391] | layer_1[368]); 
    assign layer_2[380] = layer_1[369] & ~layer_1[386]; 
    assign layer_2[381] = layer_1[382] & ~layer_1[382]; 
    assign layer_2[382] = ~layer_1[367] | (layer_1[367] & layer_1[372]); 
    assign layer_2[383] = ~layer_1[382] | (layer_1[382] & layer_1[393]); 
    assign layer_2[384] = ~layer_1[370] | (layer_1[370] & layer_1[399]); 
    assign layer_2[385] = ~layer_1[381] | (layer_1[381] & layer_1[379]); 
    assign layer_2[386] = ~(layer_1[371] | layer_1[391]); 
    assign layer_2[387] = ~(layer_1[373] ^ layer_1[392]); 
    assign layer_2[388] = layer_1[382]; 
    assign layer_2[389] = ~(layer_1[383] ^ layer_1[391]); 
    assign layer_2[390] = layer_1[394] ^ layer_1[403]; 
    assign layer_2[391] = 1'b1; 
    assign layer_2[392] = layer_1[387] | layer_1[386]; 
    assign layer_2[393] = ~(layer_1[409] & layer_1[400]); 
    assign layer_2[394] = layer_1[408] & layer_1[386]; 
    assign layer_2[395] = layer_1[406] | layer_1[393]; 
    assign layer_2[396] = 1'b0; 
    assign layer_2[397] = layer_1[393] & ~layer_1[394]; 
    assign layer_2[398] = ~(layer_1[396] & layer_1[402]); 
    assign layer_2[399] = ~layer_1[384]; 
    assign layer_2[400] = ~layer_1[399] | (layer_1[392] & layer_1[399]); 
    assign layer_2[401] = ~layer_1[415]; 
    assign layer_2[402] = layer_1[410] & ~layer_1[390]; 
    assign layer_2[403] = ~layer_1[390] | (layer_1[407] & layer_1[390]); 
    assign layer_2[404] = layer_1[394] & ~layer_1[392]; 
    assign layer_2[405] = layer_1[407] ^ layer_1[400]; 
    assign layer_2[406] = ~layer_1[407]; 
    assign layer_2[407] = ~(layer_1[396] ^ layer_1[398]); 
    assign layer_2[408] = ~(layer_1[415] | layer_1[418]); 
    assign layer_2[409] = 1'b0; 
    assign layer_2[410] = ~layer_1[415]; 
    assign layer_2[411] = layer_1[401]; 
    assign layer_2[412] = ~(layer_1[415] & layer_1[396]); 
    assign layer_2[413] = ~(layer_1[400] & layer_1[427]); 
    assign layer_2[414] = layer_1[410] & layer_1[404]; 
    assign layer_2[415] = layer_1[406]; 
    assign layer_2[416] = ~(layer_1[419] | layer_1[420]); 
    assign layer_2[417] = ~layer_1[428]; 
    assign layer_2[418] = ~layer_1[426] | (layer_1[426] & layer_1[415]); 
    assign layer_2[419] = 1'b0; 
    assign layer_2[420] = layer_1[413]; 
    assign layer_2[421] = ~(layer_1[427] & layer_1[404]); 
    assign layer_2[422] = ~layer_1[432]; 
    assign layer_2[423] = layer_1[409] ^ layer_1[433]; 
    assign layer_2[424] = ~(layer_1[419] | layer_1[438]); 
    assign layer_2[425] = layer_1[424] ^ layer_1[420]; 
    assign layer_2[426] = 1'b0; 
    assign layer_2[427] = ~layer_1[421]; 
    assign layer_2[428] = 1'b1; 
    assign layer_2[429] = ~layer_1[428]; 
    assign layer_2[430] = ~layer_1[423]; 
    assign layer_2[431] = ~layer_1[445] | (layer_1[422] & layer_1[445]); 
    assign layer_2[432] = layer_1[438] | layer_1[443]; 
    assign layer_2[433] = 1'b1; 
    assign layer_2[434] = layer_1[441] ^ layer_1[428]; 
    assign layer_2[435] = 1'b0; 
    assign layer_2[436] = layer_1[450]; 
    assign layer_2[437] = 1'b1; 
    assign layer_2[438] = ~layer_1[430] | (layer_1[441] & layer_1[430]); 
    assign layer_2[439] = 1'b0; 
    assign layer_2[440] = 1'b0; 
    assign layer_2[441] = ~layer_1[430] | (layer_1[430] & layer_1[453]); 
    assign layer_2[442] = layer_1[452] & ~layer_1[450]; 
    assign layer_2[443] = layer_1[456]; 
    assign layer_2[444] = layer_1[445] | layer_1[433]; 
    assign layer_2[445] = layer_1[439] ^ layer_1[447]; 
    assign layer_2[446] = ~layer_1[449] | (layer_1[449] & layer_1[439]); 
    assign layer_2[447] = layer_1[446] & ~layer_1[431]; 
    assign layer_2[448] = ~(layer_1[457] | layer_1[432]); 
    assign layer_2[449] = layer_1[458] | layer_1[436]; 
    assign layer_2[450] = layer_1[445]; 
    assign layer_2[451] = layer_1[457] & ~layer_1[463]; 
    assign layer_2[452] = ~(layer_1[443] ^ layer_1[451]); 
    assign layer_2[453] = ~layer_1[438] | (layer_1[438] & layer_1[443]); 
    assign layer_2[454] = 1'b1; 
    assign layer_2[455] = layer_1[471]; 
    assign layer_2[456] = 1'b0; 
    assign layer_2[457] = ~layer_1[453]; 
    assign layer_2[458] = ~layer_1[472]; 
    assign layer_2[459] = 1'b0; 
    assign layer_2[460] = ~(layer_1[463] ^ layer_1[458]); 
    assign layer_2[461] = ~(layer_1[451] ^ layer_1[450]); 
    assign layer_2[462] = ~layer_1[463] | (layer_1[477] & layer_1[463]); 
    assign layer_2[463] = 1'b0; 
    assign layer_2[464] = ~(layer_1[465] | layer_1[461]); 
    assign layer_2[465] = ~layer_1[471]; 
    assign layer_2[466] = layer_1[463] | layer_1[478]; 
    assign layer_2[467] = ~(layer_1[481] | layer_1[473]); 
    assign layer_2[468] = ~layer_1[453] | (layer_1[453] & layer_1[453]); 
    assign layer_2[469] = ~layer_1[463]; 
    assign layer_2[470] = layer_1[476] ^ layer_1[480]; 
    assign layer_2[471] = ~layer_1[487] | (layer_1[487] & layer_1[468]); 
    assign layer_2[472] = layer_1[464]; 
    assign layer_2[473] = ~(layer_1[477] & layer_1[456]); 
    assign layer_2[474] = ~(layer_1[479] | layer_1[476]); 
    assign layer_2[475] = layer_1[470] & layer_1[471]; 
    assign layer_2[476] = layer_1[490]; 
    assign layer_2[477] = ~layer_1[465] | (layer_1[465] & layer_1[466]); 
    assign layer_2[478] = layer_1[493] & ~layer_1[480]; 
    assign layer_2[479] = layer_1[493]; 
    assign layer_2[480] = 1'b0; 
    assign layer_2[481] = ~layer_1[468]; 
    assign layer_2[482] = layer_1[494] | layer_1[473]; 
    assign layer_2[483] = 1'b0; 
    assign layer_2[484] = 1'b1; 
    assign layer_2[485] = layer_1[493]; 
    assign layer_2[486] = ~(layer_1[478] & layer_1[481]); 
    assign layer_2[487] = ~layer_1[474]; 
    assign layer_2[488] = ~(layer_1[503] | layer_1[477]); 
    assign layer_2[489] = 1'b1; 
    assign layer_2[490] = ~(layer_1[485] | layer_1[485]); 
    assign layer_2[491] = ~layer_1[496] | (layer_1[496] & layer_1[503]); 
    assign layer_2[492] = ~layer_1[501] | (layer_1[501] & layer_1[490]); 
    assign layer_2[493] = 1'b1; 
    assign layer_2[494] = 1'b0; 
    assign layer_2[495] = layer_1[486] ^ layer_1[507]; 
    assign layer_2[496] = ~(layer_1[507] | layer_1[490]); 
    assign layer_2[497] = layer_1[505]; 
    assign layer_2[498] = ~layer_1[507]; 
    assign layer_2[499] = layer_1[501] & ~layer_1[494]; 
    assign layer_2[500] = ~(layer_1[488] & layer_1[492]); 
    assign layer_2[501] = layer_1[499]; 
    assign layer_2[502] = layer_1[515] ^ layer_1[499]; 
    assign layer_2[503] = ~layer_1[519] | (layer_1[519] & layer_1[491]); 
    assign layer_2[504] = layer_1[514]; 
    assign layer_2[505] = layer_1[494] | layer_1[490]; 
    assign layer_2[506] = ~(layer_1[513] ^ layer_1[516]); 
    assign layer_2[507] = ~(layer_1[521] | layer_1[496]); 
    assign layer_2[508] = layer_1[492]; 
    assign layer_2[509] = layer_1[512] & ~layer_1[497]; 
    assign layer_2[510] = layer_1[513]; 
    assign layer_2[511] = layer_1[523] ^ layer_1[514]; 
    assign layer_2[512] = ~(layer_1[508] ^ layer_1[497]); 
    assign layer_2[513] = ~layer_1[502]; 
    assign layer_2[514] = layer_1[529]; 
    assign layer_2[515] = ~layer_1[510] | (layer_1[512] & layer_1[510]); 
    assign layer_2[516] = ~layer_1[513] | (layer_1[513] & layer_1[513]); 
    assign layer_2[517] = ~layer_1[505]; 
    assign layer_2[518] = layer_1[523]; 
    assign layer_2[519] = 1'b0; 
    assign layer_2[520] = ~(layer_1[508] & layer_1[528]); 
    assign layer_2[521] = layer_1[511] & ~layer_1[527]; 
    assign layer_2[522] = ~(layer_1[510] ^ layer_1[507]); 
    assign layer_2[523] = ~(layer_1[520] | layer_1[507]); 
    assign layer_2[524] = layer_1[519] | layer_1[514]; 
    assign layer_2[525] = layer_1[530] & ~layer_1[519]; 
    assign layer_2[526] = layer_1[532]; 
    assign layer_2[527] = ~layer_1[514] | (layer_1[514] & layer_1[541]); 
    assign layer_2[528] = ~layer_1[521]; 
    assign layer_2[529] = layer_1[518] & ~layer_1[517]; 
    assign layer_2[530] = 1'b1; 
    assign layer_2[531] = layer_1[531] & ~layer_1[525]; 
    assign layer_2[532] = layer_1[539]; 
    assign layer_2[533] = ~layer_1[530]; 
    assign layer_2[534] = 1'b0; 
    assign layer_2[535] = layer_1[548] & ~layer_1[534]; 
    assign layer_2[536] = ~layer_1[546] | (layer_1[541] & layer_1[546]); 
    assign layer_2[537] = ~layer_1[552]; 
    assign layer_2[538] = ~layer_1[551]; 
    assign layer_2[539] = ~layer_1[547]; 
    assign layer_2[540] = ~layer_1[537]; 
    assign layer_2[541] = ~layer_1[527] | (layer_1[527] & layer_1[524]); 
    assign layer_2[542] = layer_1[534] ^ layer_1[536]; 
    assign layer_2[543] = layer_1[538] ^ layer_1[532]; 
    assign layer_2[544] = layer_1[542] & ~layer_1[551]; 
    assign layer_2[545] = ~layer_1[549] | (layer_1[537] & layer_1[549]); 
    assign layer_2[546] = ~layer_1[533] | (layer_1[533] & layer_1[537]); 
    assign layer_2[547] = layer_1[531] & ~layer_1[538]; 
    assign layer_2[548] = ~layer_1[559] | (layer_1[559] & layer_1[542]); 
    assign layer_2[549] = layer_1[563]; 
    assign layer_2[550] = 1'b1; 
    assign layer_2[551] = layer_1[534] & ~layer_1[537]; 
    assign layer_2[552] = 1'b0; 
    assign layer_2[553] = 1'b0; 
    assign layer_2[554] = ~(layer_1[548] | layer_1[554]); 
    assign layer_2[555] = ~layer_1[546] | (layer_1[546] & layer_1[550]); 
    assign layer_2[556] = ~layer_1[547]; 
    assign layer_2[557] = 1'b0; 
    assign layer_2[558] = ~layer_1[548]; 
    assign layer_2[559] = layer_1[564] ^ layer_1[561]; 
    assign layer_2[560] = ~(layer_1[575] & layer_1[558]); 
    assign layer_2[561] = 1'b0; 
    assign layer_2[562] = ~layer_1[562] | (layer_1[563] & layer_1[562]); 
    assign layer_2[563] = ~(layer_1[555] ^ layer_1[578]); 
    assign layer_2[564] = ~layer_1[552]; 
    assign layer_2[565] = ~layer_1[552]; 
    assign layer_2[566] = ~layer_1[552] | (layer_1[552] & layer_1[556]); 
    assign layer_2[567] = ~layer_1[570]; 
    assign layer_2[568] = layer_1[578] & ~layer_1[572]; 
    assign layer_2[569] = ~layer_1[579]; 
    assign layer_2[570] = layer_1[578]; 
    assign layer_2[571] = ~(layer_1[555] & layer_1[573]); 
    assign layer_2[572] = ~(layer_1[559] & layer_1[577]); 
    assign layer_2[573] = layer_1[573] & ~layer_1[568]; 
    assign layer_2[574] = ~(layer_1[569] | layer_1[572]); 
    assign layer_2[575] = layer_1[590]; 
    assign layer_2[576] = ~layer_1[563] | (layer_1[563] & layer_1[573]); 
    assign layer_2[577] = layer_1[561]; 
    assign layer_2[578] = 1'b1; 
    assign layer_2[579] = ~layer_1[588] | (layer_1[575] & layer_1[588]); 
    assign layer_2[580] = layer_1[586] & ~layer_1[595]; 
    assign layer_2[581] = layer_1[576] & ~layer_1[585]; 
    assign layer_2[582] = layer_1[566]; 
    assign layer_2[583] = ~(layer_1[572] ^ layer_1[585]); 
    assign layer_2[584] = ~(layer_1[598] & layer_1[580]); 
    assign layer_2[585] = ~layer_1[585] | (layer_1[582] & layer_1[585]); 
    assign layer_2[586] = layer_1[581]; 
    assign layer_2[587] = layer_1[590] & ~layer_1[588]; 
    assign layer_2[588] = 1'b0; 
    assign layer_2[589] = ~(layer_1[597] & layer_1[589]); 
    assign layer_2[590] = layer_1[597]; 
    assign layer_2[591] = layer_1[601] & ~layer_1[598]; 
    assign layer_2[592] = ~(layer_1[606] ^ layer_1[600]); 
    assign layer_2[593] = ~layer_1[583]; 
    assign layer_2[594] = layer_1[579] & layer_1[590]; 
    assign layer_2[595] = layer_1[579] ^ layer_1[589]; 
    assign layer_2[596] = layer_1[589]; 
    assign layer_2[597] = ~layer_1[587] | (layer_1[586] & layer_1[587]); 
    assign layer_2[598] = ~layer_1[588] | (layer_1[582] & layer_1[588]); 
    assign layer_2[599] = layer_1[593] & ~layer_1[601]; 
    assign layer_2[600] = layer_1[615]; 
    assign layer_2[601] = 1'b0; 
    assign layer_2[602] = layer_1[611] & layer_1[601]; 
    assign layer_2[603] = layer_1[607] & layer_1[588]; 
    assign layer_2[604] = ~layer_1[611]; 
    assign layer_2[605] = ~layer_1[620]; 
    assign layer_2[606] = ~layer_1[601] | (layer_1[601] & layer_1[609]); 
    assign layer_2[607] = layer_1[599] | layer_1[617]; 
    assign layer_2[608] = layer_1[617] & ~layer_1[604]; 
    assign layer_2[609] = layer_1[624]; 
    assign layer_2[610] = layer_1[602] ^ layer_1[605]; 
    assign layer_2[611] = layer_1[624] & layer_1[612]; 
    assign layer_2[612] = layer_1[597] & ~layer_1[614]; 
    assign layer_2[613] = layer_1[611] & ~layer_1[596]; 
    assign layer_2[614] = ~layer_1[622] | (layer_1[622] & layer_1[624]); 
    assign layer_2[615] = ~(layer_1[623] ^ layer_1[615]); 
    assign layer_2[616] = layer_1[631]; 
    assign layer_2[617] = ~layer_1[622] | (layer_1[603] & layer_1[622]); 
    assign layer_2[618] = ~(layer_1[627] ^ layer_1[624]); 
    assign layer_2[619] = ~layer_1[627]; 
    assign layer_2[620] = ~(layer_1[625] ^ layer_1[635]); 
    assign layer_2[621] = layer_1[609] | layer_1[605]; 
    assign layer_2[622] = ~layer_1[611] | (layer_1[611] & layer_1[611]); 
    assign layer_2[623] = ~(layer_1[625] & layer_1[629]); 
    assign layer_2[624] = layer_1[617] & ~layer_1[614]; 
    assign layer_2[625] = ~(layer_1[633] & layer_1[625]); 
    assign layer_2[626] = layer_1[631]; 
    assign layer_2[627] = layer_1[636] & ~layer_1[616]; 
    assign layer_2[628] = ~layer_1[632]; 
    assign layer_2[629] = layer_1[630]; 
    assign layer_2[630] = ~layer_1[622] | (layer_1[631] & layer_1[622]); 
    assign layer_2[631] = ~layer_1[621] | (layer_1[621] & layer_1[624]); 
    assign layer_2[632] = 1'b0; 
    assign layer_2[633] = 1'b1; 
    assign layer_2[634] = 1'b0; 
    assign layer_2[635] = ~layer_1[646] | (layer_1[646] & layer_1[639]); 
    assign layer_2[636] = ~layer_1[630]; 
    assign layer_2[637] = ~layer_1[647]; 
    assign layer_2[638] = layer_1[641]; 
    assign layer_2[639] = layer_1[649] & ~layer_1[632]; 
    assign layer_2[640] = ~layer_1[653]; 
    assign layer_2[641] = layer_1[632] ^ layer_1[626]; 
    assign layer_2[642] = 1'b1; 
    assign layer_2[643] = layer_1[652] | layer_1[649]; 
    assign layer_2[644] = ~layer_1[653]; 
    assign layer_2[645] = 1'b0; 
    assign layer_2[646] = layer_1[644]; 
    assign layer_2[647] = layer_1[650] & ~layer_1[638]; 
    assign layer_2[648] = ~layer_1[633] | (layer_1[643] & layer_1[633]); 
    assign layer_2[649] = ~layer_1[653]; 
    assign layer_2[650] = ~layer_1[666]; 
    assign layer_2[651] = ~layer_1[663]; 
    assign layer_2[652] = ~layer_1[645] | (layer_1[645] & layer_1[639]); 
    assign layer_2[653] = ~layer_1[647]; 
    assign layer_2[654] = layer_1[650]; 
    assign layer_2[655] = layer_1[645] & ~layer_1[663]; 
    assign layer_2[656] = ~(layer_1[659] & layer_1[649]); 
    assign layer_2[657] = ~(layer_1[662] ^ layer_1[658]); 
    assign layer_2[658] = 1'b0; 
    assign layer_2[659] = layer_1[675] & ~layer_1[649]; 
    assign layer_2[660] = layer_1[644]; 
    assign layer_2[661] = layer_1[664] & layer_1[656]; 
    assign layer_2[662] = ~(layer_1[670] & layer_1[654]); 
    assign layer_2[663] = layer_1[658] & ~layer_1[661]; 
    assign layer_2[664] = 1'b0; 
    assign layer_2[665] = ~(layer_1[654] | layer_1[648]); 
    assign layer_2[666] = layer_1[665] & ~layer_1[661]; 
    assign layer_2[667] = layer_1[654]; 
    assign layer_2[668] = ~(layer_1[663] | layer_1[678]); 
    assign layer_2[669] = ~(layer_1[673] & layer_1[675]); 
    assign layer_2[670] = layer_1[671] | layer_1[663]; 
    assign layer_2[671] = layer_1[666] | layer_1[656]; 
    assign layer_2[672] = layer_1[665]; 
    assign layer_2[673] = ~layer_1[669] | (layer_1[688] & layer_1[669]); 
    assign layer_2[674] = layer_1[670] & ~layer_1[658]; 
    assign layer_2[675] = ~(layer_1[676] | layer_1[689]); 
    assign layer_2[676] = 1'b0; 
    assign layer_2[677] = layer_1[689] & ~layer_1[677]; 
    assign layer_2[678] = ~layer_1[680]; 
    assign layer_2[679] = layer_1[685] & ~layer_1[663]; 
    assign layer_2[680] = layer_1[665] & layer_1[680]; 
    assign layer_2[681] = layer_1[674] | layer_1[681]; 
    assign layer_2[682] = layer_1[681] | layer_1[691]; 
    assign layer_2[683] = ~layer_1[693]; 
    assign layer_2[684] = layer_1[668] & layer_1[670]; 
    assign layer_2[685] = ~layer_1[699]; 
    assign layer_2[686] = layer_1[678]; 
    assign layer_2[687] = ~layer_1[695] | (layer_1[695] & layer_1[672]); 
    assign layer_2[688] = layer_1[704] ^ layer_1[702]; 
    assign layer_2[689] = layer_1[675] & ~layer_1[682]; 
    assign layer_2[690] = layer_1[681]; 
    assign layer_2[691] = ~(layer_1[679] ^ layer_1[697]); 
    assign layer_2[692] = layer_1[687] & ~layer_1[677]; 
    assign layer_2[693] = ~(layer_1[686] | layer_1[699]); 
    assign layer_2[694] = layer_1[693] ^ layer_1[698]; 
    assign layer_2[695] = ~(layer_1[702] ^ layer_1[687]); 
    assign layer_2[696] = 1'b1; 
    assign layer_2[697] = layer_1[709] & layer_1[691]; 
    assign layer_2[698] = layer_1[688] & layer_1[705]; 
    assign layer_2[699] = ~layer_1[711] | (layer_1[702] & layer_1[711]); 
    assign layer_2[700] = layer_1[690] | layer_1[697]; 
    assign layer_2[701] = layer_1[685] | layer_1[708]; 
    assign layer_2[702] = layer_1[689] & ~layer_1[690]; 
    assign layer_2[703] = ~layer_1[699] | (layer_1[701] & layer_1[699]); 
    assign layer_2[704] = 1'b0; 
    assign layer_2[705] = layer_1[691] & ~layer_1[718]; 
    assign layer_2[706] = ~layer_1[695]; 
    assign layer_2[707] = 1'b1; 
    assign layer_2[708] = layer_1[699] & ~layer_1[705]; 
    assign layer_2[709] = ~(layer_1[718] & layer_1[717]); 
    assign layer_2[710] = ~layer_1[710] | (layer_1[701] & layer_1[710]); 
    assign layer_2[711] = ~(layer_1[700] | layer_1[718]); 
    assign layer_2[712] = layer_1[710] & ~layer_1[706]; 
    assign layer_2[713] = ~(layer_1[717] ^ layer_1[714]); 
    assign layer_2[714] = 1'b0; 
    assign layer_2[715] = 1'b1; 
    assign layer_2[716] = layer_1[728]; 
    assign layer_2[717] = ~layer_1[714]; 
    assign layer_2[718] = ~(layer_1[709] ^ layer_1[701]); 
    assign layer_2[719] = ~layer_1[730] | (layer_1[730] & layer_1[702]); 
    assign layer_2[720] = layer_1[724]; 
    assign layer_2[721] = layer_1[715] ^ layer_1[709]; 
    assign layer_2[722] = layer_1[735]; 
    assign layer_2[723] = 1'b0; 
    assign layer_2[724] = ~layer_1[712]; 
    assign layer_2[725] = ~layer_1[719] | (layer_1[719] & layer_1[712]); 
    assign layer_2[726] = ~layer_1[720]; 
    assign layer_2[727] = 1'b1; 
    assign layer_2[728] = ~(layer_1[720] & layer_1[737]); 
    assign layer_2[729] = ~layer_1[738]; 
    assign layer_2[730] = ~layer_1[729] | (layer_1[737] & layer_1[729]); 
    assign layer_2[731] = ~layer_1[720] | (layer_1[720] & layer_1[741]); 
    assign layer_2[732] = ~(layer_1[744] ^ layer_1[741]); 
    assign layer_2[733] = layer_1[747] & layer_1[724]; 
    assign layer_2[734] = ~layer_1[730]; 
    assign layer_2[735] = layer_1[737] | layer_1[734]; 
    assign layer_2[736] = layer_1[730] | layer_1[722]; 
    assign layer_2[737] = layer_1[743]; 
    assign layer_2[738] = layer_1[746] & layer_1[726]; 
    assign layer_2[739] = ~layer_1[727] | (layer_1[748] & layer_1[727]); 
    assign layer_2[740] = ~layer_1[724]; 
    assign layer_2[741] = layer_1[726] | layer_1[730]; 
    assign layer_2[742] = ~(layer_1[731] ^ layer_1[753]); 
    assign layer_2[743] = layer_1[743] & layer_1[732]; 
    assign layer_2[744] = ~(layer_1[738] & layer_1[747]); 
    assign layer_2[745] = ~layer_1[739]; 
    assign layer_2[746] = layer_1[744] ^ layer_1[740]; 
    assign layer_2[747] = ~layer_1[740] | (layer_1[746] & layer_1[740]); 
    assign layer_2[748] = ~(layer_1[753] & layer_1[732]); 
    assign layer_2[749] = ~(layer_1[748] & layer_1[747]); 
    assign layer_2[750] = 1'b1; 
    assign layer_2[751] = ~(layer_1[761] & layer_1[743]); 
    assign layer_2[752] = ~(layer_1[753] & layer_1[736]); 
    assign layer_2[753] = ~(layer_1[753] ^ layer_1[754]); 
    assign layer_2[754] = layer_1[751]; 
    assign layer_2[755] = layer_1[759] | layer_1[770]; 
    assign layer_2[756] = ~layer_1[749]; 
    assign layer_2[757] = layer_1[758] | layer_1[756]; 
    assign layer_2[758] = ~layer_1[771]; 
    assign layer_2[759] = ~layer_1[753]; 
    assign layer_2[760] = ~layer_1[760] | (layer_1[760] & layer_1[760]); 
    assign layer_2[761] = ~layer_1[774]; 
    assign layer_2[762] = layer_1[761] & ~layer_1[772]; 
    assign layer_2[763] = 1'b0; 
    assign layer_2[764] = layer_1[774] | layer_1[764]; 
    assign layer_2[765] = ~layer_1[767]; 
    assign layer_2[766] = ~layer_1[769] | (layer_1[776] & layer_1[769]); 
    assign layer_2[767] = ~(layer_1[762] | layer_1[778]); 
    assign layer_2[768] = layer_1[760]; 
    assign layer_2[769] = layer_1[773] & ~layer_1[773]; 
    assign layer_2[770] = layer_1[771] ^ layer_1[780]; 
    assign layer_2[771] = ~(layer_1[768] | layer_1[757]); 
    assign layer_2[772] = ~(layer_1[761] | layer_1[766]); 
    assign layer_2[773] = ~layer_1[788] | (layer_1[788] & layer_1[759]); 
    assign layer_2[774] = layer_1[763]; 
    assign layer_2[775] = layer_1[764] ^ layer_1[762]; 
    assign layer_2[776] = layer_1[766] ^ layer_1[765]; 
    assign layer_2[777] = ~(layer_1[786] ^ layer_1[763]); 
    assign layer_2[778] = layer_1[777] & layer_1[769]; 
    assign layer_2[779] = layer_1[794] | layer_1[766]; 
    assign layer_2[780] = ~layer_1[790] | (layer_1[780] & layer_1[790]); 
    assign layer_2[781] = ~layer_1[781]; 
    assign layer_2[782] = 1'b1; 
    assign layer_2[783] = ~layer_1[798] | (layer_1[798] & layer_1[772]); 
    assign layer_2[784] = layer_1[788] & layer_1[780]; 
    assign layer_2[785] = layer_1[790] ^ layer_1[779]; 
    assign layer_2[786] = ~(layer_1[780] ^ layer_1[784]); 
    assign layer_2[787] = ~layer_1[781]; 
    assign layer_2[788] = ~layer_1[774]; 
    assign layer_2[789] = ~layer_1[772]; 
    assign layer_2[790] = layer_1[789]; 
    assign layer_2[791] = ~layer_1[801] | (layer_1[795] & layer_1[801]); 
    assign layer_2[792] = 1'b1; 
    assign layer_2[793] = ~(layer_1[781] ^ layer_1[801]); 
    assign layer_2[794] = ~layer_1[804] | (layer_1[804] & layer_1[795]); 
    assign layer_2[795] = layer_1[805]; 
    assign layer_2[796] = layer_1[787] ^ layer_1[789]; 
    assign layer_2[797] = ~layer_1[780]; 
    assign layer_2[798] = layer_1[806]; 
    assign layer_2[799] = layer_1[789] & ~layer_1[785]; 
    assign layer_2[800] = layer_1[788] | layer_1[795]; 
    assign layer_2[801] = ~layer_1[790]; 
    assign layer_2[802] = layer_1[798] | layer_1[807]; 
    assign layer_2[803] = 1'b0; 
    assign layer_2[804] = ~layer_1[805]; 
    assign layer_2[805] = ~(layer_1[805] ^ layer_1[815]); 
    assign layer_2[806] = layer_1[798] & ~layer_1[800]; 
    assign layer_2[807] = ~(layer_1[791] ^ layer_1[802]); 
    assign layer_2[808] = 1'b1; 
    assign layer_2[809] = ~(layer_1[794] ^ layer_1[797]); 
    assign layer_2[810] = layer_1[826]; 
    assign layer_2[811] = layer_1[818]; 
    assign layer_2[812] = layer_1[824] & ~layer_1[810]; 
    assign layer_2[813] = 1'b1; 
    assign layer_2[814] = layer_1[806] & layer_1[825]; 
    assign layer_2[815] = ~layer_1[812]; 
    assign layer_2[816] = 1'b0; 
    assign layer_2[817] = ~layer_1[826] | (layer_1[826] & layer_1[828]); 
    assign layer_2[818] = layer_1[826] & ~layer_1[818]; 
    assign layer_2[819] = layer_1[815] ^ layer_1[806]; 
    assign layer_2[820] = 1'b0; 
    assign layer_2[821] = ~(layer_1[830] & layer_1[821]); 
    assign layer_2[822] = ~layer_1[806] | (layer_1[838] & layer_1[806]); 
    assign layer_2[823] = layer_1[817]; 
    assign layer_2[824] = layer_1[827] | layer_1[821]; 
    assign layer_2[825] = ~(layer_1[827] | layer_1[831]); 
    assign layer_2[826] = layer_1[827] ^ layer_1[828]; 
    assign layer_2[827] = 1'b1; 
    assign layer_2[828] = ~layer_1[824]; 
    assign layer_2[829] = ~layer_1[819]; 
    assign layer_2[830] = 1'b1; 
    assign layer_2[831] = layer_1[844] ^ layer_1[833]; 
    assign layer_2[832] = ~layer_1[830] | (layer_1[843] & layer_1[830]); 
    assign layer_2[833] = 1'b0; 
    assign layer_2[834] = 1'b1; 
    assign layer_2[835] = ~layer_1[844] | (layer_1[839] & layer_1[844]); 
    assign layer_2[836] = ~layer_1[830]; 
    assign layer_2[837] = layer_1[848]; 
    assign layer_2[838] = ~(layer_1[839] & layer_1[845]); 
    assign layer_2[839] = ~layer_1[847]; 
    assign layer_2[840] = 1'b0; 
    assign layer_2[841] = 1'b0; 
    assign layer_2[842] = ~layer_1[831]; 
    assign layer_2[843] = layer_1[857] ^ layer_1[841]; 
    assign layer_2[844] = ~(layer_1[829] ^ layer_1[856]); 
    assign layer_2[845] = 1'b1; 
    assign layer_2[846] = layer_1[846]; 
    assign layer_2[847] = ~layer_1[836]; 
    assign layer_2[848] = ~layer_1[848]; 
    assign layer_2[849] = layer_1[855] & ~layer_1[842]; 
    assign layer_2[850] = layer_1[834] & ~layer_1[835]; 
    assign layer_2[851] = layer_1[857] | layer_1[860]; 
    assign layer_2[852] = ~layer_1[866] | (layer_1[866] & layer_1[860]); 
    assign layer_2[853] = 1'b0; 
    assign layer_2[854] = ~layer_1[848]; 
    assign layer_2[855] = layer_1[869] & ~layer_1[844]; 
    assign layer_2[856] = layer_1[859] ^ layer_1[850]; 
    assign layer_2[857] = ~(layer_1[872] ^ layer_1[868]); 
    assign layer_2[858] = 1'b0; 
    assign layer_2[859] = layer_1[871] & ~layer_1[848]; 
    assign layer_2[860] = layer_1[848] & layer_1[869]; 
    assign layer_2[861] = layer_1[865] ^ layer_1[859]; 
    assign layer_2[862] = layer_1[856] & ~layer_1[848]; 
    assign layer_2[863] = 1'b0; 
    assign layer_2[864] = 1'b0; 
    assign layer_2[865] = ~(layer_1[850] & layer_1[858]); 
    assign layer_2[866] = layer_1[859] ^ layer_1[864]; 
    assign layer_2[867] = ~layer_1[878] | (layer_1[855] & layer_1[878]); 
    assign layer_2[868] = ~(layer_1[866] | layer_1[881]); 
    assign layer_2[869] = layer_1[865]; 
    assign layer_2[870] = layer_1[886] & layer_1[878]; 
    assign layer_2[871] = ~layer_1[884]; 
    assign layer_2[872] = 1'b1; 
    assign layer_2[873] = ~(layer_1[874] & layer_1[887]); 
    assign layer_2[874] = ~layer_1[871]; 
    assign layer_2[875] = layer_1[870] & ~layer_1[859]; 
    assign layer_2[876] = ~layer_1[883]; 
    assign layer_2[877] = ~layer_1[890] | (layer_1[870] & layer_1[890]); 
    assign layer_2[878] = layer_1[864]; 
    assign layer_2[879] = ~layer_1[883]; 
    assign layer_2[880] = 1'b0; 
    assign layer_2[881] = ~(layer_1[869] | layer_1[881]); 
    assign layer_2[882] = 1'b0; 
    assign layer_2[883] = layer_1[867] & ~layer_1[871]; 
    assign layer_2[884] = ~layer_1[877] | (layer_1[893] & layer_1[877]); 
    assign layer_2[885] = layer_1[892] | layer_1[900]; 
    assign layer_2[886] = 1'b0; 
    assign layer_2[887] = ~(layer_1[885] | layer_1[887]); 
    assign layer_2[888] = ~layer_1[892]; 
    assign layer_2[889] = ~layer_1[901]; 
    assign layer_2[890] = ~(layer_1[902] ^ layer_1[883]); 
    assign layer_2[891] = ~layer_1[890]; 
    assign layer_2[892] = ~(layer_1[902] | layer_1[886]); 
    assign layer_2[893] = layer_1[892]; 
    assign layer_2[894] = ~layer_1[903]; 
    assign layer_2[895] = layer_1[891] & ~layer_1[882]; 
    assign layer_2[896] = 1'b0; 
    assign layer_2[897] = 1'b1; 
    assign layer_2[898] = ~layer_1[904]; 
    assign layer_2[899] = layer_1[906] & ~layer_1[895]; 
    assign layer_2[900] = ~layer_1[897]; 
    assign layer_2[901] = layer_1[907] & ~layer_1[893]; 
    assign layer_2[902] = layer_1[905] ^ layer_1[911]; 
    assign layer_2[903] = ~(layer_1[907] & layer_1[900]); 
    assign layer_2[904] = layer_1[888] & ~layer_1[891]; 
    assign layer_2[905] = ~layer_1[900] | (layer_1[906] & layer_1[900]); 
    assign layer_2[906] = layer_1[909] & layer_1[909]; 
    assign layer_2[907] = layer_1[918] & ~layer_1[902]; 
    assign layer_2[908] = layer_1[918] & ~layer_1[921]; 
    assign layer_2[909] = layer_1[917]; 
    assign layer_2[910] = 1'b1; 
    assign layer_2[911] = layer_1[926]; 
    assign layer_2[912] = ~layer_1[903] | (layer_1[903] & layer_1[905]); 
    assign layer_2[913] = layer_1[899] & ~layer_1[924]; 
    assign layer_2[914] = ~layer_1[903] | (layer_1[920] & layer_1[903]); 
    assign layer_2[915] = layer_1[919] ^ layer_1[926]; 
    assign layer_2[916] = ~layer_1[915] | (layer_1[932] & layer_1[915]); 
    assign layer_2[917] = layer_1[929] & layer_1[930]; 
    assign layer_2[918] = layer_1[926] | layer_1[904]; 
    assign layer_2[919] = ~layer_1[925] | (layer_1[923] & layer_1[925]); 
    assign layer_2[920] = ~(layer_1[917] ^ layer_1[903]); 
    assign layer_2[921] = layer_1[916]; 
    assign layer_2[922] = layer_1[918] ^ layer_1[919]; 
    assign layer_2[923] = ~layer_1[929] | (layer_1[919] & layer_1[929]); 
    assign layer_2[924] = ~layer_1[911]; 
    assign layer_2[925] = layer_1[936] ^ layer_1[932]; 
    assign layer_2[926] = layer_1[927] & ~layer_1[914]; 
    assign layer_2[927] = layer_1[913] & ~layer_1[924]; 
    assign layer_2[928] = 1'b1; 
    assign layer_2[929] = ~layer_1[924]; 
    assign layer_2[930] = ~layer_1[932]; 
    assign layer_2[931] = 1'b0; 
    assign layer_2[932] = layer_1[931] & ~layer_1[925]; 
    assign layer_2[933] = layer_1[921]; 
    assign layer_2[934] = layer_1[927] & ~layer_1[920]; 
    assign layer_2[935] = ~layer_1[942]; 
    assign layer_2[936] = ~(layer_1[921] ^ layer_1[929]); 
    assign layer_2[937] = ~(layer_1[921] | layer_1[920]); 
    assign layer_2[938] = ~layer_1[932]; 
    assign layer_2[939] = ~layer_1[929] | (layer_1[931] & layer_1[929]); 
    assign layer_2[940] = 1'b1; 
    assign layer_2[941] = ~layer_1[933]; 
    assign layer_2[942] = layer_1[953] & ~layer_1[943]; 
    assign layer_2[943] = layer_1[957] ^ layer_1[935]; 
    assign layer_2[944] = layer_1[932] & ~layer_1[932]; 
    assign layer_2[945] = ~(layer_1[953] | layer_1[941]); 
    assign layer_2[946] = layer_1[960] & layer_1[941]; 
    assign layer_2[947] = layer_1[958]; 
    assign layer_2[948] = layer_1[936]; 
    assign layer_2[949] = 1'b0; 
    assign layer_2[950] = layer_1[949]; 
    assign layer_2[951] = ~(layer_1[951] ^ layer_1[952]); 
    assign layer_2[952] = ~layer_1[953] | (layer_1[963] & layer_1[953]); 
    assign layer_2[953] = layer_1[948]; 
    assign layer_2[954] = ~(layer_1[967] | layer_1[968]); 
    assign layer_2[955] = 1'b1; 
    assign layer_2[956] = ~(layer_1[957] & layer_1[952]); 
    assign layer_2[957] = layer_1[965] ^ layer_1[949]; 
    assign layer_2[958] = layer_1[965] & ~layer_1[964]; 
    assign layer_2[959] = layer_1[964] & ~layer_1[970]; 
    assign layer_2[960] = layer_1[964] & ~layer_1[966]; 
    assign layer_2[961] = 1'b0; 
    assign layer_2[962] = layer_1[972] ^ layer_1[969]; 
    assign layer_2[963] = layer_1[965] & ~layer_1[958]; 
    assign layer_2[964] = layer_1[974] | layer_1[962]; 
    assign layer_2[965] = 1'b1; 
    assign layer_2[966] = ~layer_1[956]; 
    assign layer_2[967] = layer_1[981] & layer_1[979]; 
    assign layer_2[968] = ~layer_1[968]; 
    assign layer_2[969] = ~layer_1[984] | (layer_1[975] & layer_1[984]); 
    assign layer_2[970] = ~layer_1[961] | (layer_1[968] & layer_1[961]); 
    assign layer_2[971] = layer_1[959]; 
    assign layer_2[972] = ~layer_1[976]; 
    assign layer_2[973] = layer_1[968] & layer_1[979]; 
    assign layer_2[974] = ~(layer_1[965] | layer_1[962]); 
    assign layer_2[975] = ~layer_1[959] | (layer_1[959] & layer_1[962]); 
    assign layer_2[976] = 1'b1; 
    assign layer_2[977] = ~(layer_1[992] ^ layer_1[962]); 
    assign layer_2[978] = ~(layer_1[992] ^ layer_1[984]); 
    assign layer_2[979] = layer_1[985]; 
    assign layer_2[980] = ~layer_1[984] | (layer_1[984] & layer_1[971]); 
    assign layer_2[981] = layer_1[967] & layer_1[975]; 
    assign layer_2[982] = 1'b0; 
    assign layer_2[983] = ~(layer_1[972] ^ layer_1[977]); 
    assign layer_2[984] = layer_1[992] | layer_1[988]; 
    assign layer_2[985] = ~(layer_1[992] & layer_1[994]); 
    assign layer_2[986] = layer_1[995] & layer_1[974]; 
    assign layer_2[987] = ~(layer_1[996] & layer_1[974]); 
    assign layer_2[988] = layer_1[984] & ~layer_1[979]; 
    assign layer_2[989] = 1'b0; 
    assign layer_2[990] = 1'b1; 
    assign layer_2[991] = ~layer_1[996]; 
    assign layer_2[992] = layer_1[1007] | layer_1[1001]; 
    assign layer_2[993] = layer_1[1008] & layer_1[988]; 
    assign layer_2[994] = ~(layer_1[983] ^ layer_1[982]); 
    assign layer_2[995] = ~(layer_1[1002] ^ layer_1[1005]); 
    assign layer_2[996] = ~layer_1[1010]; 
    assign layer_2[997] = layer_1[984] ^ layer_1[998]; 
    assign layer_2[998] = layer_1[1003] ^ layer_1[1007]; 
    assign layer_2[999] = layer_1[986] | layer_1[991]; 
    assign layer_2[1000] = ~(layer_1[994] | layer_1[1005]); 
    assign layer_2[1001] = 1'b0; 
    assign layer_2[1002] = ~layer_1[1013]; 
    assign layer_2[1003] = 1'b1; 
    assign layer_2[1004] = layer_1[993] | layer_1[1015]; 
    assign layer_2[1005] = ~layer_1[1010] | (layer_1[1006] & layer_1[1010]); 
    assign layer_2[1006] = layer_1[995]; 
    assign layer_2[1007] = ~layer_1[992]; 
    assign layer_2[1008] = ~(layer_1[1003] ^ layer_1[1000]); 
    assign layer_2[1009] = layer_1[1022]; 
    assign layer_2[1010] = layer_1[995]; 
    assign layer_2[1011] = ~(layer_1[1001] | layer_1[1021]); 
    assign layer_2[1012] = layer_1[1017]; 
    assign layer_2[1013] = ~(layer_1[1013] | layer_1[1016]); 
    assign layer_2[1014] = ~layer_1[1013]; 
    assign layer_2[1015] = ~(layer_1[1009] & layer_1[1016]); 
    assign layer_2[1016] = layer_1[1007]; 
    assign layer_2[1017] = 1'b0; 
    assign layer_2[1018] = ~(layer_1[1012] | layer_1[1012]); 
    assign layer_2[1019] = layer_1[1018] & ~layer_1[1013]; 
    assign layer_2[1020] = ~layer_1[1013]; 
    assign layer_2[1021] = ~(layer_1[1011] ^ layer_1[1018]); 
    assign layer_2[1022] = layer_1[1007]; 
    assign layer_2[1023] = 1'b0; 
    // Layer 3 ============================================================
    assign layer_3[0] = layer_2[0] & ~layer_2[13]; 
    assign layer_3[1] = layer_2[3]; 
    assign layer_3[2] = layer_2[5]; 
    assign layer_3[3] = ~layer_2[5] | (layer_2[5] & layer_2[6]); 
    assign layer_3[4] = ~layer_2[2] | (layer_2[19] & layer_2[2]); 
    assign layer_3[5] = 1'b1; 
    assign layer_3[6] = ~layer_2[9] | (layer_2[9] & layer_2[7]); 
    assign layer_3[7] = 1'b0; 
    assign layer_3[8] = ~layer_2[20]; 
    assign layer_3[9] = layer_2[1]; 
    assign layer_3[10] = ~(layer_2[6] | layer_2[1]); 
    assign layer_3[11] = ~(layer_2[7] ^ layer_2[2]); 
    assign layer_3[12] = ~layer_2[26] | (layer_2[26] & layer_2[18]); 
    assign layer_3[13] = 1'b1; 
    assign layer_3[14] = ~layer_2[29]; 
    assign layer_3[15] = layer_2[4] & ~layer_2[28]; 
    assign layer_3[16] = ~(layer_2[6] | layer_2[15]); 
    assign layer_3[17] = ~layer_2[13]; 
    assign layer_3[18] = layer_2[16] & ~layer_2[12]; 
    assign layer_3[19] = ~(layer_2[3] & layer_2[18]); 
    assign layer_3[20] = ~layer_2[28] | (layer_2[34] & layer_2[28]); 
    assign layer_3[21] = ~layer_2[17]; 
    assign layer_3[22] = ~layer_2[13]; 
    assign layer_3[23] = ~layer_2[21] | (layer_2[21] & layer_2[28]); 
    assign layer_3[24] = ~layer_2[17]; 
    assign layer_3[25] = layer_2[9] & layer_2[15]; 
    assign layer_3[26] = ~layer_2[10]; 
    assign layer_3[27] = layer_2[15] & ~layer_2[15]; 
    assign layer_3[28] = layer_2[44] | layer_2[11]; 
    assign layer_3[29] = layer_2[23] & ~layer_2[24]; 
    assign layer_3[30] = layer_2[38] ^ layer_2[18]; 
    assign layer_3[31] = layer_2[28] & layer_2[20]; 
    assign layer_3[32] = ~layer_2[42]; 
    assign layer_3[33] = layer_2[17] | layer_2[26]; 
    assign layer_3[34] = layer_2[37] & ~layer_2[25]; 
    assign layer_3[35] = layer_2[50]; 
    assign layer_3[36] = ~layer_2[27] | (layer_2[24] & layer_2[27]); 
    assign layer_3[37] = ~(layer_2[33] | layer_2[23]); 
    assign layer_3[38] = layer_2[40]; 
    assign layer_3[39] = layer_2[45]; 
    assign layer_3[40] = ~layer_2[40]; 
    assign layer_3[41] = ~(layer_2[51] ^ layer_2[43]); 
    assign layer_3[42] = ~(layer_2[35] | layer_2[46]); 
    assign layer_3[43] = ~(layer_2[52] & layer_2[49]); 
    assign layer_3[44] = ~(layer_2[35] | layer_2[57]); 
    assign layer_3[45] = layer_2[38] | layer_2[58]; 
    assign layer_3[46] = layer_2[32]; 
    assign layer_3[47] = layer_2[48] | layer_2[57]; 
    assign layer_3[48] = layer_2[38] & ~layer_2[31]; 
    assign layer_3[49] = ~(layer_2[43] | layer_2[52]); 
    assign layer_3[50] = layer_2[40] & ~layer_2[52]; 
    assign layer_3[51] = 1'b0; 
    assign layer_3[52] = layer_2[59] & ~layer_2[47]; 
    assign layer_3[53] = layer_2[52] ^ layer_2[56]; 
    assign layer_3[54] = ~(layer_2[49] & layer_2[56]); 
    assign layer_3[55] = layer_2[71] & ~layer_2[54]; 
    assign layer_3[56] = layer_2[68] & layer_2[53]; 
    assign layer_3[57] = ~layer_2[56] | (layer_2[47] & layer_2[56]); 
    assign layer_3[58] = 1'b0; 
    assign layer_3[59] = ~layer_2[55]; 
    assign layer_3[60] = ~(layer_2[46] ^ layer_2[61]); 
    assign layer_3[61] = layer_2[64] ^ layer_2[53]; 
    assign layer_3[62] = ~(layer_2[78] | layer_2[46]); 
    assign layer_3[63] = layer_2[71] & ~layer_2[48]; 
    assign layer_3[64] = 1'b1; 
    assign layer_3[65] = 1'b1; 
    assign layer_3[66] = layer_2[80] & ~layer_2[60]; 
    assign layer_3[67] = ~layer_2[54] | (layer_2[54] & layer_2[52]); 
    assign layer_3[68] = ~(layer_2[84] | layer_2[53]); 
    assign layer_3[69] = layer_2[83] & layer_2[65]; 
    assign layer_3[70] = layer_2[77] ^ layer_2[66]; 
    assign layer_3[71] = ~layer_2[85]; 
    assign layer_3[72] = layer_2[80] | layer_2[61]; 
    assign layer_3[73] = layer_2[70]; 
    assign layer_3[74] = layer_2[71] & layer_2[72]; 
    assign layer_3[75] = layer_2[69] | layer_2[58]; 
    assign layer_3[76] = layer_2[82] & ~layer_2[74]; 
    assign layer_3[77] = ~(layer_2[77] ^ layer_2[69]); 
    assign layer_3[78] = ~layer_2[92]; 
    assign layer_3[79] = ~layer_2[68] | (layer_2[73] & layer_2[68]); 
    assign layer_3[80] = ~layer_2[83]; 
    assign layer_3[81] = ~(layer_2[81] | layer_2[88]); 
    assign layer_3[82] = 1'b0; 
    assign layer_3[83] = layer_2[97] & layer_2[70]; 
    assign layer_3[84] = ~(layer_2[70] & layer_2[74]); 
    assign layer_3[85] = ~(layer_2[91] & layer_2[82]); 
    assign layer_3[86] = ~(layer_2[95] ^ layer_2[76]); 
    assign layer_3[87] = layer_2[103] & ~layer_2[87]; 
    assign layer_3[88] = ~layer_2[92] | (layer_2[92] & layer_2[99]); 
    assign layer_3[89] = 1'b1; 
    assign layer_3[90] = layer_2[90] | layer_2[87]; 
    assign layer_3[91] = ~layer_2[105]; 
    assign layer_3[92] = layer_2[102]; 
    assign layer_3[93] = layer_2[102] | layer_2[88]; 
    assign layer_3[94] = layer_2[98] ^ layer_2[86]; 
    assign layer_3[95] = ~(layer_2[96] & layer_2[105]); 
    assign layer_3[96] = layer_2[112]; 
    assign layer_3[97] = ~layer_2[101]; 
    assign layer_3[98] = ~(layer_2[114] | layer_2[94]); 
    assign layer_3[99] = layer_2[88]; 
    assign layer_3[100] = ~layer_2[103] | (layer_2[103] & layer_2[89]); 
    assign layer_3[101] = layer_2[102] & ~layer_2[100]; 
    assign layer_3[102] = 1'b1; 
    assign layer_3[103] = ~(layer_2[105] ^ layer_2[118]); 
    assign layer_3[104] = layer_2[112] & ~layer_2[114]; 
    assign layer_3[105] = ~(layer_2[103] & layer_2[94]); 
    assign layer_3[106] = layer_2[119] & ~layer_2[111]; 
    assign layer_3[107] = ~(layer_2[116] & layer_2[122]); 
    assign layer_3[108] = layer_2[101] & layer_2[109]; 
    assign layer_3[109] = layer_2[105] & ~layer_2[114]; 
    assign layer_3[110] = layer_2[116] & ~layer_2[101]; 
    assign layer_3[111] = ~layer_2[95]; 
    assign layer_3[112] = ~layer_2[119]; 
    assign layer_3[113] = ~layer_2[111] | (layer_2[101] & layer_2[111]); 
    assign layer_3[114] = ~layer_2[129]; 
    assign layer_3[115] = ~layer_2[100]; 
    assign layer_3[116] = ~layer_2[110]; 
    assign layer_3[117] = layer_2[107]; 
    assign layer_3[118] = layer_2[133] ^ layer_2[124]; 
    assign layer_3[119] = layer_2[117]; 
    assign layer_3[120] = ~layer_2[128]; 
    assign layer_3[121] = ~(layer_2[118] ^ layer_2[131]); 
    assign layer_3[122] = ~layer_2[109]; 
    assign layer_3[123] = 1'b1; 
    assign layer_3[124] = ~(layer_2[134] ^ layer_2[113]); 
    assign layer_3[125] = 1'b0; 
    assign layer_3[126] = layer_2[118] | layer_2[134]; 
    assign layer_3[127] = layer_2[141]; 
    assign layer_3[128] = ~layer_2[115]; 
    assign layer_3[129] = ~(layer_2[113] | layer_2[127]); 
    assign layer_3[130] = 1'b0; 
    assign layer_3[131] = ~(layer_2[127] & layer_2[143]); 
    assign layer_3[132] = ~(layer_2[147] ^ layer_2[132]); 
    assign layer_3[133] = ~(layer_2[122] | layer_2[118]); 
    assign layer_3[134] = layer_2[133]; 
    assign layer_3[135] = ~(layer_2[121] ^ layer_2[131]); 
    assign layer_3[136] = layer_2[152] & ~layer_2[127]; 
    assign layer_3[137] = layer_2[126] & ~layer_2[142]; 
    assign layer_3[138] = layer_2[123] & layer_2[144]; 
    assign layer_3[139] = ~(layer_2[124] ^ layer_2[144]); 
    assign layer_3[140] = layer_2[135] ^ layer_2[139]; 
    assign layer_3[141] = ~(layer_2[154] & layer_2[153]); 
    assign layer_3[142] = layer_2[127] & layer_2[132]; 
    assign layer_3[143] = ~(layer_2[128] & layer_2[148]); 
    assign layer_3[144] = layer_2[135] & ~layer_2[151]; 
    assign layer_3[145] = ~layer_2[149] | (layer_2[149] & layer_2[145]); 
    assign layer_3[146] = layer_2[151] & ~layer_2[159]; 
    assign layer_3[147] = layer_2[152] | layer_2[134]; 
    assign layer_3[148] = layer_2[155] & ~layer_2[141]; 
    assign layer_3[149] = layer_2[161]; 
    assign layer_3[150] = ~(layer_2[141] | layer_2[133]); 
    assign layer_3[151] = layer_2[150] | layer_2[151]; 
    assign layer_3[152] = layer_2[141] & layer_2[141]; 
    assign layer_3[153] = layer_2[151] & ~layer_2[141]; 
    assign layer_3[154] = layer_2[170] ^ layer_2[157]; 
    assign layer_3[155] = layer_2[167] & ~layer_2[148]; 
    assign layer_3[156] = layer_2[155] ^ layer_2[156]; 
    assign layer_3[157] = layer_2[161]; 
    assign layer_3[158] = ~layer_2[163] | (layer_2[163] & layer_2[166]); 
    assign layer_3[159] = ~(layer_2[153] | layer_2[148]); 
    assign layer_3[160] = layer_2[170] | layer_2[156]; 
    assign layer_3[161] = ~(layer_2[152] | layer_2[156]); 
    assign layer_3[162] = 1'b0; 
    assign layer_3[163] = ~layer_2[155]; 
    assign layer_3[164] = layer_2[153] & ~layer_2[176]; 
    assign layer_3[165] = layer_2[177]; 
    assign layer_3[166] = ~layer_2[152] | (layer_2[154] & layer_2[152]); 
    assign layer_3[167] = layer_2[169] & layer_2[151]; 
    assign layer_3[168] = ~(layer_2[156] | layer_2[182]); 
    assign layer_3[169] = ~(layer_2[168] ^ layer_2[162]); 
    assign layer_3[170] = layer_2[174] & ~layer_2[182]; 
    assign layer_3[171] = layer_2[167] ^ layer_2[157]; 
    assign layer_3[172] = layer_2[184]; 
    assign layer_3[173] = ~layer_2[177] | (layer_2[177] & layer_2[173]); 
    assign layer_3[174] = layer_2[159] & layer_2[180]; 
    assign layer_3[175] = layer_2[180] & layer_2[164]; 
    assign layer_3[176] = 1'b0; 
    assign layer_3[177] = layer_2[192] & layer_2[173]; 
    assign layer_3[178] = layer_2[162] & ~layer_2[163]; 
    assign layer_3[179] = layer_2[163] | layer_2[183]; 
    assign layer_3[180] = 1'b1; 
    assign layer_3[181] = ~(layer_2[167] ^ layer_2[174]); 
    assign layer_3[182] = layer_2[180] & ~layer_2[165]; 
    assign layer_3[183] = layer_2[193]; 
    assign layer_3[184] = ~layer_2[185]; 
    assign layer_3[185] = layer_2[170]; 
    assign layer_3[186] = layer_2[191] | layer_2[177]; 
    assign layer_3[187] = layer_2[190] & ~layer_2[195]; 
    assign layer_3[188] = ~layer_2[183] | (layer_2[198] & layer_2[183]); 
    assign layer_3[189] = ~(layer_2[198] ^ layer_2[183]); 
    assign layer_3[190] = ~layer_2[205]; 
    assign layer_3[191] = ~layer_2[206] | (layer_2[191] & layer_2[206]); 
    assign layer_3[192] = layer_2[188] & ~layer_2[183]; 
    assign layer_3[193] = ~layer_2[186]; 
    assign layer_3[194] = layer_2[203] & layer_2[192]; 
    assign layer_3[195] = ~(layer_2[192] & layer_2[208]); 
    assign layer_3[196] = layer_2[189] & layer_2[205]; 
    assign layer_3[197] = 1'b0; 
    assign layer_3[198] = layer_2[200] & layer_2[195]; 
    assign layer_3[199] = layer_2[212] & ~layer_2[193]; 
    assign layer_3[200] = layer_2[198]; 
    assign layer_3[201] = layer_2[208] | layer_2[198]; 
    assign layer_3[202] = layer_2[190] & ~layer_2[211]; 
    assign layer_3[203] = layer_2[210] & ~layer_2[216]; 
    assign layer_3[204] = layer_2[187] & ~layer_2[216]; 
    assign layer_3[205] = ~(layer_2[213] & layer_2[203]); 
    assign layer_3[206] = layer_2[202]; 
    assign layer_3[207] = layer_2[208]; 
    assign layer_3[208] = ~(layer_2[201] ^ layer_2[191]); 
    assign layer_3[209] = ~layer_2[219]; 
    assign layer_3[210] = ~(layer_2[226] ^ layer_2[208]); 
    assign layer_3[211] = ~layer_2[206] | (layer_2[216] & layer_2[206]); 
    assign layer_3[212] = layer_2[221] & layer_2[209]; 
    assign layer_3[213] = layer_2[225] & ~layer_2[224]; 
    assign layer_3[214] = layer_2[208] & layer_2[217]; 
    assign layer_3[215] = ~(layer_2[219] & layer_2[227]); 
    assign layer_3[216] = ~layer_2[222]; 
    assign layer_3[217] = ~layer_2[219] | (layer_2[219] & layer_2[229]); 
    assign layer_3[218] = ~(layer_2[223] & layer_2[225]); 
    assign layer_3[219] = layer_2[229]; 
    assign layer_3[220] = layer_2[216] & ~layer_2[214]; 
    assign layer_3[221] = 1'b1; 
    assign layer_3[222] = layer_2[206] & ~layer_2[221]; 
    assign layer_3[223] = ~layer_2[228] | (layer_2[228] & layer_2[211]); 
    assign layer_3[224] = ~(layer_2[215] ^ layer_2[213]); 
    assign layer_3[225] = layer_2[214] & layer_2[227]; 
    assign layer_3[226] = layer_2[228] & ~layer_2[241]; 
    assign layer_3[227] = ~layer_2[227]; 
    assign layer_3[228] = ~(layer_2[237] & layer_2[239]); 
    assign layer_3[229] = 1'b0; 
    assign layer_3[230] = layer_2[230] & ~layer_2[236]; 
    assign layer_3[231] = ~layer_2[233] | (layer_2[233] & layer_2[216]); 
    assign layer_3[232] = layer_2[220]; 
    assign layer_3[233] = 1'b1; 
    assign layer_3[234] = ~layer_2[225]; 
    assign layer_3[235] = ~layer_2[230] | (layer_2[246] & layer_2[230]); 
    assign layer_3[236] = 1'b1; 
    assign layer_3[237] = ~(layer_2[249] ^ layer_2[247]); 
    assign layer_3[238] = layer_2[243] & ~layer_2[222]; 
    assign layer_3[239] = ~layer_2[240] | (layer_2[223] & layer_2[240]); 
    assign layer_3[240] = ~(layer_2[251] & layer_2[226]); 
    assign layer_3[241] = ~(layer_2[252] | layer_2[238]); 
    assign layer_3[242] = layer_2[245] & ~layer_2[236]; 
    assign layer_3[243] = 1'b1; 
    assign layer_3[244] = layer_2[254] & ~layer_2[245]; 
    assign layer_3[245] = layer_2[261] & layer_2[233]; 
    assign layer_3[246] = ~layer_2[231]; 
    assign layer_3[247] = ~layer_2[241]; 
    assign layer_3[248] = layer_2[255]; 
    assign layer_3[249] = 1'b1; 
    assign layer_3[250] = ~(layer_2[244] ^ layer_2[242]); 
    assign layer_3[251] = ~layer_2[249]; 
    assign layer_3[252] = ~layer_2[260]; 
    assign layer_3[253] = ~(layer_2[238] | layer_2[253]); 
    assign layer_3[254] = ~(layer_2[240] & layer_2[250]); 
    assign layer_3[255] = ~(layer_2[241] | layer_2[255]); 
    assign layer_3[256] = ~(layer_2[269] & layer_2[253]); 
    assign layer_3[257] = 1'b0; 
    assign layer_3[258] = ~(layer_2[245] ^ layer_2[273]); 
    assign layer_3[259] = layer_2[268] ^ layer_2[261]; 
    assign layer_3[260] = ~layer_2[275]; 
    assign layer_3[261] = ~(layer_2[256] & layer_2[248]); 
    assign layer_3[262] = layer_2[276] ^ layer_2[266]; 
    assign layer_3[263] = layer_2[275] ^ layer_2[250]; 
    assign layer_3[264] = layer_2[277] & layer_2[279]; 
    assign layer_3[265] = ~layer_2[249] | (layer_2[280] & layer_2[249]); 
    assign layer_3[266] = 1'b1; 
    assign layer_3[267] = layer_2[260] | layer_2[266]; 
    assign layer_3[268] = ~(layer_2[276] | layer_2[281]); 
    assign layer_3[269] = ~layer_2[283]; 
    assign layer_3[270] = ~layer_2[270]; 
    assign layer_3[271] = ~layer_2[259] | (layer_2[259] & layer_2[264]); 
    assign layer_3[272] = layer_2[280] | layer_2[266]; 
    assign layer_3[273] = ~layer_2[286] | (layer_2[286] & layer_2[276]); 
    assign layer_3[274] = layer_2[271]; 
    assign layer_3[275] = layer_2[276] & ~layer_2[275]; 
    assign layer_3[276] = layer_2[291] & layer_2[260]; 
    assign layer_3[277] = ~layer_2[293]; 
    assign layer_3[278] = layer_2[271] & layer_2[272]; 
    assign layer_3[279] = ~layer_2[287]; 
    assign layer_3[280] = ~layer_2[286]; 
    assign layer_3[281] = 1'b1; 
    assign layer_3[282] = 1'b1; 
    assign layer_3[283] = layer_2[294]; 
    assign layer_3[284] = layer_2[274]; 
    assign layer_3[285] = layer_2[276]; 
    assign layer_3[286] = ~layer_2[302]; 
    assign layer_3[287] = ~layer_2[279]; 
    assign layer_3[288] = ~layer_2[298] | (layer_2[298] & layer_2[271]); 
    assign layer_3[289] = ~(layer_2[290] ^ layer_2[302]); 
    assign layer_3[290] = 1'b0; 
    assign layer_3[291] = ~(layer_2[294] ^ layer_2[293]); 
    assign layer_3[292] = 1'b0; 
    assign layer_3[293] = ~layer_2[285] | (layer_2[306] & layer_2[285]); 
    assign layer_3[294] = ~(layer_2[292] | layer_2[293]); 
    assign layer_3[295] = 1'b1; 
    assign layer_3[296] = ~layer_2[305]; 
    assign layer_3[297] = ~layer_2[306] | (layer_2[306] & layer_2[285]); 
    assign layer_3[298] = layer_2[302]; 
    assign layer_3[299] = 1'b1; 
    assign layer_3[300] = ~layer_2[312]; 
    assign layer_3[301] = layer_2[291] & layer_2[293]; 
    assign layer_3[302] = ~layer_2[286] | (layer_2[293] & layer_2[286]); 
    assign layer_3[303] = layer_2[297]; 
    assign layer_3[304] = layer_2[291] & ~layer_2[313]; 
    assign layer_3[305] = layer_2[311] ^ layer_2[291]; 
    assign layer_3[306] = ~(layer_2[298] | layer_2[297]); 
    assign layer_3[307] = 1'b1; 
    assign layer_3[308] = layer_2[315] & ~layer_2[292]; 
    assign layer_3[309] = layer_2[304] & ~layer_2[300]; 
    assign layer_3[310] = ~(layer_2[296] | layer_2[324]); 
    assign layer_3[311] = ~(layer_2[299] & layer_2[317]); 
    assign layer_3[312] = layer_2[298] & ~layer_2[309]; 
    assign layer_3[313] = layer_2[316]; 
    assign layer_3[314] = 1'b0; 
    assign layer_3[315] = layer_2[310] & layer_2[320]; 
    assign layer_3[316] = layer_2[324] | layer_2[313]; 
    assign layer_3[317] = ~layer_2[314]; 
    assign layer_3[318] = ~layer_2[333] | (layer_2[334] & layer_2[333]); 
    assign layer_3[319] = ~layer_2[318]; 
    assign layer_3[320] = ~(layer_2[310] ^ layer_2[333]); 
    assign layer_3[321] = ~layer_2[309] | (layer_2[332] & layer_2[309]); 
    assign layer_3[322] = ~layer_2[312]; 
    assign layer_3[323] = layer_2[308] & layer_2[329]; 
    assign layer_3[324] = layer_2[315] & ~layer_2[334]; 
    assign layer_3[325] = 1'b1; 
    assign layer_3[326] = ~(layer_2[330] & layer_2[321]); 
    assign layer_3[327] = layer_2[319] ^ layer_2[339]; 
    assign layer_3[328] = ~layer_2[340] | (layer_2[334] & layer_2[340]); 
    assign layer_3[329] = ~layer_2[314]; 
    assign layer_3[330] = 1'b1; 
    assign layer_3[331] = ~layer_2[321]; 
    assign layer_3[332] = ~(layer_2[316] & layer_2[343]); 
    assign layer_3[333] = ~layer_2[339] | (layer_2[339] & layer_2[328]); 
    assign layer_3[334] = layer_2[325] & ~layer_2[347]; 
    assign layer_3[335] = layer_2[342] & layer_2[319]; 
    assign layer_3[336] = ~(layer_2[351] & layer_2[321]); 
    assign layer_3[337] = layer_2[351] & layer_2[349]; 
    assign layer_3[338] = layer_2[339] & layer_2[329]; 
    assign layer_3[339] = layer_2[348]; 
    assign layer_3[340] = layer_2[356] & ~layer_2[343]; 
    assign layer_3[341] = layer_2[325] & ~layer_2[329]; 
    assign layer_3[342] = ~(layer_2[348] ^ layer_2[325]); 
    assign layer_3[343] = layer_2[335] ^ layer_2[336]; 
    assign layer_3[344] = ~layer_2[343]; 
    assign layer_3[345] = ~layer_2[351] | (layer_2[333] & layer_2[351]); 
    assign layer_3[346] = ~(layer_2[348] ^ layer_2[353]); 
    assign layer_3[347] = ~layer_2[357]; 
    assign layer_3[348] = ~layer_2[344] | (layer_2[344] & layer_2[347]); 
    assign layer_3[349] = layer_2[340] & layer_2[335]; 
    assign layer_3[350] = 1'b0; 
    assign layer_3[351] = layer_2[339]; 
    assign layer_3[352] = ~layer_2[354] | (layer_2[354] & layer_2[367]); 
    assign layer_3[353] = 1'b0; 
    assign layer_3[354] = ~layer_2[363] | (layer_2[350] & layer_2[363]); 
    assign layer_3[355] = layer_2[363] ^ layer_2[346]; 
    assign layer_3[356] = layer_2[353] & ~layer_2[353]; 
    assign layer_3[357] = ~layer_2[365]; 
    assign layer_3[358] = layer_2[359]; 
    assign layer_3[359] = ~layer_2[361]; 
    assign layer_3[360] = ~layer_2[350]; 
    assign layer_3[361] = ~(layer_2[372] & layer_2[361]); 
    assign layer_3[362] = layer_2[351]; 
    assign layer_3[363] = layer_2[348]; 
    assign layer_3[364] = 1'b1; 
    assign layer_3[365] = layer_2[379] ^ layer_2[350]; 
    assign layer_3[366] = 1'b1; 
    assign layer_3[367] = layer_2[379]; 
    assign layer_3[368] = ~(layer_2[373] & layer_2[356]); 
    assign layer_3[369] = ~layer_2[357]; 
    assign layer_3[370] = layer_2[368] & ~layer_2[365]; 
    assign layer_3[371] = layer_2[386] & ~layer_2[359]; 
    assign layer_3[372] = layer_2[359] & ~layer_2[365]; 
    assign layer_3[373] = layer_2[378] & layer_2[360]; 
    assign layer_3[374] = layer_2[388] & layer_2[370]; 
    assign layer_3[375] = ~layer_2[379]; 
    assign layer_3[376] = layer_2[368]; 
    assign layer_3[377] = ~layer_2[374]; 
    assign layer_3[378] = ~(layer_2[375] ^ layer_2[378]); 
    assign layer_3[379] = ~layer_2[374]; 
    assign layer_3[380] = 1'b0; 
    assign layer_3[381] = 1'b0; 
    assign layer_3[382] = layer_2[375]; 
    assign layer_3[383] = 1'b1; 
    assign layer_3[384] = ~(layer_2[379] & layer_2[396]); 
    assign layer_3[385] = layer_2[390] | layer_2[376]; 
    assign layer_3[386] = layer_2[389] ^ layer_2[375]; 
    assign layer_3[387] = layer_2[376] & ~layer_2[374]; 
    assign layer_3[388] = ~(layer_2[403] | layer_2[388]); 
    assign layer_3[389] = layer_2[403] & layer_2[388]; 
    assign layer_3[390] = ~layer_2[385]; 
    assign layer_3[391] = layer_2[376] ^ layer_2[399]; 
    assign layer_3[392] = layer_2[377] | layer_2[380]; 
    assign layer_3[393] = 1'b1; 
    assign layer_3[394] = ~(layer_2[408] ^ layer_2[404]); 
    assign layer_3[395] = ~(layer_2[406] ^ layer_2[399]); 
    assign layer_3[396] = ~layer_2[385]; 
    assign layer_3[397] = ~(layer_2[411] ^ layer_2[391]); 
    assign layer_3[398] = layer_2[399] & layer_2[406]; 
    assign layer_3[399] = ~layer_2[403]; 
    assign layer_3[400] = ~layer_2[397] | (layer_2[397] & layer_2[407]); 
    assign layer_3[401] = layer_2[400]; 
    assign layer_3[402] = ~(layer_2[405] ^ layer_2[393]); 
    assign layer_3[403] = layer_2[412] & ~layer_2[387]; 
    assign layer_3[404] = layer_2[418] | layer_2[387]; 
    assign layer_3[405] = 1'b1; 
    assign layer_3[406] = ~layer_2[414] | (layer_2[414] & layer_2[419]); 
    assign layer_3[407] = 1'b1; 
    assign layer_3[408] = layer_2[405] | layer_2[405]; 
    assign layer_3[409] = ~layer_2[424]; 
    assign layer_3[410] = layer_2[405]; 
    assign layer_3[411] = ~(layer_2[411] ^ layer_2[407]); 
    assign layer_3[412] = layer_2[404] & layer_2[425]; 
    assign layer_3[413] = layer_2[398] & ~layer_2[402]; 
    assign layer_3[414] = layer_2[400] ^ layer_2[420]; 
    assign layer_3[415] = ~layer_2[417] | (layer_2[429] & layer_2[417]); 
    assign layer_3[416] = layer_2[401]; 
    assign layer_3[417] = ~layer_2[420] | (layer_2[420] & layer_2[401]); 
    assign layer_3[418] = layer_2[427]; 
    assign layer_3[419] = layer_2[403] & layer_2[422]; 
    assign layer_3[420] = ~layer_2[421] | (layer_2[421] & layer_2[431]); 
    assign layer_3[421] = ~layer_2[424] | (layer_2[424] & layer_2[422]); 
    assign layer_3[422] = ~layer_2[419]; 
    assign layer_3[423] = ~layer_2[415] | (layer_2[407] & layer_2[415]); 
    assign layer_3[424] = layer_2[431]; 
    assign layer_3[425] = 1'b1; 
    assign layer_3[426] = layer_2[420]; 
    assign layer_3[427] = layer_2[431]; 
    assign layer_3[428] = ~(layer_2[415] & layer_2[415]); 
    assign layer_3[429] = ~layer_2[424]; 
    assign layer_3[430] = ~(layer_2[420] ^ layer_2[428]); 
    assign layer_3[431] = 1'b0; 
    assign layer_3[432] = layer_2[436] & ~layer_2[435]; 
    assign layer_3[433] = ~layer_2[437]; 
    assign layer_3[434] = ~layer_2[439] | (layer_2[438] & layer_2[439]); 
    assign layer_3[435] = layer_2[423] & layer_2[428]; 
    assign layer_3[436] = ~layer_2[430] | (layer_2[430] & layer_2[429]); 
    assign layer_3[437] = layer_2[444]; 
    assign layer_3[438] = 1'b1; 
    assign layer_3[439] = ~layer_2[431]; 
    assign layer_3[440] = layer_2[440] ^ layer_2[444]; 
    assign layer_3[441] = ~layer_2[452]; 
    assign layer_3[442] = ~(layer_2[450] | layer_2[426]); 
    assign layer_3[443] = layer_2[458]; 
    assign layer_3[444] = ~(layer_2[446] & layer_2[432]); 
    assign layer_3[445] = 1'b1; 
    assign layer_3[446] = layer_2[431] & ~layer_2[460]; 
    assign layer_3[447] = 1'b0; 
    assign layer_3[448] = layer_2[449]; 
    assign layer_3[449] = layer_2[443] & ~layer_2[445]; 
    assign layer_3[450] = ~layer_2[444]; 
    assign layer_3[451] = 1'b0; 
    assign layer_3[452] = ~layer_2[451] | (layer_2[451] & layer_2[440]); 
    assign layer_3[453] = layer_2[456] | layer_2[449]; 
    assign layer_3[454] = layer_2[448] & ~layer_2[443]; 
    assign layer_3[455] = layer_2[458]; 
    assign layer_3[456] = 1'b1; 
    assign layer_3[457] = ~layer_2[441]; 
    assign layer_3[458] = ~layer_2[450]; 
    assign layer_3[459] = ~layer_2[471] | (layer_2[468] & layer_2[471]); 
    assign layer_3[460] = ~(layer_2[446] ^ layer_2[451]); 
    assign layer_3[461] = layer_2[461] & ~layer_2[459]; 
    assign layer_3[462] = ~layer_2[472]; 
    assign layer_3[463] = layer_2[474]; 
    assign layer_3[464] = layer_2[473] & layer_2[473]; 
    assign layer_3[465] = layer_2[448] & ~layer_2[468]; 
    assign layer_3[466] = ~layer_2[454]; 
    assign layer_3[467] = ~layer_2[471] | (layer_2[471] & layer_2[460]); 
    assign layer_3[468] = layer_2[457] ^ layer_2[464]; 
    assign layer_3[469] = ~(layer_2[462] & layer_2[472]); 
    assign layer_3[470] = ~(layer_2[486] & layer_2[472]); 
    assign layer_3[471] = layer_2[463] | layer_2[465]; 
    assign layer_3[472] = layer_2[474]; 
    assign layer_3[473] = ~layer_2[477] | (layer_2[477] & layer_2[460]); 
    assign layer_3[474] = ~layer_2[470]; 
    assign layer_3[475] = layer_2[460] & ~layer_2[484]; 
    assign layer_3[476] = 1'b0; 
    assign layer_3[477] = layer_2[482] & ~layer_2[491]; 
    assign layer_3[478] = layer_2[478] | layer_2[481]; 
    assign layer_3[479] = 1'b1; 
    assign layer_3[480] = 1'b1; 
    assign layer_3[481] = ~layer_2[486] | (layer_2[490] & layer_2[486]); 
    assign layer_3[482] = layer_2[467]; 
    assign layer_3[483] = layer_2[475] | layer_2[475]; 
    assign layer_3[484] = ~layer_2[495] | (layer_2[487] & layer_2[495]); 
    assign layer_3[485] = ~layer_2[483] | (layer_2[483] & layer_2[474]); 
    assign layer_3[486] = layer_2[490] & ~layer_2[477]; 
    assign layer_3[487] = 1'b0; 
    assign layer_3[488] = layer_2[499] & ~layer_2[474]; 
    assign layer_3[489] = 1'b0; 
    assign layer_3[490] = ~layer_2[474] | (layer_2[474] & layer_2[491]); 
    assign layer_3[491] = ~(layer_2[478] ^ layer_2[495]); 
    assign layer_3[492] = layer_2[479] ^ layer_2[478]; 
    assign layer_3[493] = ~(layer_2[485] | layer_2[485]); 
    assign layer_3[494] = ~(layer_2[507] & layer_2[488]); 
    assign layer_3[495] = layer_2[494] ^ layer_2[481]; 
    assign layer_3[496] = layer_2[486] | layer_2[508]; 
    assign layer_3[497] = layer_2[482]; 
    assign layer_3[498] = layer_2[495] | layer_2[502]; 
    assign layer_3[499] = layer_2[491]; 
    assign layer_3[500] = layer_2[494]; 
    assign layer_3[501] = ~(layer_2[508] | layer_2[512]); 
    assign layer_3[502] = layer_2[507] & layer_2[516]; 
    assign layer_3[503] = 1'b0; 
    assign layer_3[504] = ~layer_2[512] | (layer_2[512] & layer_2[510]); 
    assign layer_3[505] = layer_2[517]; 
    assign layer_3[506] = ~layer_2[504]; 
    assign layer_3[507] = ~layer_2[492] | (layer_2[492] & layer_2[500]); 
    assign layer_3[508] = layer_2[521]; 
    assign layer_3[509] = layer_2[518] & ~layer_2[524]; 
    assign layer_3[510] = layer_2[495]; 
    assign layer_3[511] = ~layer_2[513] | (layer_2[496] & layer_2[513]); 
    assign layer_3[512] = 1'b0; 
    assign layer_3[513] = layer_2[497] & ~layer_2[522]; 
    assign layer_3[514] = layer_2[514] & ~layer_2[522]; 
    assign layer_3[515] = layer_2[520] | layer_2[508]; 
    assign layer_3[516] = layer_2[528] & ~layer_2[501]; 
    assign layer_3[517] = 1'b0; 
    assign layer_3[518] = layer_2[526] & ~layer_2[512]; 
    assign layer_3[519] = ~(layer_2[519] & layer_2[530]); 
    assign layer_3[520] = 1'b0; 
    assign layer_3[521] = ~(layer_2[524] & layer_2[505]); 
    assign layer_3[522] = ~(layer_2[530] | layer_2[529]); 
    assign layer_3[523] = layer_2[523] & ~layer_2[510]; 
    assign layer_3[524] = ~(layer_2[529] | layer_2[539]); 
    assign layer_3[525] = layer_2[510] & ~layer_2[516]; 
    assign layer_3[526] = layer_2[517]; 
    assign layer_3[527] = layer_2[533] | layer_2[516]; 
    assign layer_3[528] = ~layer_2[531]; 
    assign layer_3[529] = layer_2[529] & ~layer_2[515]; 
    assign layer_3[530] = ~(layer_2[529] & layer_2[531]); 
    assign layer_3[531] = layer_2[524] & ~layer_2[524]; 
    assign layer_3[532] = layer_2[539] & ~layer_2[538]; 
    assign layer_3[533] = layer_2[547] & layer_2[534]; 
    assign layer_3[534] = layer_2[528] & layer_2[525]; 
    assign layer_3[535] = layer_2[519] ^ layer_2[544]; 
    assign layer_3[536] = ~(layer_2[535] | layer_2[522]); 
    assign layer_3[537] = ~(layer_2[545] ^ layer_2[552]); 
    assign layer_3[538] = 1'b0; 
    assign layer_3[539] = ~layer_2[534] | (layer_2[534] & layer_2[552]); 
    assign layer_3[540] = 1'b1; 
    assign layer_3[541] = ~layer_2[556]; 
    assign layer_3[542] = layer_2[556] & ~layer_2[542]; 
    assign layer_3[543] = layer_2[548]; 
    assign layer_3[544] = ~layer_2[529] | (layer_2[529] & layer_2[558]); 
    assign layer_3[545] = ~layer_2[542]; 
    assign layer_3[546] = ~layer_2[554]; 
    assign layer_3[547] = 1'b0; 
    assign layer_3[548] = layer_2[547] ^ layer_2[559]; 
    assign layer_3[549] = layer_2[548] ^ layer_2[553]; 
    assign layer_3[550] = ~layer_2[549] | (layer_2[549] & layer_2[539]); 
    assign layer_3[551] = layer_2[548]; 
    assign layer_3[552] = layer_2[560] & ~layer_2[542]; 
    assign layer_3[553] = 1'b0; 
    assign layer_3[554] = layer_2[539] & ~layer_2[540]; 
    assign layer_3[555] = 1'b0; 
    assign layer_3[556] = 1'b0; 
    assign layer_3[557] = layer_2[544] & ~layer_2[568]; 
    assign layer_3[558] = layer_2[569] & layer_2[550]; 
    assign layer_3[559] = ~(layer_2[554] & layer_2[546]); 
    assign layer_3[560] = ~layer_2[557] | (layer_2[565] & layer_2[557]); 
    assign layer_3[561] = layer_2[567] & layer_2[570]; 
    assign layer_3[562] = ~(layer_2[567] & layer_2[546]); 
    assign layer_3[563] = ~layer_2[554] | (layer_2[554] & layer_2[574]); 
    assign layer_3[564] = ~layer_2[558]; 
    assign layer_3[565] = layer_2[552]; 
    assign layer_3[566] = ~layer_2[556]; 
    assign layer_3[567] = 1'b1; 
    assign layer_3[568] = ~layer_2[575] | (layer_2[575] & layer_2[567]); 
    assign layer_3[569] = ~(layer_2[564] & layer_2[573]); 
    assign layer_3[570] = layer_2[554] ^ layer_2[556]; 
    assign layer_3[571] = ~layer_2[567] | (layer_2[567] & layer_2[573]); 
    assign layer_3[572] = 1'b1; 
    assign layer_3[573] = ~layer_2[572]; 
    assign layer_3[574] = ~layer_2[587]; 
    assign layer_3[575] = ~(layer_2[589] | layer_2[579]); 
    assign layer_3[576] = ~layer_2[577]; 
    assign layer_3[577] = layer_2[561] & ~layer_2[575]; 
    assign layer_3[578] = ~(layer_2[580] ^ layer_2[593]); 
    assign layer_3[579] = layer_2[580] & layer_2[590]; 
    assign layer_3[580] = ~(layer_2[579] & layer_2[569]); 
    assign layer_3[581] = ~(layer_2[595] | layer_2[589]); 
    assign layer_3[582] = ~(layer_2[576] & layer_2[577]); 
    assign layer_3[583] = 1'b1; 
    assign layer_3[584] = ~(layer_2[595] & layer_2[597]); 
    assign layer_3[585] = ~(layer_2[573] | layer_2[599]); 
    assign layer_3[586] = ~layer_2[584] | (layer_2[584] & layer_2[584]); 
    assign layer_3[587] = ~(layer_2[595] & layer_2[602]); 
    assign layer_3[588] = ~layer_2[597]; 
    assign layer_3[589] = ~layer_2[602] | (layer_2[577] & layer_2[602]); 
    assign layer_3[590] = ~(layer_2[578] & layer_2[602]); 
    assign layer_3[591] = ~(layer_2[595] ^ layer_2[584]); 
    assign layer_3[592] = layer_2[605] & layer_2[591]; 
    assign layer_3[593] = ~(layer_2[607] & layer_2[584]); 
    assign layer_3[594] = ~(layer_2[578] | layer_2[586]); 
    assign layer_3[595] = ~layer_2[583] | (layer_2[579] & layer_2[583]); 
    assign layer_3[596] = 1'b0; 
    assign layer_3[597] = ~(layer_2[591] ^ layer_2[584]); 
    assign layer_3[598] = ~layer_2[595]; 
    assign layer_3[599] = 1'b1; 
    assign layer_3[600] = 1'b0; 
    assign layer_3[601] = ~layer_2[611]; 
    assign layer_3[602] = 1'b0; 
    assign layer_3[603] = ~(layer_2[597] & layer_2[590]); 
    assign layer_3[604] = ~(layer_2[590] ^ layer_2[607]); 
    assign layer_3[605] = ~layer_2[591]; 
    assign layer_3[606] = 1'b1; 
    assign layer_3[607] = layer_2[621]; 
    assign layer_3[608] = layer_2[602] ^ layer_2[617]; 
    assign layer_3[609] = ~layer_2[622] | (layer_2[604] & layer_2[622]); 
    assign layer_3[610] = layer_2[607] ^ layer_2[601]; 
    assign layer_3[611] = layer_2[609] & ~layer_2[615]; 
    assign layer_3[612] = 1'b0; 
    assign layer_3[613] = layer_2[617] & ~layer_2[616]; 
    assign layer_3[614] = 1'b0; 
    assign layer_3[615] = layer_2[627] & ~layer_2[598]; 
    assign layer_3[616] = ~(layer_2[605] ^ layer_2[628]); 
    assign layer_3[617] = ~(layer_2[607] ^ layer_2[607]); 
    assign layer_3[618] = ~layer_2[611]; 
    assign layer_3[619] = ~layer_2[608] | (layer_2[615] & layer_2[608]); 
    assign layer_3[620] = ~layer_2[623] | (layer_2[623] & layer_2[617]); 
    assign layer_3[621] = layer_2[614]; 
    assign layer_3[622] = ~(layer_2[635] ^ layer_2[622]); 
    assign layer_3[623] = ~(layer_2[627] & layer_2[631]); 
    assign layer_3[624] = layer_2[608]; 
    assign layer_3[625] = layer_2[626]; 
    assign layer_3[626] = ~layer_2[611]; 
    assign layer_3[627] = 1'b1; 
    assign layer_3[628] = ~(layer_2[623] | layer_2[634]); 
    assign layer_3[629] = layer_2[616] & ~layer_2[616]; 
    assign layer_3[630] = layer_2[623] & layer_2[640]; 
    assign layer_3[631] = layer_2[643] & ~layer_2[635]; 
    assign layer_3[632] = 1'b0; 
    assign layer_3[633] = 1'b1; 
    assign layer_3[634] = layer_2[634] | layer_2[633]; 
    assign layer_3[635] = layer_2[628] & ~layer_2[626]; 
    assign layer_3[636] = ~(layer_2[629] ^ layer_2[635]); 
    assign layer_3[637] = layer_2[628] | layer_2[636]; 
    assign layer_3[638] = layer_2[645] & ~layer_2[652]; 
    assign layer_3[639] = layer_2[643] | layer_2[633]; 
    assign layer_3[640] = layer_2[651] & layer_2[637]; 
    assign layer_3[641] = layer_2[656] ^ layer_2[643]; 
    assign layer_3[642] = ~layer_2[648]; 
    assign layer_3[643] = ~layer_2[641] | (layer_2[641] & layer_2[638]); 
    assign layer_3[644] = layer_2[646] ^ layer_2[659]; 
    assign layer_3[645] = ~(layer_2[659] | layer_2[636]); 
    assign layer_3[646] = ~layer_2[631]; 
    assign layer_3[647] = layer_2[643]; 
    assign layer_3[648] = ~layer_2[655]; 
    assign layer_3[649] = layer_2[634] ^ layer_2[654]; 
    assign layer_3[650] = layer_2[647] & ~layer_2[664]; 
    assign layer_3[651] = ~(layer_2[640] | layer_2[644]); 
    assign layer_3[652] = 1'b1; 
    assign layer_3[653] = ~(layer_2[649] ^ layer_2[667]); 
    assign layer_3[654] = 1'b1; 
    assign layer_3[655] = ~(layer_2[640] | layer_2[659]); 
    assign layer_3[656] = 1'b1; 
    assign layer_3[657] = ~(layer_2[641] ^ layer_2[672]); 
    assign layer_3[658] = layer_2[672]; 
    assign layer_3[659] = 1'b1; 
    assign layer_3[660] = layer_2[660] ^ layer_2[661]; 
    assign layer_3[661] = ~layer_2[655]; 
    assign layer_3[662] = layer_2[656]; 
    assign layer_3[663] = layer_2[663] ^ layer_2[670]; 
    assign layer_3[664] = ~layer_2[672] | (layer_2[670] & layer_2[672]); 
    assign layer_3[665] = ~(layer_2[659] ^ layer_2[670]); 
    assign layer_3[666] = ~layer_2[659] | (layer_2[659] & layer_2[650]); 
    assign layer_3[667] = 1'b1; 
    assign layer_3[668] = layer_2[670]; 
    assign layer_3[669] = layer_2[660] & ~layer_2[673]; 
    assign layer_3[670] = layer_2[682] & ~layer_2[671]; 
    assign layer_3[671] = layer_2[659] & layer_2[674]; 
    assign layer_3[672] = layer_2[678]; 
    assign layer_3[673] = 1'b1; 
    assign layer_3[674] = layer_2[666] | layer_2[674]; 
    assign layer_3[675] = layer_2[659] & ~layer_2[658]; 
    assign layer_3[676] = ~layer_2[663] | (layer_2[663] & layer_2[690]); 
    assign layer_3[677] = ~layer_2[668] | (layer_2[665] & layer_2[668]); 
    assign layer_3[678] = layer_2[675] & ~layer_2[691]; 
    assign layer_3[679] = layer_2[674] & ~layer_2[691]; 
    assign layer_3[680] = ~layer_2[675] | (layer_2[675] & layer_2[682]); 
    assign layer_3[681] = ~(layer_2[667] & layer_2[686]); 
    assign layer_3[682] = 1'b0; 
    assign layer_3[683] = 1'b0; 
    assign layer_3[684] = ~layer_2[668]; 
    assign layer_3[685] = ~(layer_2[697] ^ layer_2[689]); 
    assign layer_3[686] = layer_2[688]; 
    assign layer_3[687] = layer_2[691] ^ layer_2[673]; 
    assign layer_3[688] = 1'b0; 
    assign layer_3[689] = layer_2[686] ^ layer_2[690]; 
    assign layer_3[690] = 1'b1; 
    assign layer_3[691] = layer_2[691] & layer_2[698]; 
    assign layer_3[692] = 1'b1; 
    assign layer_3[693] = ~(layer_2[679] ^ layer_2[684]); 
    assign layer_3[694] = ~layer_2[702] | (layer_2[702] & layer_2[689]); 
    assign layer_3[695] = layer_2[708] & ~layer_2[690]; 
    assign layer_3[696] = 1'b0; 
    assign layer_3[697] = ~layer_2[703]; 
    assign layer_3[698] = layer_2[701] | layer_2[697]; 
    assign layer_3[699] = ~layer_2[707] | (layer_2[707] & layer_2[712]); 
    assign layer_3[700] = ~layer_2[716]; 
    assign layer_3[701] = layer_2[692] ^ layer_2[692]; 
    assign layer_3[702] = layer_2[712] | layer_2[686]; 
    assign layer_3[703] = ~(layer_2[707] & layer_2[705]); 
    assign layer_3[704] = layer_2[689]; 
    assign layer_3[705] = ~layer_2[691] | (layer_2[711] & layer_2[691]); 
    assign layer_3[706] = 1'b1; 
    assign layer_3[707] = ~(layer_2[707] ^ layer_2[701]); 
    assign layer_3[708] = 1'b0; 
    assign layer_3[709] = ~layer_2[704] | (layer_2[704] & layer_2[722]); 
    assign layer_3[710] = layer_2[710] & ~layer_2[707]; 
    assign layer_3[711] = layer_2[706]; 
    assign layer_3[712] = ~layer_2[709] | (layer_2[708] & layer_2[709]); 
    assign layer_3[713] = ~(layer_2[710] | layer_2[726]); 
    assign layer_3[714] = layer_2[715]; 
    assign layer_3[715] = layer_2[707] | layer_2[723]; 
    assign layer_3[716] = ~layer_2[710] | (layer_2[710] & layer_2[724]); 
    assign layer_3[717] = layer_2[723] & layer_2[727]; 
    assign layer_3[718] = ~(layer_2[709] & layer_2[723]); 
    assign layer_3[719] = ~(layer_2[705] | layer_2[729]); 
    assign layer_3[720] = layer_2[718] & ~layer_2[716]; 
    assign layer_3[721] = 1'b0; 
    assign layer_3[722] = ~layer_2[711]; 
    assign layer_3[723] = 1'b1; 
    assign layer_3[724] = 1'b1; 
    assign layer_3[725] = ~layer_2[724] | (layer_2[724] & layer_2[713]); 
    assign layer_3[726] = layer_2[725]; 
    assign layer_3[727] = ~(layer_2[730] & layer_2[735]); 
    assign layer_3[728] = layer_2[734] ^ layer_2[731]; 
    assign layer_3[729] = 1'b0; 
    assign layer_3[730] = layer_2[718]; 
    assign layer_3[731] = ~layer_2[730]; 
    assign layer_3[732] = ~(layer_2[735] | layer_2[741]); 
    assign layer_3[733] = ~(layer_2[740] & layer_2[745]); 
    assign layer_3[734] = ~layer_2[722] | (layer_2[739] & layer_2[722]); 
    assign layer_3[735] = ~layer_2[733]; 
    assign layer_3[736] = 1'b1; 
    assign layer_3[737] = 1'b0; 
    assign layer_3[738] = layer_2[749]; 
    assign layer_3[739] = layer_2[734] & ~layer_2[724]; 
    assign layer_3[740] = ~(layer_2[732] | layer_2[752]); 
    assign layer_3[741] = 1'b1; 
    assign layer_3[742] = ~layer_2[744] | (layer_2[729] & layer_2[744]); 
    assign layer_3[743] = ~(layer_2[734] | layer_2[743]); 
    assign layer_3[744] = layer_2[737] & ~layer_2[731]; 
    assign layer_3[745] = ~(layer_2[737] | layer_2[753]); 
    assign layer_3[746] = ~layer_2[735] | (layer_2[736] & layer_2[735]); 
    assign layer_3[747] = ~(layer_2[739] ^ layer_2[732]); 
    assign layer_3[748] = layer_2[743] & layer_2[739]; 
    assign layer_3[749] = layer_2[758] & ~layer_2[745]; 
    assign layer_3[750] = layer_2[749] ^ layer_2[737]; 
    assign layer_3[751] = ~layer_2[736]; 
    assign layer_3[752] = layer_2[751] & ~layer_2[756]; 
    assign layer_3[753] = ~(layer_2[766] ^ layer_2[743]); 
    assign layer_3[754] = 1'b1; 
    assign layer_3[755] = ~layer_2[763] | (layer_2[763] & layer_2[746]); 
    assign layer_3[756] = layer_2[742] | layer_2[741]; 
    assign layer_3[757] = layer_2[742] & ~layer_2[752]; 
    assign layer_3[758] = ~layer_2[773]; 
    assign layer_3[759] = ~layer_2[760] | (layer_2[746] & layer_2[760]); 
    assign layer_3[760] = ~layer_2[763]; 
    assign layer_3[761] = 1'b1; 
    assign layer_3[762] = ~(layer_2[760] & layer_2[748]); 
    assign layer_3[763] = layer_2[750]; 
    assign layer_3[764] = layer_2[754] & ~layer_2[767]; 
    assign layer_3[765] = layer_2[774] & ~layer_2[769]; 
    assign layer_3[766] = ~layer_2[766]; 
    assign layer_3[767] = ~(layer_2[781] ^ layer_2[765]); 
    assign layer_3[768] = ~layer_2[775]; 
    assign layer_3[769] = ~(layer_2[770] & layer_2[778]); 
    assign layer_3[770] = layer_2[777] & layer_2[761]; 
    assign layer_3[771] = layer_2[768] & ~layer_2[781]; 
    assign layer_3[772] = ~layer_2[766]; 
    assign layer_3[773] = layer_2[779] ^ layer_2[781]; 
    assign layer_3[774] = layer_2[759] & ~layer_2[788]; 
    assign layer_3[775] = ~(layer_2[764] & layer_2[787]); 
    assign layer_3[776] = ~(layer_2[791] & layer_2[772]); 
    assign layer_3[777] = layer_2[783] | layer_2[769]; 
    assign layer_3[778] = ~layer_2[776] | (layer_2[776] & layer_2[780]); 
    assign layer_3[779] = 1'b1; 
    assign layer_3[780] = ~layer_2[784] | (layer_2[784] & layer_2[774]); 
    assign layer_3[781] = ~layer_2[773] | (layer_2[777] & layer_2[773]); 
    assign layer_3[782] = layer_2[775]; 
    assign layer_3[783] = layer_2[767]; 
    assign layer_3[784] = ~(layer_2[788] ^ layer_2[772]); 
    assign layer_3[785] = ~layer_2[786] | (layer_2[800] & layer_2[786]); 
    assign layer_3[786] = 1'b1; 
    assign layer_3[787] = layer_2[777] ^ layer_2[799]; 
    assign layer_3[788] = ~layer_2[782] | (layer_2[782] & layer_2[772]); 
    assign layer_3[789] = ~(layer_2[775] ^ layer_2[791]); 
    assign layer_3[790] = ~layer_2[800]; 
    assign layer_3[791] = 1'b1; 
    assign layer_3[792] = ~layer_2[802] | (layer_2[782] & layer_2[802]); 
    assign layer_3[793] = 1'b1; 
    assign layer_3[794] = layer_2[804] ^ layer_2[788]; 
    assign layer_3[795] = ~layer_2[787] | (layer_2[787] & layer_2[784]); 
    assign layer_3[796] = layer_2[804] & ~layer_2[810]; 
    assign layer_3[797] = ~layer_2[799] | (layer_2[802] & layer_2[799]); 
    assign layer_3[798] = layer_2[801] & ~layer_2[797]; 
    assign layer_3[799] = layer_2[790] ^ layer_2[804]; 
    assign layer_3[800] = ~layer_2[809]; 
    assign layer_3[801] = ~layer_2[786] | (layer_2[796] & layer_2[786]); 
    assign layer_3[802] = layer_2[801] | layer_2[812]; 
    assign layer_3[803] = ~(layer_2[801] & layer_2[809]); 
    assign layer_3[804] = 1'b1; 
    assign layer_3[805] = 1'b1; 
    assign layer_3[806] = ~(layer_2[805] | layer_2[814]); 
    assign layer_3[807] = layer_2[822] & ~layer_2[803]; 
    assign layer_3[808] = ~layer_2[805] | (layer_2[805] & layer_2[794]); 
    assign layer_3[809] = 1'b0; 
    assign layer_3[810] = ~layer_2[826] | (layer_2[826] & layer_2[812]); 
    assign layer_3[811] = layer_2[816] & layer_2[813]; 
    assign layer_3[812] = layer_2[817] & ~layer_2[803]; 
    assign layer_3[813] = layer_2[824] ^ layer_2[803]; 
    assign layer_3[814] = ~(layer_2[798] | layer_2[814]); 
    assign layer_3[815] = ~layer_2[826]; 
    assign layer_3[816] = layer_2[805] & ~layer_2[809]; 
    assign layer_3[817] = layer_2[809] & ~layer_2[804]; 
    assign layer_3[818] = ~(layer_2[819] ^ layer_2[821]); 
    assign layer_3[819] = ~(layer_2[816] | layer_2[827]); 
    assign layer_3[820] = 1'b0; 
    assign layer_3[821] = layer_2[805] | layer_2[829]; 
    assign layer_3[822] = ~(layer_2[820] | layer_2[825]); 
    assign layer_3[823] = layer_2[831] & ~layer_2[835]; 
    assign layer_3[824] = ~(layer_2[822] | layer_2[815]); 
    assign layer_3[825] = ~layer_2[822] | (layer_2[821] & layer_2[822]); 
    assign layer_3[826] = layer_2[840]; 
    assign layer_3[827] = ~layer_2[819]; 
    assign layer_3[828] = ~layer_2[838]; 
    assign layer_3[829] = ~(layer_2[841] & layer_2[838]); 
    assign layer_3[830] = ~layer_2[814] | (layer_2[814] & layer_2[828]); 
    assign layer_3[831] = layer_2[819]; 
    assign layer_3[832] = layer_2[830]; 
    assign layer_3[833] = ~(layer_2[818] & layer_2[821]); 
    assign layer_3[834] = layer_2[819] | layer_2[843]; 
    assign layer_3[835] = layer_2[823] | layer_2[850]; 
    assign layer_3[836] = layer_2[831] ^ layer_2[849]; 
    assign layer_3[837] = ~layer_2[839] | (layer_2[850] & layer_2[839]); 
    assign layer_3[838] = layer_2[822] | layer_2[850]; 
    assign layer_3[839] = layer_2[833] | layer_2[854]; 
    assign layer_3[840] = layer_2[826] & ~layer_2[845]; 
    assign layer_3[841] = layer_2[855] ^ layer_2[824]; 
    assign layer_3[842] = 1'b0; 
    assign layer_3[843] = layer_2[846]; 
    assign layer_3[844] = ~layer_2[853] | (layer_2[854] & layer_2[853]); 
    assign layer_3[845] = layer_2[852] ^ layer_2[845]; 
    assign layer_3[846] = ~(layer_2[835] & layer_2[850]); 
    assign layer_3[847] = ~layer_2[860]; 
    assign layer_3[848] = ~layer_2[861] | (layer_2[864] & layer_2[861]); 
    assign layer_3[849] = ~layer_2[864] | (layer_2[864] & layer_2[841]); 
    assign layer_3[850] = ~layer_2[864]; 
    assign layer_3[851] = layer_2[836]; 
    assign layer_3[852] = layer_2[847] & ~layer_2[836]; 
    assign layer_3[853] = ~layer_2[855] | (layer_2[853] & layer_2[855]); 
    assign layer_3[854] = layer_2[843] & ~layer_2[861]; 
    assign layer_3[855] = layer_2[866] & ~layer_2[854]; 
    assign layer_3[856] = layer_2[851] | layer_2[869]; 
    assign layer_3[857] = 1'b1; 
    assign layer_3[858] = layer_2[843]; 
    assign layer_3[859] = 1'b1; 
    assign layer_3[860] = ~(layer_2[858] | layer_2[866]); 
    assign layer_3[861] = ~layer_2[873]; 
    assign layer_3[862] = ~layer_2[866]; 
    assign layer_3[863] = ~layer_2[847]; 
    assign layer_3[864] = 1'b1; 
    assign layer_3[865] = layer_2[850] & ~layer_2[864]; 
    assign layer_3[866] = layer_2[876] & ~layer_2[864]; 
    assign layer_3[867] = 1'b1; 
    assign layer_3[868] = layer_2[861] ^ layer_2[868]; 
    assign layer_3[869] = layer_2[879] & layer_2[874]; 
    assign layer_3[870] = layer_2[856] | layer_2[869]; 
    assign layer_3[871] = ~layer_2[871]; 
    assign layer_3[872] = ~layer_2[857]; 
    assign layer_3[873] = 1'b1; 
    assign layer_3[874] = layer_2[888] | layer_2[859]; 
    assign layer_3[875] = layer_2[864] & ~layer_2[889]; 
    assign layer_3[876] = ~layer_2[861] | (layer_2[872] & layer_2[861]); 
    assign layer_3[877] = ~layer_2[873]; 
    assign layer_3[878] = layer_2[881]; 
    assign layer_3[879] = layer_2[866]; 
    assign layer_3[880] = ~(layer_2[871] & layer_2[881]); 
    assign layer_3[881] = 1'b1; 
    assign layer_3[882] = ~(layer_2[867] | layer_2[887]); 
    assign layer_3[883] = ~(layer_2[867] ^ layer_2[875]); 
    assign layer_3[884] = ~(layer_2[885] & layer_2[898]); 
    assign layer_3[885] = ~(layer_2[897] & layer_2[878]); 
    assign layer_3[886] = ~layer_2[876]; 
    assign layer_3[887] = 1'b1; 
    assign layer_3[888] = 1'b0; 
    assign layer_3[889] = ~layer_2[897]; 
    assign layer_3[890] = ~(layer_2[877] | layer_2[890]); 
    assign layer_3[891] = layer_2[878] | layer_2[883]; 
    assign layer_3[892] = ~layer_2[877] | (layer_2[905] & layer_2[877]); 
    assign layer_3[893] = ~layer_2[909]; 
    assign layer_3[894] = 1'b1; 
    assign layer_3[895] = layer_2[893] & ~layer_2[894]; 
    assign layer_3[896] = ~layer_2[900] | (layer_2[900] & layer_2[884]); 
    assign layer_3[897] = ~(layer_2[908] & layer_2[905]); 
    assign layer_3[898] = ~layer_2[885] | (layer_2[885] & layer_2[884]); 
    assign layer_3[899] = layer_2[914] & layer_2[903]; 
    assign layer_3[900] = ~(layer_2[901] | layer_2[897]); 
    assign layer_3[901] = 1'b1; 
    assign layer_3[902] = layer_2[892] ^ layer_2[900]; 
    assign layer_3[903] = ~(layer_2[906] | layer_2[905]); 
    assign layer_3[904] = layer_2[903] & ~layer_2[893]; 
    assign layer_3[905] = ~(layer_2[895] ^ layer_2[890]); 
    assign layer_3[906] = layer_2[922] & layer_2[892]; 
    assign layer_3[907] = 1'b1; 
    assign layer_3[908] = layer_2[899] | layer_2[900]; 
    assign layer_3[909] = ~layer_2[922] | (layer_2[922] & layer_2[920]); 
    assign layer_3[910] = layer_2[919]; 
    assign layer_3[911] = layer_2[915]; 
    assign layer_3[912] = 1'b1; 
    assign layer_3[913] = layer_2[899] & ~layer_2[924]; 
    assign layer_3[914] = ~(layer_2[917] | layer_2[898]); 
    assign layer_3[915] = layer_2[911] & ~layer_2[923]; 
    assign layer_3[916] = ~layer_2[931]; 
    assign layer_3[917] = layer_2[931] & ~layer_2[918]; 
    assign layer_3[918] = ~(layer_2[903] & layer_2[932]); 
    assign layer_3[919] = ~(layer_2[906] | layer_2[931]); 
    assign layer_3[920] = layer_2[919] | layer_2[910]; 
    assign layer_3[921] = ~(layer_2[932] & layer_2[924]); 
    assign layer_3[922] = ~layer_2[912] | (layer_2[912] & layer_2[924]); 
    assign layer_3[923] = layer_2[909] & ~layer_2[910]; 
    assign layer_3[924] = ~layer_2[915] | (layer_2[920] & layer_2[915]); 
    assign layer_3[925] = ~layer_2[924]; 
    assign layer_3[926] = 1'b1; 
    assign layer_3[927] = layer_2[926]; 
    assign layer_3[928] = ~layer_2[912] | (layer_2[940] & layer_2[912]); 
    assign layer_3[929] = layer_2[920] & layer_2[918]; 
    assign layer_3[930] = ~layer_2[944]; 
    assign layer_3[931] = ~layer_2[919]; 
    assign layer_3[932] = ~(layer_2[946] & layer_2[941]); 
    assign layer_3[933] = layer_2[945]; 
    assign layer_3[934] = ~(layer_2[943] ^ layer_2[936]); 
    assign layer_3[935] = ~(layer_2[929] & layer_2[948]); 
    assign layer_3[936] = ~layer_2[932]; 
    assign layer_3[937] = layer_2[943]; 
    assign layer_3[938] = layer_2[939]; 
    assign layer_3[939] = ~layer_2[943]; 
    assign layer_3[940] = layer_2[938] | layer_2[950]; 
    assign layer_3[941] = ~(layer_2[930] ^ layer_2[954]); 
    assign layer_3[942] = ~layer_2[932]; 
    assign layer_3[943] = ~(layer_2[934] | layer_2[926]); 
    assign layer_3[944] = ~layer_2[955] | (layer_2[940] & layer_2[955]); 
    assign layer_3[945] = layer_2[944] ^ layer_2[931]; 
    assign layer_3[946] = layer_2[934] & ~layer_2[960]; 
    assign layer_3[947] = layer_2[952]; 
    assign layer_3[948] = ~(layer_2[934] | layer_2[949]); 
    assign layer_3[949] = 1'b0; 
    assign layer_3[950] = layer_2[952]; 
    assign layer_3[951] = layer_2[937] ^ layer_2[952]; 
    assign layer_3[952] = 1'b0; 
    assign layer_3[953] = layer_2[957] & layer_2[948]; 
    assign layer_3[954] = 1'b1; 
    assign layer_3[955] = layer_2[970]; 
    assign layer_3[956] = ~layer_2[959] | (layer_2[948] & layer_2[959]); 
    assign layer_3[957] = layer_2[965] | layer_2[971]; 
    assign layer_3[958] = 1'b1; 
    assign layer_3[959] = layer_2[974] | layer_2[955]; 
    assign layer_3[960] = ~layer_2[949]; 
    assign layer_3[961] = layer_2[948]; 
    assign layer_3[962] = 1'b1; 
    assign layer_3[963] = layer_2[967]; 
    assign layer_3[964] = ~layer_2[966] | (layer_2[975] & layer_2[966]); 
    assign layer_3[965] = ~(layer_2[960] ^ layer_2[975]); 
    assign layer_3[966] = layer_2[972] & ~layer_2[957]; 
    assign layer_3[967] = ~(layer_2[982] ^ layer_2[954]); 
    assign layer_3[968] = layer_2[970] & ~layer_2[958]; 
    assign layer_3[969] = ~layer_2[957] | (layer_2[967] & layer_2[957]); 
    assign layer_3[970] = ~layer_2[973] | (layer_2[973] & layer_2[968]); 
    assign layer_3[971] = layer_2[978] & ~layer_2[968]; 
    assign layer_3[972] = ~(layer_2[979] | layer_2[968]); 
    assign layer_3[973] = layer_2[956]; 
    assign layer_3[974] = layer_2[971] ^ layer_2[981]; 
    assign layer_3[975] = ~layer_2[965] | (layer_2[965] & layer_2[979]); 
    assign layer_3[976] = ~layer_2[970] | (layer_2[986] & layer_2[970]); 
    assign layer_3[977] = layer_2[972] ^ layer_2[982]; 
    assign layer_3[978] = layer_2[973] | layer_2[968]; 
    assign layer_3[979] = layer_2[982] & ~layer_2[977]; 
    assign layer_3[980] = ~(layer_2[974] ^ layer_2[986]); 
    assign layer_3[981] = ~(layer_2[974] ^ layer_2[985]); 
    assign layer_3[982] = ~layer_2[974]; 
    assign layer_3[983] = ~(layer_2[994] | layer_2[983]); 
    assign layer_3[984] = layer_2[994]; 
    assign layer_3[985] = ~layer_2[970] | (layer_2[970] & layer_2[986]); 
    assign layer_3[986] = layer_2[996] | layer_2[985]; 
    assign layer_3[987] = layer_2[975]; 
    assign layer_3[988] = ~(layer_2[998] ^ layer_2[988]); 
    assign layer_3[989] = ~(layer_2[973] | layer_2[991]); 
    assign layer_3[990] = layer_2[980] & ~layer_2[977]; 
    assign layer_3[991] = ~layer_2[997] | (layer_2[997] & layer_2[976]); 
    assign layer_3[992] = layer_2[1002] ^ layer_2[991]; 
    assign layer_3[993] = ~layer_2[1006]; 
    assign layer_3[994] = 1'b1; 
    assign layer_3[995] = layer_2[997] & ~layer_2[998]; 
    assign layer_3[996] = ~(layer_2[992] | layer_2[1000]); 
    assign layer_3[997] = ~(layer_2[993] & layer_2[1002]); 
    assign layer_3[998] = ~layer_2[1008]; 
    assign layer_3[999] = ~layer_2[1012]; 
    assign layer_3[1000] = layer_2[997]; 
    assign layer_3[1001] = ~layer_2[998] | (layer_2[1010] & layer_2[998]); 
    assign layer_3[1002] = layer_2[994] ^ layer_2[1005]; 
    assign layer_3[1003] = ~layer_2[1003]; 
    assign layer_3[1004] = ~(layer_2[1010] & layer_2[996]); 
    assign layer_3[1005] = layer_2[993]; 
    assign layer_3[1006] = layer_2[996]; 
    assign layer_3[1007] = layer_2[1020]; 
    assign layer_3[1008] = ~(layer_2[1012] & layer_2[993]); 
    assign layer_3[1009] = 1'b0; 
    assign layer_3[1010] = layer_2[1022]; 
    assign layer_3[1011] = ~layer_2[1008] | (layer_2[1008] & layer_2[1022]); 
    assign layer_3[1012] = 1'b1; 
    assign layer_3[1013] = ~layer_2[1006] | (layer_2[1006] & layer_2[1009]); 
    assign layer_3[1014] = layer_2[1001] | layer_2[1018]; 
    assign layer_3[1015] = ~layer_2[1003]; 
    assign layer_3[1016] = 1'b0; 
    assign layer_3[1017] = ~layer_2[1021]; 
    assign layer_3[1018] = 1'b0; 
    assign layer_3[1019] = 1'b0; 
    assign layer_3[1020] = layer_2[1021]; 
    assign layer_3[1021] = 1'b0; 
    assign layer_3[1022] = 1'b1; 
    assign layer_3[1023] = layer_2[1015] & layer_2[1017]; 
    // Layer 4 ============================================================
    assign layer_4[0] = ~layer_3[13] | (layer_3[13] & layer_3[3]); 
    assign layer_4[1] = ~layer_3[7]; 
    assign layer_4[2] = layer_3[6] & ~layer_3[1]; 
    assign layer_4[3] = layer_3[17] | layer_3[3]; 
    assign layer_4[4] = layer_3[2] | layer_3[4]; 
    assign layer_4[5] = layer_3[13]; 
    assign layer_4[6] = 1'b1; 
    assign layer_4[7] = layer_3[18]; 
    assign layer_4[8] = ~layer_3[14]; 
    assign layer_4[9] = ~(layer_3[4] | layer_3[6]); 
    assign layer_4[10] = ~layer_3[4]; 
    assign layer_4[11] = layer_3[20]; 
    assign layer_4[12] = ~layer_3[9] | (layer_3[21] & layer_3[9]); 
    assign layer_4[13] = ~(layer_3[18] & layer_3[14]); 
    assign layer_4[14] = ~(layer_3[16] ^ layer_3[7]); 
    assign layer_4[15] = 1'b0; 
    assign layer_4[16] = layer_3[25] & ~layer_3[2]; 
    assign layer_4[17] = 1'b1; 
    assign layer_4[18] = layer_3[19] & layer_3[26]; 
    assign layer_4[19] = 1'b1; 
    assign layer_4[20] = ~layer_3[12]; 
    assign layer_4[21] = layer_3[12] & layer_3[13]; 
    assign layer_4[22] = layer_3[28]; 
    assign layer_4[23] = layer_3[31]; 
    assign layer_4[24] = ~(layer_3[29] & layer_3[8]); 
    assign layer_4[25] = layer_3[12]; 
    assign layer_4[26] = layer_3[40] | layer_3[19]; 
    assign layer_4[27] = 1'b0; 
    assign layer_4[28] = ~layer_3[21] | (layer_3[16] & layer_3[21]); 
    assign layer_4[29] = ~(layer_3[30] & layer_3[33]); 
    assign layer_4[30] = layer_3[16] ^ layer_3[15]; 
    assign layer_4[31] = layer_3[26] & ~layer_3[43]; 
    assign layer_4[32] = layer_3[46]; 
    assign layer_4[33] = ~(layer_3[24] | layer_3[35]); 
    assign layer_4[34] = layer_3[27] ^ layer_3[35]; 
    assign layer_4[35] = ~layer_3[22] | (layer_3[45] & layer_3[22]); 
    assign layer_4[36] = layer_3[41] & layer_3[48]; 
    assign layer_4[37] = layer_3[40] & ~layer_3[39]; 
    assign layer_4[38] = ~layer_3[24] | (layer_3[24] & layer_3[42]); 
    assign layer_4[39] = layer_3[53] ^ layer_3[26]; 
    assign layer_4[40] = layer_3[41]; 
    assign layer_4[41] = ~(layer_3[32] ^ layer_3[55]); 
    assign layer_4[42] = ~layer_3[46] | (layer_3[41] & layer_3[46]); 
    assign layer_4[43] = layer_3[57] & ~layer_3[31]; 
    assign layer_4[44] = ~(layer_3[44] | layer_3[28]); 
    assign layer_4[45] = 1'b1; 
    assign layer_4[46] = 1'b1; 
    assign layer_4[47] = ~layer_3[60]; 
    assign layer_4[48] = layer_3[34] ^ layer_3[47]; 
    assign layer_4[49] = 1'b1; 
    assign layer_4[50] = layer_3[38]; 
    assign layer_4[51] = ~(layer_3[59] | layer_3[54]); 
    assign layer_4[52] = ~layer_3[45]; 
    assign layer_4[53] = ~(layer_3[37] ^ layer_3[52]); 
    assign layer_4[54] = layer_3[37]; 
    assign layer_4[55] = 1'b1; 
    assign layer_4[56] = ~(layer_3[58] & layer_3[61]); 
    assign layer_4[57] = layer_3[57] & ~layer_3[54]; 
    assign layer_4[58] = layer_3[71]; 
    assign layer_4[59] = layer_3[53]; 
    assign layer_4[60] = ~layer_3[58] | (layer_3[58] & layer_3[43]); 
    assign layer_4[61] = ~(layer_3[57] ^ layer_3[50]); 
    assign layer_4[62] = ~(layer_3[55] & layer_3[68]); 
    assign layer_4[63] = layer_3[68] ^ layer_3[65]; 
    assign layer_4[64] = layer_3[72]; 
    assign layer_4[65] = layer_3[64]; 
    assign layer_4[66] = 1'b1; 
    assign layer_4[67] = 1'b0; 
    assign layer_4[68] = ~layer_3[79] | (layer_3[72] & layer_3[79]); 
    assign layer_4[69] = ~layer_3[56]; 
    assign layer_4[70] = layer_3[80] & ~layer_3[57]; 
    assign layer_4[71] = layer_3[86]; 
    assign layer_4[72] = layer_3[66] & layer_3[65]; 
    assign layer_4[73] = layer_3[87]; 
    assign layer_4[74] = ~layer_3[87]; 
    assign layer_4[75] = layer_3[72] & ~layer_3[89]; 
    assign layer_4[76] = ~layer_3[63] | (layer_3[63] & layer_3[63]); 
    assign layer_4[77] = ~(layer_3[83] ^ layer_3[89]); 
    assign layer_4[78] = ~layer_3[63]; 
    assign layer_4[79] = layer_3[78] ^ layer_3[81]; 
    assign layer_4[80] = layer_3[65] & ~layer_3[94]; 
    assign layer_4[81] = layer_3[85] & ~layer_3[88]; 
    assign layer_4[82] = ~(layer_3[93] | layer_3[82]); 
    assign layer_4[83] = ~layer_3[73] | (layer_3[73] & layer_3[85]); 
    assign layer_4[84] = layer_3[85]; 
    assign layer_4[85] = 1'b1; 
    assign layer_4[86] = ~layer_3[78]; 
    assign layer_4[87] = ~layer_3[100] | (layer_3[87] & layer_3[100]); 
    assign layer_4[88] = layer_3[81] & layer_3[71]; 
    assign layer_4[89] = ~(layer_3[85] & layer_3[84]); 
    assign layer_4[90] = ~(layer_3[97] ^ layer_3[83]); 
    assign layer_4[91] = 1'b1; 
    assign layer_4[92] = layer_3[82] & layer_3[84]; 
    assign layer_4[93] = layer_3[105]; 
    assign layer_4[94] = ~layer_3[109]; 
    assign layer_4[95] = ~layer_3[88] | (layer_3[88] & layer_3[96]); 
    assign layer_4[96] = 1'b0; 
    assign layer_4[97] = ~(layer_3[83] | layer_3[83]); 
    assign layer_4[98] = ~layer_3[91]; 
    assign layer_4[99] = layer_3[92] & ~layer_3[106]; 
    assign layer_4[100] = 1'b0; 
    assign layer_4[101] = ~(layer_3[103] & layer_3[85]); 
    assign layer_4[102] = layer_3[101] & layer_3[86]; 
    assign layer_4[103] = ~layer_3[101] | (layer_3[113] & layer_3[101]); 
    assign layer_4[104] = ~layer_3[117] | (layer_3[117] & layer_3[117]); 
    assign layer_4[105] = ~layer_3[95]; 
    assign layer_4[106] = 1'b0; 
    assign layer_4[107] = ~(layer_3[105] ^ layer_3[119]); 
    assign layer_4[108] = 1'b0; 
    assign layer_4[109] = layer_3[96] & ~layer_3[124]; 
    assign layer_4[110] = layer_3[99] & layer_3[115]; 
    assign layer_4[111] = layer_3[124]; 
    assign layer_4[112] = layer_3[116] & layer_3[103]; 
    assign layer_4[113] = layer_3[107] ^ layer_3[106]; 
    assign layer_4[114] = ~layer_3[103]; 
    assign layer_4[115] = layer_3[117] ^ layer_3[112]; 
    assign layer_4[116] = ~(layer_3[115] & layer_3[111]); 
    assign layer_4[117] = ~(layer_3[117] & layer_3[114]); 
    assign layer_4[118] = 1'b1; 
    assign layer_4[119] = ~layer_3[134]; 
    assign layer_4[120] = layer_3[135]; 
    assign layer_4[121] = layer_3[136]; 
    assign layer_4[122] = layer_3[135] & ~layer_3[129]; 
    assign layer_4[123] = ~layer_3[132] | (layer_3[134] & layer_3[132]); 
    assign layer_4[124] = layer_3[118]; 
    assign layer_4[125] = ~layer_3[127]; 
    assign layer_4[126] = ~layer_3[120] | (layer_3[120] & layer_3[116]); 
    assign layer_4[127] = ~(layer_3[132] ^ layer_3[124]); 
    assign layer_4[128] = layer_3[135] & layer_3[134]; 
    assign layer_4[129] = ~(layer_3[143] ^ layer_3[113]); 
    assign layer_4[130] = ~(layer_3[115] & layer_3[131]); 
    assign layer_4[131] = ~(layer_3[121] & layer_3[134]); 
    assign layer_4[132] = layer_3[117]; 
    assign layer_4[133] = layer_3[142] | layer_3[122]; 
    assign layer_4[134] = layer_3[149] & ~layer_3[132]; 
    assign layer_4[135] = ~(layer_3[119] | layer_3[141]); 
    assign layer_4[136] = ~(layer_3[149] | layer_3[120]); 
    assign layer_4[137] = ~(layer_3[131] | layer_3[122]); 
    assign layer_4[138] = ~layer_3[148] | (layer_3[132] & layer_3[148]); 
    assign layer_4[139] = 1'b1; 
    assign layer_4[140] = layer_3[137] & ~layer_3[129]; 
    assign layer_4[141] = 1'b0; 
    assign layer_4[142] = ~layer_3[141]; 
    assign layer_4[143] = 1'b1; 
    assign layer_4[144] = 1'b0; 
    assign layer_4[145] = 1'b0; 
    assign layer_4[146] = ~(layer_3[161] ^ layer_3[145]); 
    assign layer_4[147] = ~layer_3[151] | (layer_3[136] & layer_3[151]); 
    assign layer_4[148] = ~layer_3[158]; 
    assign layer_4[149] = layer_3[137] & ~layer_3[140]; 
    assign layer_4[150] = ~layer_3[157] | (layer_3[159] & layer_3[157]); 
    assign layer_4[151] = ~layer_3[143] | (layer_3[143] & layer_3[137]); 
    assign layer_4[152] = layer_3[142]; 
    assign layer_4[153] = ~(layer_3[167] ^ layer_3[142]); 
    assign layer_4[154] = ~(layer_3[162] | layer_3[140]); 
    assign layer_4[155] = layer_3[140] & layer_3[169]; 
    assign layer_4[156] = ~layer_3[139]; 
    assign layer_4[157] = layer_3[167] | layer_3[167]; 
    assign layer_4[158] = layer_3[143] | layer_3[159]; 
    assign layer_4[159] = ~layer_3[160] | (layer_3[165] & layer_3[160]); 
    assign layer_4[160] = layer_3[155] & ~layer_3[150]; 
    assign layer_4[161] = layer_3[162] ^ layer_3[168]; 
    assign layer_4[162] = ~layer_3[148] | (layer_3[153] & layer_3[148]); 
    assign layer_4[163] = layer_3[155]; 
    assign layer_4[164] = 1'b1; 
    assign layer_4[165] = ~layer_3[158]; 
    assign layer_4[166] = layer_3[169] | layer_3[155]; 
    assign layer_4[167] = layer_3[153] ^ layer_3[162]; 
    assign layer_4[168] = layer_3[155] & ~layer_3[171]; 
    assign layer_4[169] = layer_3[158]; 
    assign layer_4[170] = ~(layer_3[157] ^ layer_3[158]); 
    assign layer_4[171] = layer_3[161] ^ layer_3[185]; 
    assign layer_4[172] = 1'b0; 
    assign layer_4[173] = ~layer_3[161]; 
    assign layer_4[174] = ~layer_3[163] | (layer_3[163] & layer_3[172]); 
    assign layer_4[175] = 1'b1; 
    assign layer_4[176] = ~(layer_3[190] ^ layer_3[182]); 
    assign layer_4[177] = layer_3[189]; 
    assign layer_4[178] = ~(layer_3[180] | layer_3[172]); 
    assign layer_4[179] = layer_3[188] & ~layer_3[173]; 
    assign layer_4[180] = ~(layer_3[192] | layer_3[170]); 
    assign layer_4[181] = 1'b1; 
    assign layer_4[182] = layer_3[178] & ~layer_3[192]; 
    assign layer_4[183] = 1'b1; 
    assign layer_4[184] = layer_3[181]; 
    assign layer_4[185] = ~layer_3[192]; 
    assign layer_4[186] = layer_3[196] ^ layer_3[179]; 
    assign layer_4[187] = ~layer_3[202] | (layer_3[202] & layer_3[196]); 
    assign layer_4[188] = ~(layer_3[182] | layer_3[187]); 
    assign layer_4[189] = ~layer_3[177] | (layer_3[177] & layer_3[200]); 
    assign layer_4[190] = layer_3[191] & ~layer_3[201]; 
    assign layer_4[191] = layer_3[185] & layer_3[182]; 
    assign layer_4[192] = ~(layer_3[196] | layer_3[206]); 
    assign layer_4[193] = layer_3[182] & ~layer_3[185]; 
    assign layer_4[194] = ~layer_3[193] | (layer_3[193] & layer_3[209]); 
    assign layer_4[195] = ~layer_3[190] | (layer_3[204] & layer_3[190]); 
    assign layer_4[196] = ~(layer_3[182] & layer_3[180]); 
    assign layer_4[197] = ~(layer_3[201] ^ layer_3[196]); 
    assign layer_4[198] = ~layer_3[195] | (layer_3[214] & layer_3[195]); 
    assign layer_4[199] = layer_3[203] & ~layer_3[214]; 
    assign layer_4[200] = layer_3[186]; 
    assign layer_4[201] = ~(layer_3[206] ^ layer_3[204]); 
    assign layer_4[202] = layer_3[193] ^ layer_3[202]; 
    assign layer_4[203] = ~(layer_3[194] & layer_3[211]); 
    assign layer_4[204] = layer_3[206]; 
    assign layer_4[205] = ~(layer_3[216] & layer_3[217]); 
    assign layer_4[206] = ~layer_3[193]; 
    assign layer_4[207] = ~layer_3[194] | (layer_3[222] & layer_3[194]); 
    assign layer_4[208] = layer_3[224] & layer_3[214]; 
    assign layer_4[209] = ~layer_3[193] | (layer_3[193] & layer_3[210]); 
    assign layer_4[210] = 1'b0; 
    assign layer_4[211] = layer_3[207] ^ layer_3[221]; 
    assign layer_4[212] = ~(layer_3[205] & layer_3[196]); 
    assign layer_4[213] = layer_3[199] & layer_3[222]; 
    assign layer_4[214] = ~(layer_3[211] ^ layer_3[197]); 
    assign layer_4[215] = layer_3[221]; 
    assign layer_4[216] = 1'b0; 
    assign layer_4[217] = ~(layer_3[213] ^ layer_3[217]); 
    assign layer_4[218] = ~layer_3[227]; 
    assign layer_4[219] = layer_3[220] & layer_3[213]; 
    assign layer_4[220] = ~(layer_3[210] | layer_3[208]); 
    assign layer_4[221] = ~layer_3[237]; 
    assign layer_4[222] = layer_3[215] | layer_3[222]; 
    assign layer_4[223] = layer_3[218] & layer_3[237]; 
    assign layer_4[224] = ~layer_3[240] | (layer_3[240] & layer_3[236]); 
    assign layer_4[225] = ~(layer_3[215] & layer_3[227]); 
    assign layer_4[226] = layer_3[226]; 
    assign layer_4[227] = layer_3[237]; 
    assign layer_4[228] = ~layer_3[240]; 
    assign layer_4[229] = layer_3[213]; 
    assign layer_4[230] = ~(layer_3[246] & layer_3[244]); 
    assign layer_4[231] = layer_3[221] | layer_3[234]; 
    assign layer_4[232] = ~(layer_3[235] & layer_3[226]); 
    assign layer_4[233] = ~layer_3[234]; 
    assign layer_4[234] = layer_3[246] & ~layer_3[223]; 
    assign layer_4[235] = ~layer_3[225]; 
    assign layer_4[236] = ~layer_3[232] | (layer_3[232] & layer_3[251]); 
    assign layer_4[237] = ~layer_3[227]; 
    assign layer_4[238] = ~layer_3[235]; 
    assign layer_4[239] = ~(layer_3[247] | layer_3[224]); 
    assign layer_4[240] = layer_3[240] | layer_3[247]; 
    assign layer_4[241] = ~layer_3[244]; 
    assign layer_4[242] = layer_3[229]; 
    assign layer_4[243] = layer_3[237] ^ layer_3[246]; 
    assign layer_4[244] = layer_3[236] | layer_3[228]; 
    assign layer_4[245] = 1'b0; 
    assign layer_4[246] = ~(layer_3[247] & layer_3[248]); 
    assign layer_4[247] = layer_3[259]; 
    assign layer_4[248] = ~layer_3[259] | (layer_3[259] & layer_3[231]); 
    assign layer_4[249] = layer_3[242] & layer_3[262]; 
    assign layer_4[250] = ~layer_3[241]; 
    assign layer_4[251] = ~(layer_3[251] ^ layer_3[237]); 
    assign layer_4[252] = layer_3[254] | layer_3[237]; 
    assign layer_4[253] = layer_3[266] | layer_3[241]; 
    assign layer_4[254] = ~(layer_3[254] & layer_3[266]); 
    assign layer_4[255] = layer_3[240]; 
    assign layer_4[256] = ~layer_3[241]; 
    assign layer_4[257] = ~layer_3[251] | (layer_3[251] & layer_3[267]); 
    assign layer_4[258] = layer_3[268] ^ layer_3[272]; 
    assign layer_4[259] = ~layer_3[266] | (layer_3[267] & layer_3[266]); 
    assign layer_4[260] = ~(layer_3[271] & layer_3[260]); 
    assign layer_4[261] = layer_3[253]; 
    assign layer_4[262] = ~(layer_3[278] | layer_3[264]); 
    assign layer_4[263] = layer_3[276] & ~layer_3[248]; 
    assign layer_4[264] = ~layer_3[274] | (layer_3[274] & layer_3[253]); 
    assign layer_4[265] = ~(layer_3[266] ^ layer_3[279]); 
    assign layer_4[266] = ~layer_3[267]; 
    assign layer_4[267] = layer_3[257] | layer_3[255]; 
    assign layer_4[268] = 1'b0; 
    assign layer_4[269] = layer_3[263] & layer_3[253]; 
    assign layer_4[270] = ~(layer_3[278] ^ layer_3[260]); 
    assign layer_4[271] = layer_3[278]; 
    assign layer_4[272] = ~layer_3[285]; 
    assign layer_4[273] = ~layer_3[287]; 
    assign layer_4[274] = layer_3[285]; 
    assign layer_4[275] = ~layer_3[282]; 
    assign layer_4[276] = ~layer_3[281]; 
    assign layer_4[277] = 1'b1; 
    assign layer_4[278] = ~layer_3[278] | (layer_3[288] & layer_3[278]); 
    assign layer_4[279] = layer_3[280] & layer_3[286]; 
    assign layer_4[280] = layer_3[292] & ~layer_3[284]; 
    assign layer_4[281] = layer_3[294] & ~layer_3[290]; 
    assign layer_4[282] = layer_3[288] & ~layer_3[279]; 
    assign layer_4[283] = layer_3[292] & ~layer_3[289]; 
    assign layer_4[284] = layer_3[295] | layer_3[277]; 
    assign layer_4[285] = 1'b1; 
    assign layer_4[286] = layer_3[299] & layer_3[276]; 
    assign layer_4[287] = layer_3[301] & ~layer_3[277]; 
    assign layer_4[288] = ~layer_3[296]; 
    assign layer_4[289] = ~layer_3[278]; 
    assign layer_4[290] = ~layer_3[279]; 
    assign layer_4[291] = ~(layer_3[287] & layer_3[282]); 
    assign layer_4[292] = layer_3[293] | layer_3[287]; 
    assign layer_4[293] = ~(layer_3[308] & layer_3[300]); 
    assign layer_4[294] = ~layer_3[299] | (layer_3[299] & layer_3[297]); 
    assign layer_4[295] = layer_3[310] & layer_3[288]; 
    assign layer_4[296] = layer_3[312]; 
    assign layer_4[297] = layer_3[283] ^ layer_3[289]; 
    assign layer_4[298] = layer_3[303] & ~layer_3[307]; 
    assign layer_4[299] = ~layer_3[314]; 
    assign layer_4[300] = ~layer_3[295]; 
    assign layer_4[301] = layer_3[285] | layer_3[294]; 
    assign layer_4[302] = 1'b0; 
    assign layer_4[303] = layer_3[291] | layer_3[296]; 
    assign layer_4[304] = ~layer_3[310]; 
    assign layer_4[305] = layer_3[293]; 
    assign layer_4[306] = ~layer_3[320]; 
    assign layer_4[307] = ~(layer_3[314] | layer_3[308]); 
    assign layer_4[308] = layer_3[312] & layer_3[316]; 
    assign layer_4[309] = ~(layer_3[322] ^ layer_3[304]); 
    assign layer_4[310] = layer_3[316] & ~layer_3[321]; 
    assign layer_4[311] = ~layer_3[300] | (layer_3[311] & layer_3[300]); 
    assign layer_4[312] = ~(layer_3[309] & layer_3[302]); 
    assign layer_4[313] = ~layer_3[323] | (layer_3[323] & layer_3[303]); 
    assign layer_4[314] = ~layer_3[317] | (layer_3[300] & layer_3[317]); 
    assign layer_4[315] = layer_3[307] ^ layer_3[302]; 
    assign layer_4[316] = layer_3[301] | layer_3[322]; 
    assign layer_4[317] = ~(layer_3[327] & layer_3[315]); 
    assign layer_4[318] = ~(layer_3[307] ^ layer_3[307]); 
    assign layer_4[319] = layer_3[328] ^ layer_3[334]; 
    assign layer_4[320] = ~layer_3[308]; 
    assign layer_4[321] = ~layer_3[326] | (layer_3[326] & layer_3[313]); 
    assign layer_4[322] = 1'b0; 
    assign layer_4[323] = ~layer_3[313]; 
    assign layer_4[324] = layer_3[330] | layer_3[317]; 
    assign layer_4[325] = ~layer_3[316] | (layer_3[320] & layer_3[316]); 
    assign layer_4[326] = ~(layer_3[329] ^ layer_3[338]); 
    assign layer_4[327] = layer_3[332] & ~layer_3[331]; 
    assign layer_4[328] = layer_3[320] | layer_3[315]; 
    assign layer_4[329] = layer_3[318]; 
    assign layer_4[330] = layer_3[328] & ~layer_3[326]; 
    assign layer_4[331] = ~layer_3[331] | (layer_3[331] & layer_3[344]); 
    assign layer_4[332] = layer_3[340]; 
    assign layer_4[333] = ~layer_3[321]; 
    assign layer_4[334] = ~(layer_3[323] ^ layer_3[342]); 
    assign layer_4[335] = layer_3[322] | layer_3[322]; 
    assign layer_4[336] = 1'b0; 
    assign layer_4[337] = ~(layer_3[348] & layer_3[346]); 
    assign layer_4[338] = ~(layer_3[350] & layer_3[334]); 
    assign layer_4[339] = 1'b0; 
    assign layer_4[340] = layer_3[329] | layer_3[326]; 
    assign layer_4[341] = ~layer_3[353]; 
    assign layer_4[342] = layer_3[333] ^ layer_3[332]; 
    assign layer_4[343] = ~(layer_3[333] | layer_3[357]); 
    assign layer_4[344] = ~(layer_3[336] ^ layer_3[348]); 
    assign layer_4[345] = 1'b1; 
    assign layer_4[346] = ~layer_3[350]; 
    assign layer_4[347] = layer_3[346] & ~layer_3[335]; 
    assign layer_4[348] = layer_3[338] | layer_3[334]; 
    assign layer_4[349] = 1'b0; 
    assign layer_4[350] = ~layer_3[353] | (layer_3[353] & layer_3[338]); 
    assign layer_4[351] = ~(layer_3[335] & layer_3[366]); 
    assign layer_4[352] = ~(layer_3[353] ^ layer_3[353]); 
    assign layer_4[353] = ~(layer_3[365] & layer_3[368]); 
    assign layer_4[354] = ~layer_3[344]; 
    assign layer_4[355] = ~(layer_3[358] | layer_3[356]); 
    assign layer_4[356] = ~(layer_3[355] | layer_3[360]); 
    assign layer_4[357] = layer_3[372] & ~layer_3[343]; 
    assign layer_4[358] = ~layer_3[358] | (layer_3[358] & layer_3[343]); 
    assign layer_4[359] = ~(layer_3[360] | layer_3[357]); 
    assign layer_4[360] = layer_3[371] & layer_3[367]; 
    assign layer_4[361] = layer_3[375]; 
    assign layer_4[362] = layer_3[351] | layer_3[348]; 
    assign layer_4[363] = layer_3[375] & layer_3[354]; 
    assign layer_4[364] = ~layer_3[371] | (layer_3[379] & layer_3[371]); 
    assign layer_4[365] = ~(layer_3[364] | layer_3[354]); 
    assign layer_4[366] = ~layer_3[381]; 
    assign layer_4[367] = ~layer_3[360]; 
    assign layer_4[368] = ~(layer_3[359] ^ layer_3[358]); 
    assign layer_4[369] = layer_3[366]; 
    assign layer_4[370] = layer_3[363] ^ layer_3[360]; 
    assign layer_4[371] = ~layer_3[364] | (layer_3[364] & layer_3[369]); 
    assign layer_4[372] = ~layer_3[364]; 
    assign layer_4[373] = layer_3[365] & layer_3[364]; 
    assign layer_4[374] = ~layer_3[380] | (layer_3[380] & layer_3[385]); 
    assign layer_4[375] = ~(layer_3[385] ^ layer_3[358]); 
    assign layer_4[376] = layer_3[372] & ~layer_3[367]; 
    assign layer_4[377] = layer_3[375] | layer_3[362]; 
    assign layer_4[378] = layer_3[371] ^ layer_3[381]; 
    assign layer_4[379] = ~layer_3[381]; 
    assign layer_4[380] = ~layer_3[366]; 
    assign layer_4[381] = ~(layer_3[373] | layer_3[380]); 
    assign layer_4[382] = ~layer_3[370]; 
    assign layer_4[383] = layer_3[373]; 
    assign layer_4[384] = ~layer_3[387] | (layer_3[387] & layer_3[394]); 
    assign layer_4[385] = layer_3[377] & ~layer_3[370]; 
    assign layer_4[386] = ~layer_3[387]; 
    assign layer_4[387] = ~layer_3[378] | (layer_3[398] & layer_3[378]); 
    assign layer_4[388] = ~(layer_3[392] | layer_3[396]); 
    assign layer_4[389] = ~layer_3[393] | (layer_3[403] & layer_3[393]); 
    assign layer_4[390] = 1'b0; 
    assign layer_4[391] = ~(layer_3[404] ^ layer_3[384]); 
    assign layer_4[392] = ~layer_3[404] | (layer_3[404] & layer_3[375]); 
    assign layer_4[393] = layer_3[381] & ~layer_3[390]; 
    assign layer_4[394] = layer_3[379] & ~layer_3[392]; 
    assign layer_4[395] = ~layer_3[386] | (layer_3[386] & layer_3[384]); 
    assign layer_4[396] = ~(layer_3[398] & layer_3[382]); 
    assign layer_4[397] = 1'b0; 
    assign layer_4[398] = layer_3[411] & ~layer_3[399]; 
    assign layer_4[399] = ~(layer_3[409] ^ layer_3[401]); 
    assign layer_4[400] = layer_3[389] & layer_3[384]; 
    assign layer_4[401] = layer_3[386] & layer_3[395]; 
    assign layer_4[402] = layer_3[398] & layer_3[388]; 
    assign layer_4[403] = layer_3[388] & ~layer_3[396]; 
    assign layer_4[404] = ~(layer_3[396] | layer_3[390]); 
    assign layer_4[405] = layer_3[394] | layer_3[415]; 
    assign layer_4[406] = layer_3[408] & ~layer_3[399]; 
    assign layer_4[407] = ~(layer_3[402] | layer_3[408]); 
    assign layer_4[408] = ~(layer_3[399] | layer_3[410]); 
    assign layer_4[409] = ~layer_3[419]; 
    assign layer_4[410] = layer_3[411]; 
    assign layer_4[411] = 1'b0; 
    assign layer_4[412] = 1'b0; 
    assign layer_4[413] = layer_3[424] & ~layer_3[411]; 
    assign layer_4[414] = ~(layer_3[408] & layer_3[417]); 
    assign layer_4[415] = ~layer_3[409]; 
    assign layer_4[416] = ~layer_3[409] | (layer_3[409] & layer_3[405]); 
    assign layer_4[417] = layer_3[429]; 
    assign layer_4[418] = 1'b1; 
    assign layer_4[419] = layer_3[418] | layer_3[424]; 
    assign layer_4[420] = 1'b1; 
    assign layer_4[421] = 1'b0; 
    assign layer_4[422] = layer_3[418]; 
    assign layer_4[423] = layer_3[437] & ~layer_3[419]; 
    assign layer_4[424] = layer_3[419] & ~layer_3[408]; 
    assign layer_4[425] = ~(layer_3[439] ^ layer_3[409]); 
    assign layer_4[426] = layer_3[435] & ~layer_3[414]; 
    assign layer_4[427] = 1'b0; 
    assign layer_4[428] = ~layer_3[413] | (layer_3[413] & layer_3[417]); 
    assign layer_4[429] = layer_3[444] ^ layer_3[434]; 
    assign layer_4[430] = ~(layer_3[415] | layer_3[427]); 
    assign layer_4[431] = 1'b0; 
    assign layer_4[432] = ~layer_3[447] | (layer_3[438] & layer_3[447]); 
    assign layer_4[433] = layer_3[426] & layer_3[439]; 
    assign layer_4[434] = layer_3[435] & ~layer_3[426]; 
    assign layer_4[435] = 1'b1; 
    assign layer_4[436] = layer_3[431]; 
    assign layer_4[437] = 1'b1; 
    assign layer_4[438] = ~layer_3[445] | (layer_3[450] & layer_3[445]); 
    assign layer_4[439] = 1'b0; 
    assign layer_4[440] = ~layer_3[445]; 
    assign layer_4[441] = ~(layer_3[431] | layer_3[456]); 
    assign layer_4[442] = layer_3[430] & layer_3[441]; 
    assign layer_4[443] = layer_3[438] | layer_3[441]; 
    assign layer_4[444] = ~layer_3[431] | (layer_3[431] & layer_3[430]); 
    assign layer_4[445] = ~layer_3[437] | (layer_3[454] & layer_3[437]); 
    assign layer_4[446] = ~layer_3[444] | (layer_3[444] & layer_3[450]); 
    assign layer_4[447] = layer_3[453]; 
    assign layer_4[448] = layer_3[458] & ~layer_3[447]; 
    assign layer_4[449] = layer_3[462]; 
    assign layer_4[450] = layer_3[436]; 
    assign layer_4[451] = 1'b1; 
    assign layer_4[452] = layer_3[436] & layer_3[463]; 
    assign layer_4[453] = ~layer_3[459] | (layer_3[459] & layer_3[455]); 
    assign layer_4[454] = layer_3[462]; 
    assign layer_4[455] = ~(layer_3[452] & layer_3[461]); 
    assign layer_4[456] = layer_3[444]; 
    assign layer_4[457] = layer_3[450] & layer_3[448]; 
    assign layer_4[458] = ~layer_3[460] | (layer_3[460] & layer_3[465]); 
    assign layer_4[459] = layer_3[455] ^ layer_3[474]; 
    assign layer_4[460] = layer_3[466] | layer_3[455]; 
    assign layer_4[461] = layer_3[464] & ~layer_3[455]; 
    assign layer_4[462] = ~layer_3[454]; 
    assign layer_4[463] = layer_3[470] | layer_3[458]; 
    assign layer_4[464] = layer_3[471] & layer_3[463]; 
    assign layer_4[465] = layer_3[462] & ~layer_3[472]; 
    assign layer_4[466] = layer_3[451]; 
    assign layer_4[467] = ~layer_3[451] | (layer_3[451] & layer_3[461]); 
    assign layer_4[468] = layer_3[466] | layer_3[476]; 
    assign layer_4[469] = ~(layer_3[471] | layer_3[458]); 
    assign layer_4[470] = layer_3[484]; 
    assign layer_4[471] = layer_3[467]; 
    assign layer_4[472] = layer_3[484] & ~layer_3[461]; 
    assign layer_4[473] = ~(layer_3[476] ^ layer_3[458]); 
    assign layer_4[474] = layer_3[478] & layer_3[468]; 
    assign layer_4[475] = layer_3[473] ^ layer_3[485]; 
    assign layer_4[476] = layer_3[472] | layer_3[480]; 
    assign layer_4[477] = 1'b0; 
    assign layer_4[478] = ~(layer_3[480] & layer_3[469]); 
    assign layer_4[479] = layer_3[485]; 
    assign layer_4[480] = ~layer_3[467]; 
    assign layer_4[481] = ~layer_3[492]; 
    assign layer_4[482] = ~layer_3[465]; 
    assign layer_4[483] = ~layer_3[471]; 
    assign layer_4[484] = layer_3[483] ^ layer_3[486]; 
    assign layer_4[485] = layer_3[501] | layer_3[483]; 
    assign layer_4[486] = layer_3[492] | layer_3[501]; 
    assign layer_4[487] = 1'b1; 
    assign layer_4[488] = ~(layer_3[485] & layer_3[489]); 
    assign layer_4[489] = layer_3[498] & ~layer_3[490]; 
    assign layer_4[490] = ~layer_3[475] | (layer_3[476] & layer_3[475]); 
    assign layer_4[491] = layer_3[493]; 
    assign layer_4[492] = layer_3[476] & layer_3[477]; 
    assign layer_4[493] = 1'b1; 
    assign layer_4[494] = layer_3[487] & ~layer_3[494]; 
    assign layer_4[495] = layer_3[494]; 
    assign layer_4[496] = layer_3[511] | layer_3[508]; 
    assign layer_4[497] = 1'b0; 
    assign layer_4[498] = ~layer_3[494]; 
    assign layer_4[499] = layer_3[486]; 
    assign layer_4[500] = ~layer_3[500] | (layer_3[484] & layer_3[500]); 
    assign layer_4[501] = ~(layer_3[490] & layer_3[485]); 
    assign layer_4[502] = layer_3[495]; 
    assign layer_4[503] = layer_3[515] & ~layer_3[514]; 
    assign layer_4[504] = layer_3[488] & ~layer_3[491]; 
    assign layer_4[505] = layer_3[509] & ~layer_3[519]; 
    assign layer_4[506] = layer_3[516] & ~layer_3[507]; 
    assign layer_4[507] = layer_3[513]; 
    assign layer_4[508] = ~(layer_3[524] & layer_3[513]); 
    assign layer_4[509] = layer_3[506] ^ layer_3[515]; 
    assign layer_4[510] = 1'b1; 
    assign layer_4[511] = layer_3[513] ^ layer_3[514]; 
    assign layer_4[512] = layer_3[511] & layer_3[511]; 
    assign layer_4[513] = ~layer_3[526] | (layer_3[511] & layer_3[526]); 
    assign layer_4[514] = ~(layer_3[501] | layer_3[506]); 
    assign layer_4[515] = layer_3[510]; 
    assign layer_4[516] = layer_3[510]; 
    assign layer_4[517] = layer_3[520] | layer_3[500]; 
    assign layer_4[518] = ~layer_3[529] | (layer_3[529] & layer_3[532]); 
    assign layer_4[519] = ~layer_3[525] | (layer_3[525] & layer_3[503]); 
    assign layer_4[520] = ~(layer_3[517] ^ layer_3[504]); 
    assign layer_4[521] = layer_3[514] ^ layer_3[529]; 
    assign layer_4[522] = layer_3[512] ^ layer_3[513]; 
    assign layer_4[523] = ~layer_3[538] | (layer_3[515] & layer_3[538]); 
    assign layer_4[524] = 1'b0; 
    assign layer_4[525] = 1'b0; 
    assign layer_4[526] = 1'b1; 
    assign layer_4[527] = layer_3[526] & layer_3[528]; 
    assign layer_4[528] = ~(layer_3[523] | layer_3[539]); 
    assign layer_4[529] = ~layer_3[523] | (layer_3[534] & layer_3[523]); 
    assign layer_4[530] = ~layer_3[527]; 
    assign layer_4[531] = layer_3[532]; 
    assign layer_4[532] = ~layer_3[527] | (layer_3[527] & layer_3[526]); 
    assign layer_4[533] = ~(layer_3[519] ^ layer_3[542]); 
    assign layer_4[534] = ~layer_3[540] | (layer_3[520] & layer_3[540]); 
    assign layer_4[535] = 1'b0; 
    assign layer_4[536] = layer_3[542]; 
    assign layer_4[537] = layer_3[541]; 
    assign layer_4[538] = layer_3[550] & ~layer_3[531]; 
    assign layer_4[539] = ~(layer_3[531] | layer_3[522]); 
    assign layer_4[540] = layer_3[551]; 
    assign layer_4[541] = layer_3[548] ^ layer_3[526]; 
    assign layer_4[542] = 1'b0; 
    assign layer_4[543] = layer_3[535] ^ layer_3[531]; 
    assign layer_4[544] = ~(layer_3[534] & layer_3[540]); 
    assign layer_4[545] = ~layer_3[536] | (layer_3[536] & layer_3[533]); 
    assign layer_4[546] = layer_3[535] & ~layer_3[546]; 
    assign layer_4[547] = layer_3[553]; 
    assign layer_4[548] = ~layer_3[536] | (layer_3[555] & layer_3[536]); 
    assign layer_4[549] = layer_3[534] ^ layer_3[554]; 
    assign layer_4[550] = ~layer_3[542] | (layer_3[542] & layer_3[543]); 
    assign layer_4[551] = layer_3[543] & layer_3[553]; 
    assign layer_4[552] = layer_3[553] & ~layer_3[556]; 
    assign layer_4[553] = ~(layer_3[541] & layer_3[556]); 
    assign layer_4[554] = layer_3[543] ^ layer_3[550]; 
    assign layer_4[555] = layer_3[544] & layer_3[542]; 
    assign layer_4[556] = layer_3[547] | layer_3[558]; 
    assign layer_4[557] = ~(layer_3[556] & layer_3[555]); 
    assign layer_4[558] = layer_3[573]; 
    assign layer_4[559] = ~(layer_3[565] | layer_3[545]); 
    assign layer_4[560] = ~layer_3[557] | (layer_3[551] & layer_3[557]); 
    assign layer_4[561] = ~layer_3[573] | (layer_3[573] & layer_3[573]); 
    assign layer_4[562] = ~(layer_3[570] ^ layer_3[566]); 
    assign layer_4[563] = layer_3[554] & layer_3[548]; 
    assign layer_4[564] = layer_3[577] & layer_3[557]; 
    assign layer_4[565] = ~(layer_3[566] ^ layer_3[552]); 
    assign layer_4[566] = ~layer_3[572] | (layer_3[572] & layer_3[557]); 
    assign layer_4[567] = ~layer_3[569]; 
    assign layer_4[568] = ~layer_3[578] | (layer_3[578] & layer_3[555]); 
    assign layer_4[569] = ~layer_3[566]; 
    assign layer_4[570] = ~layer_3[573] | (layer_3[578] & layer_3[573]); 
    assign layer_4[571] = layer_3[558] | layer_3[557]; 
    assign layer_4[572] = ~layer_3[558] | (layer_3[568] & layer_3[558]); 
    assign layer_4[573] = ~(layer_3[580] | layer_3[586]); 
    assign layer_4[574] = layer_3[567] | layer_3[582]; 
    assign layer_4[575] = layer_3[563]; 
    assign layer_4[576] = layer_3[561]; 
    assign layer_4[577] = ~(layer_3[573] ^ layer_3[563]); 
    assign layer_4[578] = ~layer_3[577]; 
    assign layer_4[579] = layer_3[565] ^ layer_3[586]; 
    assign layer_4[580] = 1'b1; 
    assign layer_4[581] = ~layer_3[580] | (layer_3[585] & layer_3[580]); 
    assign layer_4[582] = layer_3[592]; 
    assign layer_4[583] = 1'b1; 
    assign layer_4[584] = layer_3[569] & ~layer_3[572]; 
    assign layer_4[585] = 1'b0; 
    assign layer_4[586] = ~layer_3[582] | (layer_3[582] & layer_3[593]); 
    assign layer_4[587] = ~(layer_3[596] | layer_3[594]); 
    assign layer_4[588] = 1'b0; 
    assign layer_4[589] = ~layer_3[575]; 
    assign layer_4[590] = layer_3[598] & ~layer_3[578]; 
    assign layer_4[591] = ~layer_3[577]; 
    assign layer_4[592] = layer_3[600] & ~layer_3[583]; 
    assign layer_4[593] = layer_3[595] & layer_3[604]; 
    assign layer_4[594] = ~(layer_3[602] ^ layer_3[593]); 
    assign layer_4[595] = layer_3[605] | layer_3[597]; 
    assign layer_4[596] = layer_3[602] ^ layer_3[605]; 
    assign layer_4[597] = ~(layer_3[589] ^ layer_3[610]); 
    assign layer_4[598] = ~layer_3[602] | (layer_3[598] & layer_3[602]); 
    assign layer_4[599] = layer_3[610]; 
    assign layer_4[600] = layer_3[588] | layer_3[593]; 
    assign layer_4[601] = layer_3[596] & ~layer_3[601]; 
    assign layer_4[602] = 1'b0; 
    assign layer_4[603] = layer_3[618] & ~layer_3[607]; 
    assign layer_4[604] = ~(layer_3[609] ^ layer_3[617]); 
    assign layer_4[605] = ~(layer_3[607] ^ layer_3[614]); 
    assign layer_4[606] = layer_3[604] | layer_3[589]; 
    assign layer_4[607] = layer_3[612] & ~layer_3[602]; 
    assign layer_4[608] = 1'b1; 
    assign layer_4[609] = ~(layer_3[594] & layer_3[620]); 
    assign layer_4[610] = layer_3[596] | layer_3[614]; 
    assign layer_4[611] = ~(layer_3[597] & layer_3[616]); 
    assign layer_4[612] = 1'b1; 
    assign layer_4[613] = ~(layer_3[606] ^ layer_3[598]); 
    assign layer_4[614] = ~(layer_3[616] ^ layer_3[618]); 
    assign layer_4[615] = layer_3[628] & layer_3[606]; 
    assign layer_4[616] = layer_3[613] & ~layer_3[620]; 
    assign layer_4[617] = ~(layer_3[631] | layer_3[629]); 
    assign layer_4[618] = ~layer_3[611] | (layer_3[631] & layer_3[611]); 
    assign layer_4[619] = ~(layer_3[627] | layer_3[628]); 
    assign layer_4[620] = layer_3[627] ^ layer_3[622]; 
    assign layer_4[621] = ~(layer_3[619] ^ layer_3[624]); 
    assign layer_4[622] = layer_3[629] & ~layer_3[609]; 
    assign layer_4[623] = ~layer_3[616]; 
    assign layer_4[624] = ~layer_3[617]; 
    assign layer_4[625] = layer_3[612] & ~layer_3[611]; 
    assign layer_4[626] = layer_3[624] & ~layer_3[613]; 
    assign layer_4[627] = layer_3[612] | layer_3[636]; 
    assign layer_4[628] = 1'b1; 
    assign layer_4[629] = ~(layer_3[642] | layer_3[639]); 
    assign layer_4[630] = ~layer_3[613]; 
    assign layer_4[631] = layer_3[637] & ~layer_3[623]; 
    assign layer_4[632] = ~layer_3[633] | (layer_3[633] & layer_3[635]); 
    assign layer_4[633] = layer_3[627]; 
    assign layer_4[634] = ~layer_3[640] | (layer_3[618] & layer_3[640]); 
    assign layer_4[635] = layer_3[633] | layer_3[645]; 
    assign layer_4[636] = layer_3[640]; 
    assign layer_4[637] = ~(layer_3[640] & layer_3[638]); 
    assign layer_4[638] = layer_3[635] | layer_3[650]; 
    assign layer_4[639] = ~layer_3[642]; 
    assign layer_4[640] = ~(layer_3[651] | layer_3[646]); 
    assign layer_4[641] = layer_3[632] & ~layer_3[641]; 
    assign layer_4[642] = layer_3[650] & layer_3[636]; 
    assign layer_4[643] = layer_3[636]; 
    assign layer_4[644] = layer_3[639] & ~layer_3[658]; 
    assign layer_4[645] = ~layer_3[654] | (layer_3[658] & layer_3[654]); 
    assign layer_4[646] = 1'b0; 
    assign layer_4[647] = ~layer_3[635]; 
    assign layer_4[648] = ~(layer_3[637] ^ layer_3[642]); 
    assign layer_4[649] = ~layer_3[646]; 
    assign layer_4[650] = ~(layer_3[659] & layer_3[647]); 
    assign layer_4[651] = layer_3[639] ^ layer_3[644]; 
    assign layer_4[652] = 1'b1; 
    assign layer_4[653] = ~layer_3[668] | (layer_3[654] & layer_3[668]); 
    assign layer_4[654] = ~layer_3[657] | (layer_3[669] & layer_3[657]); 
    assign layer_4[655] = ~(layer_3[660] & layer_3[656]); 
    assign layer_4[656] = layer_3[655] & layer_3[660]; 
    assign layer_4[657] = layer_3[658] & ~layer_3[668]; 
    assign layer_4[658] = ~layer_3[645]; 
    assign layer_4[659] = ~(layer_3[672] & layer_3[644]); 
    assign layer_4[660] = layer_3[666]; 
    assign layer_4[661] = ~layer_3[655]; 
    assign layer_4[662] = ~(layer_3[659] | layer_3[665]); 
    assign layer_4[663] = layer_3[679] ^ layer_3[659]; 
    assign layer_4[664] = ~layer_3[655] | (layer_3[655] & layer_3[648]); 
    assign layer_4[665] = layer_3[649] & ~layer_3[659]; 
    assign layer_4[666] = 1'b1; 
    assign layer_4[667] = layer_3[658]; 
    assign layer_4[668] = layer_3[684] | layer_3[654]; 
    assign layer_4[669] = layer_3[657]; 
    assign layer_4[670] = ~(layer_3[678] & layer_3[670]); 
    assign layer_4[671] = layer_3[671] & ~layer_3[679]; 
    assign layer_4[672] = ~(layer_3[674] & layer_3[683]); 
    assign layer_4[673] = ~layer_3[673]; 
    assign layer_4[674] = ~(layer_3[661] ^ layer_3[684]); 
    assign layer_4[675] = ~(layer_3[659] ^ layer_3[680]); 
    assign layer_4[676] = ~layer_3[668] | (layer_3[668] & layer_3[680]); 
    assign layer_4[677] = ~(layer_3[668] & layer_3[675]); 
    assign layer_4[678] = ~(layer_3[672] & layer_3[681]); 
    assign layer_4[679] = ~layer_3[674]; 
    assign layer_4[680] = ~(layer_3[679] | layer_3[690]); 
    assign layer_4[681] = ~layer_3[668]; 
    assign layer_4[682] = layer_3[678]; 
    assign layer_4[683] = layer_3[667] & ~layer_3[694]; 
    assign layer_4[684] = ~layer_3[668]; 
    assign layer_4[685] = ~(layer_3[686] & layer_3[695]); 
    assign layer_4[686] = 1'b0; 
    assign layer_4[687] = ~layer_3[700] | (layer_3[700] & layer_3[699]); 
    assign layer_4[688] = layer_3[687]; 
    assign layer_4[689] = ~layer_3[685] | (layer_3[685] & layer_3[700]); 
    assign layer_4[690] = ~(layer_3[694] & layer_3[694]); 
    assign layer_4[691] = ~(layer_3[698] | layer_3[702]); 
    assign layer_4[692] = 1'b1; 
    assign layer_4[693] = ~(layer_3[692] | layer_3[677]); 
    assign layer_4[694] = ~(layer_3[699] ^ layer_3[699]); 
    assign layer_4[695] = layer_3[700] & ~layer_3[678]; 
    assign layer_4[696] = 1'b0; 
    assign layer_4[697] = layer_3[696]; 
    assign layer_4[698] = layer_3[696] ^ layer_3[683]; 
    assign layer_4[699] = layer_3[695]; 
    assign layer_4[700] = layer_3[693] | layer_3[694]; 
    assign layer_4[701] = layer_3[707] | layer_3[685]; 
    assign layer_4[702] = 1'b0; 
    assign layer_4[703] = layer_3[716] & ~layer_3[708]; 
    assign layer_4[704] = layer_3[718] & ~layer_3[705]; 
    assign layer_4[705] = layer_3[721] & ~layer_3[703]; 
    assign layer_4[706] = layer_3[719] & ~layer_3[696]; 
    assign layer_4[707] = layer_3[708] & ~layer_3[700]; 
    assign layer_4[708] = 1'b1; 
    assign layer_4[709] = layer_3[719]; 
    assign layer_4[710] = layer_3[706] | layer_3[716]; 
    assign layer_4[711] = layer_3[706] & layer_3[722]; 
    assign layer_4[712] = ~(layer_3[721] & layer_3[726]); 
    assign layer_4[713] = layer_3[712]; 
    assign layer_4[714] = layer_3[713] & ~layer_3[718]; 
    assign layer_4[715] = layer_3[731] & layer_3[701]; 
    assign layer_4[716] = ~(layer_3[724] & layer_3[729]); 
    assign layer_4[717] = layer_3[730] ^ layer_3[724]; 
    assign layer_4[718] = layer_3[703] ^ layer_3[724]; 
    assign layer_4[719] = ~layer_3[722] | (layer_3[722] & layer_3[728]); 
    assign layer_4[720] = ~layer_3[711] | (layer_3[711] & layer_3[724]); 
    assign layer_4[721] = layer_3[729] & ~layer_3[705]; 
    assign layer_4[722] = ~layer_3[721]; 
    assign layer_4[723] = 1'b0; 
    assign layer_4[724] = layer_3[730] & ~layer_3[734]; 
    assign layer_4[725] = layer_3[734] ^ layer_3[718]; 
    assign layer_4[726] = ~layer_3[710] | (layer_3[710] & layer_3[715]); 
    assign layer_4[727] = ~(layer_3[718] & layer_3[726]); 
    assign layer_4[728] = layer_3[737] & layer_3[722]; 
    assign layer_4[729] = ~(layer_3[718] ^ layer_3[742]); 
    assign layer_4[730] = ~(layer_3[728] | layer_3[733]); 
    assign layer_4[731] = ~(layer_3[715] ^ layer_3[746]); 
    assign layer_4[732] = layer_3[737] & layer_3[732]; 
    assign layer_4[733] = 1'b0; 
    assign layer_4[734] = layer_3[742] & ~layer_3[749]; 
    assign layer_4[735] = layer_3[719] & layer_3[718]; 
    assign layer_4[736] = layer_3[734]; 
    assign layer_4[737] = layer_3[735] | layer_3[738]; 
    assign layer_4[738] = layer_3[750]; 
    assign layer_4[739] = ~layer_3[749] | (layer_3[749] & layer_3[751]); 
    assign layer_4[740] = 1'b0; 
    assign layer_4[741] = 1'b0; 
    assign layer_4[742] = ~layer_3[735]; 
    assign layer_4[743] = 1'b1; 
    assign layer_4[744] = layer_3[757]; 
    assign layer_4[745] = ~layer_3[729] | (layer_3[746] & layer_3[729]); 
    assign layer_4[746] = ~(layer_3[744] & layer_3[755]); 
    assign layer_4[747] = ~(layer_3[741] | layer_3[753]); 
    assign layer_4[748] = ~layer_3[761] | (layer_3[761] & layer_3[755]); 
    assign layer_4[749] = ~(layer_3[762] | layer_3[739]); 
    assign layer_4[750] = layer_3[762] & layer_3[761]; 
    assign layer_4[751] = layer_3[735] ^ layer_3[745]; 
    assign layer_4[752] = layer_3[760] & ~layer_3[748]; 
    assign layer_4[753] = ~(layer_3[758] ^ layer_3[736]); 
    assign layer_4[754] = ~layer_3[747] | (layer_3[747] & layer_3[743]); 
    assign layer_4[755] = layer_3[765] & ~layer_3[744]; 
    assign layer_4[756] = 1'b1; 
    assign layer_4[757] = layer_3[764] & layer_3[751]; 
    assign layer_4[758] = 1'b1; 
    assign layer_4[759] = ~(layer_3[768] & layer_3[773]); 
    assign layer_4[760] = ~layer_3[772]; 
    assign layer_4[761] = ~layer_3[746] | (layer_3[772] & layer_3[746]); 
    assign layer_4[762] = layer_3[769] & layer_3[764]; 
    assign layer_4[763] = layer_3[761]; 
    assign layer_4[764] = ~layer_3[779]; 
    assign layer_4[765] = ~layer_3[754] | (layer_3[758] & layer_3[754]); 
    assign layer_4[766] = ~(layer_3[763] ^ layer_3[776]); 
    assign layer_4[767] = layer_3[779] ^ layer_3[771]; 
    assign layer_4[768] = layer_3[767] | layer_3[767]; 
    assign layer_4[769] = ~(layer_3[779] | layer_3[752]); 
    assign layer_4[770] = layer_3[763]; 
    assign layer_4[771] = layer_3[761]; 
    assign layer_4[772] = 1'b1; 
    assign layer_4[773] = ~layer_3[766] | (layer_3[766] & layer_3[765]); 
    assign layer_4[774] = layer_3[758]; 
    assign layer_4[775] = ~layer_3[784] | (layer_3[787] & layer_3[784]); 
    assign layer_4[776] = ~(layer_3[790] ^ layer_3[772]); 
    assign layer_4[777] = ~(layer_3[792] ^ layer_3[773]); 
    assign layer_4[778] = layer_3[780]; 
    assign layer_4[779] = ~(layer_3[786] ^ layer_3[789]); 
    assign layer_4[780] = ~layer_3[778] | (layer_3[778] & layer_3[767]); 
    assign layer_4[781] = ~layer_3[767] | (layer_3[778] & layer_3[767]); 
    assign layer_4[782] = ~layer_3[794]; 
    assign layer_4[783] = ~(layer_3[776] | layer_3[781]); 
    assign layer_4[784] = layer_3[774] | layer_3[791]; 
    assign layer_4[785] = ~(layer_3[769] | layer_3[793]); 
    assign layer_4[786] = ~(layer_3[786] ^ layer_3[778]); 
    assign layer_4[787] = ~layer_3[785] | (layer_3[789] & layer_3[785]); 
    assign layer_4[788] = layer_3[777] & ~layer_3[802]; 
    assign layer_4[789] = layer_3[796] & layer_3[790]; 
    assign layer_4[790] = layer_3[790]; 
    assign layer_4[791] = layer_3[781]; 
    assign layer_4[792] = ~(layer_3[795] ^ layer_3[776]); 
    assign layer_4[793] = layer_3[806] & ~layer_3[785]; 
    assign layer_4[794] = layer_3[795] & ~layer_3[795]; 
    assign layer_4[795] = ~(layer_3[806] ^ layer_3[810]); 
    assign layer_4[796] = ~layer_3[796]; 
    assign layer_4[797] = layer_3[808]; 
    assign layer_4[798] = ~(layer_3[784] | layer_3[790]); 
    assign layer_4[799] = ~(layer_3[804] | layer_3[804]); 
    assign layer_4[800] = ~layer_3[810] | (layer_3[810] & layer_3[813]); 
    assign layer_4[801] = layer_3[810] ^ layer_3[789]; 
    assign layer_4[802] = ~layer_3[811] | (layer_3[811] & layer_3[807]); 
    assign layer_4[803] = layer_3[793] & ~layer_3[787]; 
    assign layer_4[804] = ~layer_3[788] | (layer_3[807] & layer_3[788]); 
    assign layer_4[805] = 1'b0; 
    assign layer_4[806] = ~(layer_3[797] & layer_3[808]); 
    assign layer_4[807] = layer_3[802] | layer_3[809]; 
    assign layer_4[808] = ~(layer_3[795] | layer_3[802]); 
    assign layer_4[809] = ~layer_3[819]; 
    assign layer_4[810] = ~layer_3[806]; 
    assign layer_4[811] = 1'b1; 
    assign layer_4[812] = layer_3[799] & layer_3[800]; 
    assign layer_4[813] = ~layer_3[827] | (layer_3[827] & layer_3[817]); 
    assign layer_4[814] = 1'b0; 
    assign layer_4[815] = layer_3[814]; 
    assign layer_4[816] = layer_3[806]; 
    assign layer_4[817] = layer_3[823]; 
    assign layer_4[818] = ~layer_3[805] | (layer_3[805] & layer_3[822]); 
    assign layer_4[819] = layer_3[824] & ~layer_3[824]; 
    assign layer_4[820] = ~layer_3[807]; 
    assign layer_4[821] = ~(layer_3[815] ^ layer_3[810]); 
    assign layer_4[822] = 1'b0; 
    assign layer_4[823] = ~layer_3[834]; 
    assign layer_4[824] = 1'b0; 
    assign layer_4[825] = layer_3[824] & ~layer_3[819]; 
    assign layer_4[826] = layer_3[820] & ~layer_3[816]; 
    assign layer_4[827] = layer_3[814] & ~layer_3[818]; 
    assign layer_4[828] = layer_3[813] & ~layer_3[813]; 
    assign layer_4[829] = layer_3[828] & layer_3[837]; 
    assign layer_4[830] = 1'b0; 
    assign layer_4[831] = layer_3[820]; 
    assign layer_4[832] = layer_3[841] & layer_3[815]; 
    assign layer_4[833] = layer_3[827] & ~layer_3[834]; 
    assign layer_4[834] = layer_3[839] | layer_3[831]; 
    assign layer_4[835] = layer_3[849]; 
    assign layer_4[836] = ~layer_3[823] | (layer_3[823] & layer_3[832]); 
    assign layer_4[837] = ~(layer_3[848] & layer_3[833]); 
    assign layer_4[838] = layer_3[834] & ~layer_3[853]; 
    assign layer_4[839] = 1'b0; 
    assign layer_4[840] = ~(layer_3[855] & layer_3[839]); 
    assign layer_4[841] = 1'b1; 
    assign layer_4[842] = ~layer_3[830]; 
    assign layer_4[843] = ~layer_3[849]; 
    assign layer_4[844] = layer_3[856]; 
    assign layer_4[845] = ~(layer_3[830] & layer_3[857]); 
    assign layer_4[846] = layer_3[843] & ~layer_3[833]; 
    assign layer_4[847] = layer_3[848]; 
    assign layer_4[848] = layer_3[856] | layer_3[858]; 
    assign layer_4[849] = layer_3[862] | layer_3[841]; 
    assign layer_4[850] = layer_3[864] | layer_3[852]; 
    assign layer_4[851] = layer_3[836]; 
    assign layer_4[852] = layer_3[839] | layer_3[843]; 
    assign layer_4[853] = ~(layer_3[867] | layer_3[839]); 
    assign layer_4[854] = layer_3[844] & ~layer_3[861]; 
    assign layer_4[855] = layer_3[864] & ~layer_3[842]; 
    assign layer_4[856] = layer_3[854]; 
    assign layer_4[857] = layer_3[851]; 
    assign layer_4[858] = ~(layer_3[861] | layer_3[851]); 
    assign layer_4[859] = ~layer_3[871] | (layer_3[871] & layer_3[846]); 
    assign layer_4[860] = ~layer_3[869]; 
    assign layer_4[861] = layer_3[873] & ~layer_3[847]; 
    assign layer_4[862] = ~layer_3[874]; 
    assign layer_4[863] = layer_3[855] | layer_3[869]; 
    assign layer_4[864] = layer_3[878] ^ layer_3[848]; 
    assign layer_4[865] = layer_3[870] & ~layer_3[875]; 
    assign layer_4[866] = ~(layer_3[882] ^ layer_3[855]); 
    assign layer_4[867] = layer_3[883] | layer_3[855]; 
    assign layer_4[868] = layer_3[870] ^ layer_3[857]; 
    assign layer_4[869] = ~(layer_3[853] ^ layer_3[879]); 
    assign layer_4[870] = ~(layer_3[865] & layer_3[876]); 
    assign layer_4[871] = ~(layer_3[887] ^ layer_3[881]); 
    assign layer_4[872] = ~layer_3[870]; 
    assign layer_4[873] = ~(layer_3[867] ^ layer_3[883]); 
    assign layer_4[874] = layer_3[881] & ~layer_3[873]; 
    assign layer_4[875] = layer_3[883] & ~layer_3[883]; 
    assign layer_4[876] = layer_3[873] & ~layer_3[887]; 
    assign layer_4[877] = layer_3[871] ^ layer_3[885]; 
    assign layer_4[878] = layer_3[872] ^ layer_3[890]; 
    assign layer_4[879] = ~(layer_3[869] | layer_3[884]); 
    assign layer_4[880] = layer_3[863] & ~layer_3[865]; 
    assign layer_4[881] = 1'b1; 
    assign layer_4[882] = layer_3[877] & ~layer_3[879]; 
    assign layer_4[883] = ~layer_3[868] | (layer_3[868] & layer_3[886]); 
    assign layer_4[884] = layer_3[874] & ~layer_3[897]; 
    assign layer_4[885] = ~(layer_3[890] | layer_3[876]); 
    assign layer_4[886] = layer_3[871] & layer_3[872]; 
    assign layer_4[887] = layer_3[889] ^ layer_3[873]; 
    assign layer_4[888] = layer_3[883] ^ layer_3[877]; 
    assign layer_4[889] = 1'b0; 
    assign layer_4[890] = ~layer_3[899]; 
    assign layer_4[891] = ~layer_3[889] | (layer_3[889] & layer_3[900]); 
    assign layer_4[892] = ~(layer_3[896] ^ layer_3[894]); 
    assign layer_4[893] = layer_3[894]; 
    assign layer_4[894] = ~layer_3[892]; 
    assign layer_4[895] = ~layer_3[884] | (layer_3[892] & layer_3[884]); 
    assign layer_4[896] = layer_3[906]; 
    assign layer_4[897] = ~(layer_3[907] & layer_3[907]); 
    assign layer_4[898] = ~layer_3[888]; 
    assign layer_4[899] = 1'b0; 
    assign layer_4[900] = ~layer_3[906]; 
    assign layer_4[901] = layer_3[884] & ~layer_3[900]; 
    assign layer_4[902] = layer_3[915] & ~layer_3[901]; 
    assign layer_4[903] = layer_3[898] & ~layer_3[905]; 
    assign layer_4[904] = ~layer_3[894]; 
    assign layer_4[905] = ~layer_3[905]; 
    assign layer_4[906] = ~layer_3[909]; 
    assign layer_4[907] = layer_3[904]; 
    assign layer_4[908] = layer_3[919] & ~layer_3[893]; 
    assign layer_4[909] = layer_3[908]; 
    assign layer_4[910] = ~(layer_3[902] ^ layer_3[903]); 
    assign layer_4[911] = ~(layer_3[899] ^ layer_3[904]); 
    assign layer_4[912] = ~layer_3[920] | (layer_3[920] & layer_3[922]); 
    assign layer_4[913] = ~layer_3[904] | (layer_3[904] & layer_3[919]); 
    assign layer_4[914] = layer_3[904] & ~layer_3[905]; 
    assign layer_4[915] = layer_3[913] & ~layer_3[904]; 
    assign layer_4[916] = layer_3[922] & ~layer_3[925]; 
    assign layer_4[917] = layer_3[904] | layer_3[909]; 
    assign layer_4[918] = ~(layer_3[930] | layer_3[914]); 
    assign layer_4[919] = ~layer_3[926] | (layer_3[924] & layer_3[926]); 
    assign layer_4[920] = ~layer_3[932] | (layer_3[934] & layer_3[932]); 
    assign layer_4[921] = layer_3[924] & ~layer_3[917]; 
    assign layer_4[922] = ~(layer_3[911] ^ layer_3[928]); 
    assign layer_4[923] = layer_3[909] & ~layer_3[914]; 
    assign layer_4[924] = ~(layer_3[922] | layer_3[933]); 
    assign layer_4[925] = ~(layer_3[909] | layer_3[917]); 
    assign layer_4[926] = layer_3[941]; 
    assign layer_4[927] = layer_3[912]; 
    assign layer_4[928] = ~(layer_3[944] ^ layer_3[940]); 
    assign layer_4[929] = ~(layer_3[917] | layer_3[941]); 
    assign layer_4[930] = layer_3[918] & ~layer_3[916]; 
    assign layer_4[931] = layer_3[927] & ~layer_3[929]; 
    assign layer_4[932] = 1'b1; 
    assign layer_4[933] = ~(layer_3[948] ^ layer_3[918]); 
    assign layer_4[934] = 1'b1; 
    assign layer_4[935] = ~(layer_3[946] & layer_3[945]); 
    assign layer_4[936] = ~layer_3[929] | (layer_3[945] & layer_3[929]); 
    assign layer_4[937] = layer_3[946]; 
    assign layer_4[938] = layer_3[952] & ~layer_3[950]; 
    assign layer_4[939] = layer_3[933] & ~layer_3[942]; 
    assign layer_4[940] = ~layer_3[932] | (layer_3[932] & layer_3[954]); 
    assign layer_4[941] = layer_3[947] & layer_3[925]; 
    assign layer_4[942] = ~layer_3[955] | (layer_3[934] & layer_3[955]); 
    assign layer_4[943] = ~layer_3[936]; 
    assign layer_4[944] = ~layer_3[948] | (layer_3[948] & layer_3[953]); 
    assign layer_4[945] = ~layer_3[956]; 
    assign layer_4[946] = ~(layer_3[939] | layer_3[959]); 
    assign layer_4[947] = layer_3[963] & layer_3[940]; 
    assign layer_4[948] = ~layer_3[941]; 
    assign layer_4[949] = layer_3[937] | layer_3[936]; 
    assign layer_4[950] = layer_3[940] | layer_3[962]; 
    assign layer_4[951] = layer_3[961] & ~layer_3[950]; 
    assign layer_4[952] = ~layer_3[955]; 
    assign layer_4[953] = 1'b0; 
    assign layer_4[954] = layer_3[948]; 
    assign layer_4[955] = 1'b1; 
    assign layer_4[956] = layer_3[969] & layer_3[947]; 
    assign layer_4[957] = layer_3[965] ^ layer_3[943]; 
    assign layer_4[958] = layer_3[953] | layer_3[942]; 
    assign layer_4[959] = ~(layer_3[955] | layer_3[967]); 
    assign layer_4[960] = layer_3[955] & ~layer_3[947]; 
    assign layer_4[961] = layer_3[970] ^ layer_3[957]; 
    assign layer_4[962] = ~layer_3[953]; 
    assign layer_4[963] = layer_3[977] ^ layer_3[949]; 
    assign layer_4[964] = ~layer_3[977] | (layer_3[980] & layer_3[977]); 
    assign layer_4[965] = layer_3[959]; 
    assign layer_4[966] = layer_3[968] & layer_3[976]; 
    assign layer_4[967] = ~layer_3[982]; 
    assign layer_4[968] = 1'b1; 
    assign layer_4[969] = layer_3[979] & ~layer_3[979]; 
    assign layer_4[970] = ~layer_3[971] | (layer_3[971] & layer_3[966]); 
    assign layer_4[971] = ~layer_3[955]; 
    assign layer_4[972] = layer_3[973]; 
    assign layer_4[973] = layer_3[976] & ~layer_3[961]; 
    assign layer_4[974] = layer_3[974] ^ layer_3[971]; 
    assign layer_4[975] = layer_3[986] | layer_3[981]; 
    assign layer_4[976] = layer_3[965] & ~layer_3[984]; 
    assign layer_4[977] = layer_3[968] | layer_3[983]; 
    assign layer_4[978] = layer_3[974] & ~layer_3[962]; 
    assign layer_4[979] = layer_3[978]; 
    assign layer_4[980] = ~(layer_3[972] | layer_3[987]); 
    assign layer_4[981] = 1'b1; 
    assign layer_4[982] = layer_3[997] & ~layer_3[995]; 
    assign layer_4[983] = ~layer_3[968]; 
    assign layer_4[984] = layer_3[994] ^ layer_3[997]; 
    assign layer_4[985] = 1'b1; 
    assign layer_4[986] = ~layer_3[995]; 
    assign layer_4[987] = ~layer_3[981]; 
    assign layer_4[988] = layer_3[987] & ~layer_3[1003]; 
    assign layer_4[989] = 1'b1; 
    assign layer_4[990] = 1'b0; 
    assign layer_4[991] = ~layer_3[1000] | (layer_3[993] & layer_3[1000]); 
    assign layer_4[992] = layer_3[991]; 
    assign layer_4[993] = ~layer_3[994] | (layer_3[994] & layer_3[985]); 
    assign layer_4[994] = layer_3[989] & layer_3[987]; 
    assign layer_4[995] = layer_3[986] & ~layer_3[979]; 
    assign layer_4[996] = layer_3[1002] & layer_3[1000]; 
    assign layer_4[997] = layer_3[1004] | layer_3[980]; 
    assign layer_4[998] = ~layer_3[1005] | (layer_3[1006] & layer_3[1005]); 
    assign layer_4[999] = ~layer_3[985] | (layer_3[985] & layer_3[985]); 
    assign layer_4[1000] = layer_3[1014] & ~layer_3[1001]; 
    assign layer_4[1001] = 1'b0; 
    assign layer_4[1002] = ~(layer_3[987] ^ layer_3[1017]); 
    assign layer_4[1003] = ~layer_3[987] | (layer_3[1009] & layer_3[987]); 
    assign layer_4[1004] = 1'b1; 
    assign layer_4[1005] = layer_3[997]; 
    assign layer_4[1006] = layer_3[1009] & ~layer_3[999]; 
    assign layer_4[1007] = ~layer_3[1001] | (layer_3[1001] & layer_3[999]); 
    assign layer_4[1008] = layer_3[1021] ^ layer_3[1009]; 
    assign layer_4[1009] = layer_3[1014] & ~layer_3[1000]; 
    assign layer_4[1010] = layer_3[1014] | layer_3[1011]; 
    assign layer_4[1011] = layer_3[1001] & ~layer_3[997]; 
    assign layer_4[1012] = layer_3[1002]; 
    assign layer_4[1013] = 1'b1; 
    assign layer_4[1014] = ~layer_3[1005]; 
    assign layer_4[1015] = layer_3[1017] & ~layer_3[1003]; 
    assign layer_4[1016] = ~layer_3[1019] | (layer_3[1023] & layer_3[1019]); 
    assign layer_4[1017] = layer_3[1015]; 
    assign layer_4[1018] = 1'b1; 
    assign layer_4[1019] = ~(layer_3[1014] ^ layer_3[1011]); 
    assign layer_4[1020] = layer_3[1013] & ~layer_3[1022]; 
    assign layer_4[1021] = layer_3[1005]; 
    assign layer_4[1022] = layer_3[1015]; 
    assign layer_4[1023] = ~(layer_3[1008] ^ layer_3[1021]); 
    // Layer 5 ============================================================
    assign layer_5[0] = ~layer_4[14] | (layer_4[14] & layer_4[9]); 
    assign layer_5[1] = ~layer_4[4]; 
    assign layer_5[2] = ~(layer_4[17] & layer_4[0]); 
    assign layer_5[3] = layer_4[9] & ~layer_4[2]; 
    assign layer_5[4] = ~layer_4[11]; 
    assign layer_5[5] = 1'b1; 
    assign layer_5[6] = ~(layer_4[14] | layer_4[5]); 
    assign layer_5[7] = ~(layer_4[15] ^ layer_4[6]); 
    assign layer_5[8] = 1'b0; 
    assign layer_5[9] = ~(layer_4[3] & layer_4[8]); 
    assign layer_5[10] = ~layer_4[9] | (layer_4[13] & layer_4[9]); 
    assign layer_5[11] = layer_4[3]; 
    assign layer_5[12] = 1'b0; 
    assign layer_5[13] = ~layer_4[3] | (layer_4[21] & layer_4[3]); 
    assign layer_5[14] = 1'b0; 
    assign layer_5[15] = ~layer_4[30]; 
    assign layer_5[16] = 1'b1; 
    assign layer_5[17] = ~layer_4[5] | (layer_4[5] & layer_4[20]); 
    assign layer_5[18] = layer_4[5] & layer_4[9]; 
    assign layer_5[19] = layer_4[17] & layer_4[14]; 
    assign layer_5[20] = ~layer_4[10] | (layer_4[10] & layer_4[22]); 
    assign layer_5[21] = ~(layer_4[23] & layer_4[27]); 
    assign layer_5[22] = ~layer_4[24]; 
    assign layer_5[23] = ~(layer_4[38] ^ layer_4[33]); 
    assign layer_5[24] = layer_4[11] & ~layer_4[13]; 
    assign layer_5[25] = layer_4[10]; 
    assign layer_5[26] = layer_4[24]; 
    assign layer_5[27] = ~(layer_4[14] | layer_4[20]); 
    assign layer_5[28] = layer_4[21] ^ layer_4[40]; 
    assign layer_5[29] = layer_4[14]; 
    assign layer_5[30] = ~layer_4[37] | (layer_4[19] & layer_4[37]); 
    assign layer_5[31] = ~(layer_4[28] ^ layer_4[31]); 
    assign layer_5[32] = ~(layer_4[43] ^ layer_4[27]); 
    assign layer_5[33] = layer_4[44] | layer_4[37]; 
    assign layer_5[34] = ~layer_4[29] | (layer_4[29] & layer_4[25]); 
    assign layer_5[35] = layer_4[29] & ~layer_4[32]; 
    assign layer_5[36] = ~(layer_4[22] ^ layer_4[30]); 
    assign layer_5[37] = layer_4[30] & ~layer_4[24]; 
    assign layer_5[38] = layer_4[45] & ~layer_4[28]; 
    assign layer_5[39] = layer_4[26] & ~layer_4[46]; 
    assign layer_5[40] = layer_4[50] | layer_4[23]; 
    assign layer_5[41] = layer_4[26]; 
    assign layer_5[42] = ~(layer_4[52] & layer_4[50]); 
    assign layer_5[43] = ~layer_4[41] | (layer_4[51] & layer_4[41]); 
    assign layer_5[44] = layer_4[40] | layer_4[52]; 
    assign layer_5[45] = ~(layer_4[30] ^ layer_4[37]); 
    assign layer_5[46] = ~(layer_4[32] ^ layer_4[50]); 
    assign layer_5[47] = ~layer_4[61] | (layer_4[61] & layer_4[53]); 
    assign layer_5[48] = layer_4[45] & ~layer_4[45]; 
    assign layer_5[49] = ~layer_4[53]; 
    assign layer_5[50] = ~(layer_4[47] | layer_4[38]); 
    assign layer_5[51] = ~(layer_4[40] | layer_4[66]); 
    assign layer_5[52] = ~layer_4[41]; 
    assign layer_5[53] = ~layer_4[63] | (layer_4[62] & layer_4[63]); 
    assign layer_5[54] = layer_4[46] & ~layer_4[54]; 
    assign layer_5[55] = layer_4[60] | layer_4[42]; 
    assign layer_5[56] = ~layer_4[70] | (layer_4[70] & layer_4[43]); 
    assign layer_5[57] = layer_4[59]; 
    assign layer_5[58] = layer_4[49] & ~layer_4[60]; 
    assign layer_5[59] = ~layer_4[69] | (layer_4[69] & layer_4[72]); 
    assign layer_5[60] = layer_4[73]; 
    assign layer_5[61] = ~layer_4[68]; 
    assign layer_5[62] = 1'b1; 
    assign layer_5[63] = ~(layer_4[67] & layer_4[62]); 
    assign layer_5[64] = layer_4[61] & ~layer_4[51]; 
    assign layer_5[65] = layer_4[58] ^ layer_4[51]; 
    assign layer_5[66] = layer_4[56] | layer_4[61]; 
    assign layer_5[67] = layer_4[56] & ~layer_4[58]; 
    assign layer_5[68] = layer_4[58]; 
    assign layer_5[69] = 1'b0; 
    assign layer_5[70] = ~layer_4[70]; 
    assign layer_5[71] = layer_4[56] & ~layer_4[64]; 
    assign layer_5[72] = layer_4[72] & ~layer_4[60]; 
    assign layer_5[73] = layer_4[84] ^ layer_4[79]; 
    assign layer_5[74] = layer_4[72] | layer_4[76]; 
    assign layer_5[75] = layer_4[69] & ~layer_4[66]; 
    assign layer_5[76] = ~layer_4[64] | (layer_4[70] & layer_4[64]); 
    assign layer_5[77] = layer_4[68] & layer_4[74]; 
    assign layer_5[78] = layer_4[80] ^ layer_4[73]; 
    assign layer_5[79] = layer_4[92] ^ layer_4[75]; 
    assign layer_5[80] = layer_4[67] ^ layer_4[71]; 
    assign layer_5[81] = ~layer_4[90]; 
    assign layer_5[82] = layer_4[80] & ~layer_4[85]; 
    assign layer_5[83] = 1'b0; 
    assign layer_5[84] = layer_4[81] ^ layer_4[85]; 
    assign layer_5[85] = 1'b1; 
    assign layer_5[86] = ~(layer_4[75] & layer_4[84]); 
    assign layer_5[87] = ~layer_4[77]; 
    assign layer_5[88] = layer_4[73] & ~layer_4[98]; 
    assign layer_5[89] = layer_4[81] & ~layer_4[78]; 
    assign layer_5[90] = layer_4[88] & ~layer_4[84]; 
    assign layer_5[91] = ~(layer_4[105] & layer_4[106]); 
    assign layer_5[92] = 1'b0; 
    assign layer_5[93] = layer_4[107] & ~layer_4[86]; 
    assign layer_5[94] = ~layer_4[89]; 
    assign layer_5[95] = layer_4[102] & ~layer_4[111]; 
    assign layer_5[96] = ~(layer_4[99] ^ layer_4[86]); 
    assign layer_5[97] = ~(layer_4[91] & layer_4[87]); 
    assign layer_5[98] = 1'b0; 
    assign layer_5[99] = 1'b1; 
    assign layer_5[100] = ~layer_4[97]; 
    assign layer_5[101] = ~layer_4[116] | (layer_4[107] & layer_4[116]); 
    assign layer_5[102] = ~layer_4[96]; 
    assign layer_5[103] = ~layer_4[108]; 
    assign layer_5[104] = layer_4[115] & ~layer_4[119]; 
    assign layer_5[105] = 1'b1; 
    assign layer_5[106] = layer_4[101]; 
    assign layer_5[107] = 1'b1; 
    assign layer_5[108] = layer_4[94] | layer_4[105]; 
    assign layer_5[109] = layer_4[120] | layer_4[121]; 
    assign layer_5[110] = layer_4[114]; 
    assign layer_5[111] = layer_4[104]; 
    assign layer_5[112] = layer_4[106] & ~layer_4[102]; 
    assign layer_5[113] = ~layer_4[102] | (layer_4[113] & layer_4[102]); 
    assign layer_5[114] = layer_4[123] & layer_4[113]; 
    assign layer_5[115] = 1'b0; 
    assign layer_5[116] = 1'b1; 
    assign layer_5[117] = ~layer_4[110]; 
    assign layer_5[118] = ~(layer_4[132] | layer_4[124]); 
    assign layer_5[119] = ~(layer_4[124] ^ layer_4[119]); 
    assign layer_5[120] = 1'b1; 
    assign layer_5[121] = ~layer_4[130] | (layer_4[132] & layer_4[130]); 
    assign layer_5[122] = ~layer_4[132] | (layer_4[132] & layer_4[127]); 
    assign layer_5[123] = ~(layer_4[135] ^ layer_4[113]); 
    assign layer_5[124] = layer_4[119] & layer_4[134]; 
    assign layer_5[125] = layer_4[135] & layer_4[134]; 
    assign layer_5[126] = ~layer_4[135] | (layer_4[135] & layer_4[135]); 
    assign layer_5[127] = 1'b0; 
    assign layer_5[128] = 1'b1; 
    assign layer_5[129] = layer_4[130] | layer_4[120]; 
    assign layer_5[130] = ~(layer_4[115] ^ layer_4[127]); 
    assign layer_5[131] = ~(layer_4[136] ^ layer_4[118]); 
    assign layer_5[132] = ~layer_4[143] | (layer_4[143] & layer_4[139]); 
    assign layer_5[133] = layer_4[123] & layer_4[128]; 
    assign layer_5[134] = ~(layer_4[127] ^ layer_4[120]); 
    assign layer_5[135] = layer_4[149] & ~layer_4[120]; 
    assign layer_5[136] = ~(layer_4[151] | layer_4[144]); 
    assign layer_5[137] = ~(layer_4[151] | layer_4[147]); 
    assign layer_5[138] = layer_4[142]; 
    assign layer_5[139] = ~layer_4[154]; 
    assign layer_5[140] = ~layer_4[133]; 
    assign layer_5[141] = ~layer_4[137] | (layer_4[137] & layer_4[124]); 
    assign layer_5[142] = layer_4[138] | layer_4[151]; 
    assign layer_5[143] = layer_4[138]; 
    assign layer_5[144] = layer_4[140] ^ layer_4[131]; 
    assign layer_5[145] = layer_4[148]; 
    assign layer_5[146] = ~layer_4[147]; 
    assign layer_5[147] = layer_4[133] | layer_4[147]; 
    assign layer_5[148] = ~layer_4[153]; 
    assign layer_5[149] = ~layer_4[132] | (layer_4[134] & layer_4[132]); 
    assign layer_5[150] = ~layer_4[153] | (layer_4[149] & layer_4[153]); 
    assign layer_5[151] = ~(layer_4[165] ^ layer_4[151]); 
    assign layer_5[152] = layer_4[167]; 
    assign layer_5[153] = 1'b1; 
    assign layer_5[154] = ~(layer_4[148] ^ layer_4[168]); 
    assign layer_5[155] = ~(layer_4[153] ^ layer_4[149]); 
    assign layer_5[156] = layer_4[146] & ~layer_4[158]; 
    assign layer_5[157] = layer_4[154] | layer_4[156]; 
    assign layer_5[158] = layer_4[173] ^ layer_4[168]; 
    assign layer_5[159] = layer_4[166] & ~layer_4[158]; 
    assign layer_5[160] = ~layer_4[176] | (layer_4[176] & layer_4[151]); 
    assign layer_5[161] = ~layer_4[172] | (layer_4[172] & layer_4[153]); 
    assign layer_5[162] = 1'b1; 
    assign layer_5[163] = layer_4[157] & ~layer_4[162]; 
    assign layer_5[164] = ~(layer_4[179] | layer_4[167]); 
    assign layer_5[165] = layer_4[178] & layer_4[164]; 
    assign layer_5[166] = ~(layer_4[168] & layer_4[167]); 
    assign layer_5[167] = layer_4[168]; 
    assign layer_5[168] = layer_4[162] & ~layer_4[168]; 
    assign layer_5[169] = 1'b0; 
    assign layer_5[170] = ~layer_4[170]; 
    assign layer_5[171] = layer_4[183]; 
    assign layer_5[172] = layer_4[168] | layer_4[181]; 
    assign layer_5[173] = layer_4[173] & ~layer_4[157]; 
    assign layer_5[174] = ~(layer_4[184] | layer_4[183]); 
    assign layer_5[175] = ~(layer_4[169] | layer_4[167]); 
    assign layer_5[176] = ~(layer_4[178] | layer_4[173]); 
    assign layer_5[177] = layer_4[191] & ~layer_4[164]; 
    assign layer_5[178] = ~(layer_4[165] ^ layer_4[163]); 
    assign layer_5[179] = layer_4[182] & ~layer_4[167]; 
    assign layer_5[180] = ~layer_4[172] | (layer_4[182] & layer_4[172]); 
    assign layer_5[181] = ~layer_4[175]; 
    assign layer_5[182] = ~layer_4[177]; 
    assign layer_5[183] = layer_4[179] ^ layer_4[176]; 
    assign layer_5[184] = ~layer_4[184] | (layer_4[168] & layer_4[184]); 
    assign layer_5[185] = 1'b0; 
    assign layer_5[186] = ~(layer_4[183] | layer_4[182]); 
    assign layer_5[187] = ~layer_4[174]; 
    assign layer_5[188] = layer_4[178]; 
    assign layer_5[189] = ~(layer_4[175] | layer_4[201]); 
    assign layer_5[190] = ~layer_4[184]; 
    assign layer_5[191] = layer_4[188] & ~layer_4[203]; 
    assign layer_5[192] = ~layer_4[203]; 
    assign layer_5[193] = layer_4[206] & layer_4[198]; 
    assign layer_5[194] = ~layer_4[209]; 
    assign layer_5[195] = ~layer_4[192] | (layer_4[192] & layer_4[207]); 
    assign layer_5[196] = layer_4[208] & layer_4[195]; 
    assign layer_5[197] = ~(layer_4[201] ^ layer_4[196]); 
    assign layer_5[198] = ~(layer_4[206] ^ layer_4[209]); 
    assign layer_5[199] = layer_4[192] ^ layer_4[198]; 
    assign layer_5[200] = layer_4[190]; 
    assign layer_5[201] = 1'b0; 
    assign layer_5[202] = ~(layer_4[203] ^ layer_4[189]); 
    assign layer_5[203] = ~(layer_4[204] | layer_4[186]); 
    assign layer_5[204] = ~layer_4[194]; 
    assign layer_5[205] = layer_4[191] ^ layer_4[219]; 
    assign layer_5[206] = layer_4[191] | layer_4[218]; 
    assign layer_5[207] = 1'b1; 
    assign layer_5[208] = layer_4[195] & ~layer_4[203]; 
    assign layer_5[209] = ~layer_4[199]; 
    assign layer_5[210] = 1'b0; 
    assign layer_5[211] = layer_4[218]; 
    assign layer_5[212] = ~(layer_4[224] | layer_4[226]); 
    assign layer_5[213] = ~layer_4[212] | (layer_4[202] & layer_4[212]); 
    assign layer_5[214] = layer_4[206] & layer_4[218]; 
    assign layer_5[215] = layer_4[227] & ~layer_4[204]; 
    assign layer_5[216] = layer_4[217]; 
    assign layer_5[217] = layer_4[203] & ~layer_4[224]; 
    assign layer_5[218] = ~layer_4[231]; 
    assign layer_5[219] = ~layer_4[232]; 
    assign layer_5[220] = layer_4[210] & ~layer_4[224]; 
    assign layer_5[221] = 1'b1; 
    assign layer_5[222] = layer_4[220]; 
    assign layer_5[223] = layer_4[214] & ~layer_4[229]; 
    assign layer_5[224] = layer_4[219]; 
    assign layer_5[225] = layer_4[219]; 
    assign layer_5[226] = ~layer_4[225] | (layer_4[240] & layer_4[225]); 
    assign layer_5[227] = layer_4[230] & layer_4[235]; 
    assign layer_5[228] = layer_4[213]; 
    assign layer_5[229] = layer_4[235] & ~layer_4[214]; 
    assign layer_5[230] = ~layer_4[220] | (layer_4[242] & layer_4[220]); 
    assign layer_5[231] = layer_4[231] & ~layer_4[221]; 
    assign layer_5[232] = ~layer_4[229]; 
    assign layer_5[233] = layer_4[220] & ~layer_4[243]; 
    assign layer_5[234] = ~(layer_4[250] & layer_4[244]); 
    assign layer_5[235] = ~layer_4[218]; 
    assign layer_5[236] = 1'b1; 
    assign layer_5[237] = layer_4[225]; 
    assign layer_5[238] = layer_4[244] | layer_4[228]; 
    assign layer_5[239] = layer_4[246]; 
    assign layer_5[240] = ~(layer_4[251] | layer_4[239]); 
    assign layer_5[241] = ~(layer_4[242] ^ layer_4[241]); 
    assign layer_5[242] = 1'b0; 
    assign layer_5[243] = layer_4[241] | layer_4[229]; 
    assign layer_5[244] = 1'b0; 
    assign layer_5[245] = layer_4[253]; 
    assign layer_5[246] = ~layer_4[236] | (layer_4[233] & layer_4[236]); 
    assign layer_5[247] = layer_4[252] & ~layer_4[242]; 
    assign layer_5[248] = ~layer_4[258]; 
    assign layer_5[249] = ~(layer_4[239] | layer_4[253]); 
    assign layer_5[250] = layer_4[247] & ~layer_4[263]; 
    assign layer_5[251] = layer_4[246] & ~layer_4[250]; 
    assign layer_5[252] = layer_4[236] | layer_4[245]; 
    assign layer_5[253] = layer_4[263] | layer_4[259]; 
    assign layer_5[254] = ~(layer_4[244] & layer_4[252]); 
    assign layer_5[255] = ~(layer_4[262] | layer_4[242]); 
    assign layer_5[256] = layer_4[244] & ~layer_4[265]; 
    assign layer_5[257] = ~layer_4[241]; 
    assign layer_5[258] = ~(layer_4[245] | layer_4[261]); 
    assign layer_5[259] = ~layer_4[250]; 
    assign layer_5[260] = ~layer_4[268]; 
    assign layer_5[261] = layer_4[250] | layer_4[251]; 
    assign layer_5[262] = layer_4[249] ^ layer_4[275]; 
    assign layer_5[263] = layer_4[273]; 
    assign layer_5[264] = ~layer_4[254] | (layer_4[254] & layer_4[248]); 
    assign layer_5[265] = layer_4[280] & layer_4[278]; 
    assign layer_5[266] = layer_4[251] & ~layer_4[272]; 
    assign layer_5[267] = layer_4[274]; 
    assign layer_5[268] = ~layer_4[279]; 
    assign layer_5[269] = ~layer_4[268] | (layer_4[268] & layer_4[263]); 
    assign layer_5[270] = ~(layer_4[279] | layer_4[279]); 
    assign layer_5[271] = layer_4[262] ^ layer_4[283]; 
    assign layer_5[272] = ~layer_4[261]; 
    assign layer_5[273] = ~(layer_4[286] & layer_4[259]); 
    assign layer_5[274] = ~layer_4[260]; 
    assign layer_5[275] = layer_4[282] & ~layer_4[271]; 
    assign layer_5[276] = 1'b0; 
    assign layer_5[277] = ~layer_4[287]; 
    assign layer_5[278] = layer_4[290] & ~layer_4[265]; 
    assign layer_5[279] = ~(layer_4[283] & layer_4[276]); 
    assign layer_5[280] = layer_4[290]; 
    assign layer_5[281] = 1'b0; 
    assign layer_5[282] = layer_4[280]; 
    assign layer_5[283] = layer_4[298]; 
    assign layer_5[284] = ~(layer_4[275] & layer_4[275]); 
    assign layer_5[285] = layer_4[272] ^ layer_4[280]; 
    assign layer_5[286] = layer_4[276] ^ layer_4[289]; 
    assign layer_5[287] = layer_4[280] ^ layer_4[273]; 
    assign layer_5[288] = ~layer_4[284]; 
    assign layer_5[289] = layer_4[286] | layer_4[298]; 
    assign layer_5[290] = layer_4[282]; 
    assign layer_5[291] = ~layer_4[301] | (layer_4[283] & layer_4[301]); 
    assign layer_5[292] = layer_4[282] | layer_4[300]; 
    assign layer_5[293] = layer_4[298] & layer_4[290]; 
    assign layer_5[294] = 1'b1; 
    assign layer_5[295] = ~layer_4[302] | (layer_4[291] & layer_4[302]); 
    assign layer_5[296] = layer_4[290]; 
    assign layer_5[297] = ~layer_4[300] | (layer_4[300] & layer_4[294]); 
    assign layer_5[298] = ~layer_4[291] | (layer_4[306] & layer_4[291]); 
    assign layer_5[299] = ~layer_4[294]; 
    assign layer_5[300] = ~(layer_4[292] | layer_4[300]); 
    assign layer_5[301] = layer_4[296] & ~layer_4[292]; 
    assign layer_5[302] = ~layer_4[285] | (layer_4[289] & layer_4[285]); 
    assign layer_5[303] = ~(layer_4[299] ^ layer_4[318]); 
    assign layer_5[304] = layer_4[315] & ~layer_4[313]; 
    assign layer_5[305] = ~(layer_4[312] | layer_4[290]); 
    assign layer_5[306] = layer_4[292] & ~layer_4[318]; 
    assign layer_5[307] = ~(layer_4[292] | layer_4[301]); 
    assign layer_5[308] = ~layer_4[323] | (layer_4[302] & layer_4[323]); 
    assign layer_5[309] = layer_4[293] & layer_4[302]; 
    assign layer_5[310] = layer_4[302] & layer_4[300]; 
    assign layer_5[311] = layer_4[319] & layer_4[324]; 
    assign layer_5[312] = ~(layer_4[314] & layer_4[296]); 
    assign layer_5[313] = ~layer_4[309] | (layer_4[309] & layer_4[316]); 
    assign layer_5[314] = 1'b1; 
    assign layer_5[315] = ~layer_4[326] | (layer_4[326] & layer_4[321]); 
    assign layer_5[316] = ~(layer_4[301] | layer_4[308]); 
    assign layer_5[317] = layer_4[309]; 
    assign layer_5[318] = ~layer_4[305]; 
    assign layer_5[319] = ~layer_4[307] | (layer_4[330] & layer_4[307]); 
    assign layer_5[320] = layer_4[327] ^ layer_4[312]; 
    assign layer_5[321] = layer_4[312] & ~layer_4[316]; 
    assign layer_5[322] = ~layer_4[319]; 
    assign layer_5[323] = ~layer_4[326] | (layer_4[326] & layer_4[329]); 
    assign layer_5[324] = layer_4[318] | layer_4[323]; 
    assign layer_5[325] = layer_4[325]; 
    assign layer_5[326] = ~(layer_4[311] & layer_4[319]); 
    assign layer_5[327] = ~layer_4[330] | (layer_4[330] & layer_4[318]); 
    assign layer_5[328] = layer_4[325] & layer_4[341]; 
    assign layer_5[329] = ~(layer_4[338] & layer_4[320]); 
    assign layer_5[330] = 1'b0; 
    assign layer_5[331] = layer_4[329] & ~layer_4[345]; 
    assign layer_5[332] = ~layer_4[335]; 
    assign layer_5[333] = 1'b0; 
    assign layer_5[334] = layer_4[336]; 
    assign layer_5[335] = ~(layer_4[338] | layer_4[337]); 
    assign layer_5[336] = layer_4[348]; 
    assign layer_5[337] = layer_4[347] & ~layer_4[348]; 
    assign layer_5[338] = layer_4[322] & ~layer_4[351]; 
    assign layer_5[339] = ~(layer_4[336] ^ layer_4[345]); 
    assign layer_5[340] = ~(layer_4[333] ^ layer_4[323]); 
    assign layer_5[341] = ~layer_4[341]; 
    assign layer_5[342] = layer_4[350]; 
    assign layer_5[343] = layer_4[335] & ~layer_4[330]; 
    assign layer_5[344] = layer_4[329] ^ layer_4[327]; 
    assign layer_5[345] = ~layer_4[338]; 
    assign layer_5[346] = ~(layer_4[361] & layer_4[336]); 
    assign layer_5[347] = ~(layer_4[363] & layer_4[340]); 
    assign layer_5[348] = layer_4[348] & layer_4[339]; 
    assign layer_5[349] = ~layer_4[334]; 
    assign layer_5[350] = ~(layer_4[343] | layer_4[338]); 
    assign layer_5[351] = layer_4[346]; 
    assign layer_5[352] = layer_4[336] & layer_4[340]; 
    assign layer_5[353] = layer_4[367] & layer_4[349]; 
    assign layer_5[354] = layer_4[346]; 
    assign layer_5[355] = layer_4[358] ^ layer_4[343]; 
    assign layer_5[356] = ~(layer_4[365] | layer_4[359]); 
    assign layer_5[357] = layer_4[350] & ~layer_4[364]; 
    assign layer_5[358] = ~layer_4[352] | (layer_4[352] & layer_4[352]); 
    assign layer_5[359] = ~(layer_4[373] ^ layer_4[352]); 
    assign layer_5[360] = 1'b1; 
    assign layer_5[361] = layer_4[358] ^ layer_4[358]; 
    assign layer_5[362] = ~(layer_4[358] | layer_4[374]); 
    assign layer_5[363] = 1'b1; 
    assign layer_5[364] = layer_4[359]; 
    assign layer_5[365] = layer_4[360] ^ layer_4[348]; 
    assign layer_5[366] = layer_4[352]; 
    assign layer_5[367] = layer_4[361]; 
    assign layer_5[368] = layer_4[370] | layer_4[367]; 
    assign layer_5[369] = layer_4[379] | layer_4[358]; 
    assign layer_5[370] = 1'b0; 
    assign layer_5[371] = layer_4[376] & ~layer_4[365]; 
    assign layer_5[372] = layer_4[371] | layer_4[375]; 
    assign layer_5[373] = ~layer_4[364] | (layer_4[389] & layer_4[364]); 
    assign layer_5[374] = layer_4[380]; 
    assign layer_5[375] = 1'b1; 
    assign layer_5[376] = ~(layer_4[367] & layer_4[362]); 
    assign layer_5[377] = layer_4[389] & layer_4[360]; 
    assign layer_5[378] = ~(layer_4[362] ^ layer_4[392]); 
    assign layer_5[379] = layer_4[393]; 
    assign layer_5[380] = ~(layer_4[392] | layer_4[388]); 
    assign layer_5[381] = layer_4[375] & layer_4[375]; 
    assign layer_5[382] = ~layer_4[384] | (layer_4[386] & layer_4[384]); 
    assign layer_5[383] = 1'b1; 
    assign layer_5[384] = layer_4[394] & ~layer_4[377]; 
    assign layer_5[385] = layer_4[372] | layer_4[386]; 
    assign layer_5[386] = layer_4[393] & ~layer_4[375]; 
    assign layer_5[387] = layer_4[396] & layer_4[392]; 
    assign layer_5[388] = ~(layer_4[393] & layer_4[382]); 
    assign layer_5[389] = layer_4[373] ^ layer_4[394]; 
    assign layer_5[390] = layer_4[387]; 
    assign layer_5[391] = ~layer_4[406]; 
    assign layer_5[392] = layer_4[403] ^ layer_4[405]; 
    assign layer_5[393] = layer_4[402] & layer_4[402]; 
    assign layer_5[394] = ~(layer_4[407] | layer_4[393]); 
    assign layer_5[395] = layer_4[381] & layer_4[405]; 
    assign layer_5[396] = layer_4[398]; 
    assign layer_5[397] = layer_4[388] | layer_4[412]; 
    assign layer_5[398] = ~layer_4[405] | (layer_4[396] & layer_4[405]); 
    assign layer_5[399] = ~(layer_4[408] ^ layer_4[392]); 
    assign layer_5[400] = ~(layer_4[412] | layer_4[415]); 
    assign layer_5[401] = layer_4[412]; 
    assign layer_5[402] = ~(layer_4[392] ^ layer_4[413]); 
    assign layer_5[403] = ~(layer_4[414] ^ layer_4[416]); 
    assign layer_5[404] = ~layer_4[420]; 
    assign layer_5[405] = layer_4[415] & ~layer_4[410]; 
    assign layer_5[406] = ~layer_4[399] | (layer_4[399] & layer_4[420]); 
    assign layer_5[407] = layer_4[402] & ~layer_4[394]; 
    assign layer_5[408] = ~layer_4[392]; 
    assign layer_5[409] = ~layer_4[399] | (layer_4[399] & layer_4[410]); 
    assign layer_5[410] = ~(layer_4[416] ^ layer_4[409]); 
    assign layer_5[411] = ~(layer_4[408] ^ layer_4[402]); 
    assign layer_5[412] = layer_4[416] & ~layer_4[417]; 
    assign layer_5[413] = layer_4[429] | layer_4[410]; 
    assign layer_5[414] = layer_4[405] | layer_4[418]; 
    assign layer_5[415] = layer_4[420] ^ layer_4[426]; 
    assign layer_5[416] = ~(layer_4[416] & layer_4[411]); 
    assign layer_5[417] = layer_4[403]; 
    assign layer_5[418] = layer_4[427] ^ layer_4[403]; 
    assign layer_5[419] = layer_4[409] & layer_4[408]; 
    assign layer_5[420] = layer_4[411] ^ layer_4[429]; 
    assign layer_5[421] = layer_4[431] | layer_4[424]; 
    assign layer_5[422] = ~layer_4[422] | (layer_4[422] & layer_4[414]); 
    assign layer_5[423] = ~(layer_4[429] & layer_4[417]); 
    assign layer_5[424] = 1'b1; 
    assign layer_5[425] = layer_4[435] & layer_4[419]; 
    assign layer_5[426] = ~layer_4[418]; 
    assign layer_5[427] = 1'b1; 
    assign layer_5[428] = ~(layer_4[435] & layer_4[442]); 
    assign layer_5[429] = ~(layer_4[430] | layer_4[434]); 
    assign layer_5[430] = layer_4[422] & ~layer_4[420]; 
    assign layer_5[431] = ~(layer_4[447] ^ layer_4[425]); 
    assign layer_5[432] = ~layer_4[430] | (layer_4[447] & layer_4[430]); 
    assign layer_5[433] = 1'b0; 
    assign layer_5[434] = layer_4[434]; 
    assign layer_5[435] = ~layer_4[444]; 
    assign layer_5[436] = layer_4[429]; 
    assign layer_5[437] = 1'b1; 
    assign layer_5[438] = ~layer_4[439] | (layer_4[439] & layer_4[430]); 
    assign layer_5[439] = 1'b0; 
    assign layer_5[440] = 1'b0; 
    assign layer_5[441] = layer_4[454] & ~layer_4[440]; 
    assign layer_5[442] = ~layer_4[433]; 
    assign layer_5[443] = ~layer_4[427] | (layer_4[427] & layer_4[427]); 
    assign layer_5[444] = ~(layer_4[454] ^ layer_4[428]); 
    assign layer_5[445] = layer_4[436]; 
    assign layer_5[446] = ~layer_4[460]; 
    assign layer_5[447] = 1'b1; 
    assign layer_5[448] = ~(layer_4[459] ^ layer_4[450]); 
    assign layer_5[449] = ~(layer_4[439] | layer_4[441]); 
    assign layer_5[450] = layer_4[437] & ~layer_4[442]; 
    assign layer_5[451] = layer_4[457] & ~layer_4[463]; 
    assign layer_5[452] = ~layer_4[460]; 
    assign layer_5[453] = layer_4[453]; 
    assign layer_5[454] = layer_4[450]; 
    assign layer_5[455] = ~(layer_4[449] | layer_4[457]); 
    assign layer_5[456] = ~layer_4[448]; 
    assign layer_5[457] = layer_4[471] & layer_4[459]; 
    assign layer_5[458] = layer_4[456] | layer_4[446]; 
    assign layer_5[459] = 1'b1; 
    assign layer_5[460] = layer_4[463] & layer_4[471]; 
    assign layer_5[461] = ~layer_4[475] | (layer_4[475] & layer_4[470]); 
    assign layer_5[462] = ~(layer_4[478] ^ layer_4[455]); 
    assign layer_5[463] = layer_4[474]; 
    assign layer_5[464] = ~layer_4[450] | (layer_4[470] & layer_4[450]); 
    assign layer_5[465] = ~layer_4[453]; 
    assign layer_5[466] = layer_4[473] & layer_4[450]; 
    assign layer_5[467] = ~(layer_4[466] | layer_4[475]); 
    assign layer_5[468] = ~layer_4[481]; 
    assign layer_5[469] = ~layer_4[481] | (layer_4[462] & layer_4[481]); 
    assign layer_5[470] = layer_4[478] ^ layer_4[458]; 
    assign layer_5[471] = ~layer_4[457] | (layer_4[457] & layer_4[480]); 
    assign layer_5[472] = ~layer_4[459]; 
    assign layer_5[473] = ~(layer_4[484] & layer_4[480]); 
    assign layer_5[474] = layer_4[472] | layer_4[482]; 
    assign layer_5[475] = ~layer_4[462] | (layer_4[472] & layer_4[462]); 
    assign layer_5[476] = layer_4[479] | layer_4[491]; 
    assign layer_5[477] = ~layer_4[462]; 
    assign layer_5[478] = layer_4[472]; 
    assign layer_5[479] = ~(layer_4[494] | layer_4[486]); 
    assign layer_5[480] = ~layer_4[496] | (layer_4[496] & layer_4[480]); 
    assign layer_5[481] = ~(layer_4[497] | layer_4[490]); 
    assign layer_5[482] = layer_4[480] & layer_4[497]; 
    assign layer_5[483] = 1'b0; 
    assign layer_5[484] = layer_4[477] ^ layer_4[469]; 
    assign layer_5[485] = ~(layer_4[479] ^ layer_4[496]); 
    assign layer_5[486] = ~(layer_4[500] | layer_4[501]); 
    assign layer_5[487] = ~(layer_4[489] | layer_4[473]); 
    assign layer_5[488] = ~(layer_4[503] ^ layer_4[479]); 
    assign layer_5[489] = ~(layer_4[487] ^ layer_4[501]); 
    assign layer_5[490] = 1'b1; 
    assign layer_5[491] = 1'b1; 
    assign layer_5[492] = ~layer_4[490]; 
    assign layer_5[493] = layer_4[505]; 
    assign layer_5[494] = layer_4[490] & ~layer_4[500]; 
    assign layer_5[495] = layer_4[488] | layer_4[490]; 
    assign layer_5[496] = layer_4[512] | layer_4[496]; 
    assign layer_5[497] = layer_4[510] | layer_4[493]; 
    assign layer_5[498] = layer_4[483] ^ layer_4[482]; 
    assign layer_5[499] = ~layer_4[510]; 
    assign layer_5[500] = layer_4[508]; 
    assign layer_5[501] = layer_4[497] | layer_4[511]; 
    assign layer_5[502] = layer_4[505] & ~layer_4[515]; 
    assign layer_5[503] = layer_4[491] & ~layer_4[505]; 
    assign layer_5[504] = ~layer_4[514]; 
    assign layer_5[505] = layer_4[489] & ~layer_4[489]; 
    assign layer_5[506] = ~(layer_4[503] ^ layer_4[517]); 
    assign layer_5[507] = layer_4[513] & ~layer_4[505]; 
    assign layer_5[508] = layer_4[522] & ~layer_4[509]; 
    assign layer_5[509] = layer_4[496] & ~layer_4[524]; 
    assign layer_5[510] = ~(layer_4[514] | layer_4[508]); 
    assign layer_5[511] = layer_4[511] ^ layer_4[496]; 
    assign layer_5[512] = ~(layer_4[500] & layer_4[501]); 
    assign layer_5[513] = 1'b1; 
    assign layer_5[514] = ~layer_4[511]; 
    assign layer_5[515] = 1'b0; 
    assign layer_5[516] = 1'b1; 
    assign layer_5[517] = 1'b1; 
    assign layer_5[518] = ~layer_4[532]; 
    assign layer_5[519] = layer_4[524] & ~layer_4[523]; 
    assign layer_5[520] = layer_4[507] & ~layer_4[535]; 
    assign layer_5[521] = 1'b0; 
    assign layer_5[522] = layer_4[520] ^ layer_4[518]; 
    assign layer_5[523] = ~layer_4[526] | (layer_4[526] & layer_4[515]); 
    assign layer_5[524] = 1'b0; 
    assign layer_5[525] = layer_4[517] & ~layer_4[540]; 
    assign layer_5[526] = ~layer_4[533]; 
    assign layer_5[527] = ~(layer_4[531] & layer_4[526]); 
    assign layer_5[528] = layer_4[539] & layer_4[528]; 
    assign layer_5[529] = ~(layer_4[529] ^ layer_4[515]); 
    assign layer_5[530] = ~(layer_4[531] | layer_4[513]); 
    assign layer_5[531] = ~layer_4[544]; 
    assign layer_5[532] = layer_4[541] & ~layer_4[545]; 
    assign layer_5[533] = layer_4[526] & ~layer_4[522]; 
    assign layer_5[534] = layer_4[545] & ~layer_4[519]; 
    assign layer_5[535] = ~layer_4[549] | (layer_4[520] & layer_4[549]); 
    assign layer_5[536] = layer_4[538] & ~layer_4[547]; 
    assign layer_5[537] = 1'b1; 
    assign layer_5[538] = 1'b0; 
    assign layer_5[539] = layer_4[548] | layer_4[528]; 
    assign layer_5[540] = ~layer_4[526]; 
    assign layer_5[541] = layer_4[539] | layer_4[553]; 
    assign layer_5[542] = layer_4[547]; 
    assign layer_5[543] = layer_4[530] | layer_4[539]; 
    assign layer_5[544] = ~(layer_4[553] | layer_4[550]); 
    assign layer_5[545] = ~layer_4[533] | (layer_4[551] & layer_4[533]); 
    assign layer_5[546] = ~layer_4[531]; 
    assign layer_5[547] = ~layer_4[547]; 
    assign layer_5[548] = ~layer_4[555] | (layer_4[534] & layer_4[555]); 
    assign layer_5[549] = layer_4[552] & ~layer_4[558]; 
    assign layer_5[550] = ~(layer_4[536] ^ layer_4[547]); 
    assign layer_5[551] = layer_4[551] & layer_4[557]; 
    assign layer_5[552] = ~(layer_4[564] & layer_4[541]); 
    assign layer_5[553] = layer_4[541] & ~layer_4[565]; 
    assign layer_5[554] = layer_4[547] | layer_4[562]; 
    assign layer_5[555] = layer_4[550]; 
    assign layer_5[556] = ~layer_4[550]; 
    assign layer_5[557] = layer_4[552]; 
    assign layer_5[558] = ~layer_4[548] | (layer_4[570] & layer_4[548]); 
    assign layer_5[559] = layer_4[552] & ~layer_4[550]; 
    assign layer_5[560] = ~(layer_4[554] & layer_4[547]); 
    assign layer_5[561] = layer_4[567]; 
    assign layer_5[562] = layer_4[573]; 
    assign layer_5[563] = ~(layer_4[577] ^ layer_4[571]); 
    assign layer_5[564] = ~layer_4[567]; 
    assign layer_5[565] = layer_4[580] | layer_4[549]; 
    assign layer_5[566] = layer_4[574] & ~layer_4[567]; 
    assign layer_5[567] = ~(layer_4[561] | layer_4[571]); 
    assign layer_5[568] = ~(layer_4[572] ^ layer_4[564]); 
    assign layer_5[569] = ~layer_4[583]; 
    assign layer_5[570] = 1'b0; 
    assign layer_5[571] = layer_4[560] & layer_4[586]; 
    assign layer_5[572] = ~(layer_4[573] ^ layer_4[566]); 
    assign layer_5[573] = ~(layer_4[566] | layer_4[557]); 
    assign layer_5[574] = layer_4[584]; 
    assign layer_5[575] = layer_4[578]; 
    assign layer_5[576] = ~layer_4[581] | (layer_4[581] & layer_4[562]); 
    assign layer_5[577] = ~(layer_4[593] | layer_4[586]); 
    assign layer_5[578] = ~(layer_4[572] | layer_4[577]); 
    assign layer_5[579] = 1'b0; 
    assign layer_5[580] = ~(layer_4[588] | layer_4[566]); 
    assign layer_5[581] = ~(layer_4[589] & layer_4[582]); 
    assign layer_5[582] = 1'b1; 
    assign layer_5[583] = ~layer_4[598] | (layer_4[598] & layer_4[581]); 
    assign layer_5[584] = ~(layer_4[589] & layer_4[580]); 
    assign layer_5[585] = 1'b0; 
    assign layer_5[586] = ~layer_4[586]; 
    assign layer_5[587] = layer_4[590] & ~layer_4[600]; 
    assign layer_5[588] = layer_4[592]; 
    assign layer_5[589] = ~(layer_4[605] | layer_4[589]); 
    assign layer_5[590] = layer_4[585]; 
    assign layer_5[591] = ~layer_4[586] | (layer_4[586] & layer_4[600]); 
    assign layer_5[592] = ~layer_4[607]; 
    assign layer_5[593] = layer_4[581] & layer_4[604]; 
    assign layer_5[594] = 1'b1; 
    assign layer_5[595] = ~layer_4[585]; 
    assign layer_5[596] = ~(layer_4[587] ^ layer_4[609]); 
    assign layer_5[597] = layer_4[601] & layer_4[581]; 
    assign layer_5[598] = ~(layer_4[597] ^ layer_4[606]); 
    assign layer_5[599] = ~layer_4[613] | (layer_4[613] & layer_4[602]); 
    assign layer_5[600] = layer_4[586] ^ layer_4[611]; 
    assign layer_5[601] = layer_4[589]; 
    assign layer_5[602] = layer_4[616] | layer_4[587]; 
    assign layer_5[603] = 1'b1; 
    assign layer_5[604] = ~layer_4[608] | (layer_4[608] & layer_4[606]); 
    assign layer_5[605] = 1'b0; 
    assign layer_5[606] = layer_4[600] & layer_4[595]; 
    assign layer_5[607] = ~(layer_4[607] ^ layer_4[593]); 
    assign layer_5[608] = ~layer_4[593] | (layer_4[593] & layer_4[593]); 
    assign layer_5[609] = layer_4[607] ^ layer_4[610]; 
    assign layer_5[610] = layer_4[606] & ~layer_4[614]; 
    assign layer_5[611] = layer_4[616]; 
    assign layer_5[612] = layer_4[613]; 
    assign layer_5[613] = layer_4[619]; 
    assign layer_5[614] = layer_4[610]; 
    assign layer_5[615] = ~layer_4[630] | (layer_4[607] & layer_4[630]); 
    assign layer_5[616] = layer_4[599] & ~layer_4[605]; 
    assign layer_5[617] = ~(layer_4[615] ^ layer_4[609]); 
    assign layer_5[618] = 1'b1; 
    assign layer_5[619] = layer_4[630] & ~layer_4[627]; 
    assign layer_5[620] = ~(layer_4[635] | layer_4[620]); 
    assign layer_5[621] = layer_4[605]; 
    assign layer_5[622] = layer_4[630] | layer_4[623]; 
    assign layer_5[623] = layer_4[607] & layer_4[608]; 
    assign layer_5[624] = layer_4[631] | layer_4[634]; 
    assign layer_5[625] = ~(layer_4[614] ^ layer_4[635]); 
    assign layer_5[626] = layer_4[637] | layer_4[612]; 
    assign layer_5[627] = ~(layer_4[625] & layer_4[627]); 
    assign layer_5[628] = ~(layer_4[621] ^ layer_4[625]); 
    assign layer_5[629] = layer_4[639] ^ layer_4[622]; 
    assign layer_5[630] = layer_4[631] & ~layer_4[618]; 
    assign layer_5[631] = ~(layer_4[627] & layer_4[623]); 
    assign layer_5[632] = 1'b1; 
    assign layer_5[633] = ~layer_4[642] | (layer_4[640] & layer_4[642]); 
    assign layer_5[634] = layer_4[647] & ~layer_4[625]; 
    assign layer_5[635] = ~layer_4[625]; 
    assign layer_5[636] = 1'b1; 
    assign layer_5[637] = layer_4[649] | layer_4[648]; 
    assign layer_5[638] = ~layer_4[644] | (layer_4[641] & layer_4[644]); 
    assign layer_5[639] = ~(layer_4[624] & layer_4[629]); 
    assign layer_5[640] = layer_4[652] & ~layer_4[655]; 
    assign layer_5[641] = ~(layer_4[632] & layer_4[656]); 
    assign layer_5[642] = layer_4[634] & ~layer_4[635]; 
    assign layer_5[643] = layer_4[653] & ~layer_4[631]; 
    assign layer_5[644] = layer_4[643] | layer_4[650]; 
    assign layer_5[645] = layer_4[653] & ~layer_4[659]; 
    assign layer_5[646] = layer_4[634] & ~layer_4[638]; 
    assign layer_5[647] = ~(layer_4[647] | layer_4[655]); 
    assign layer_5[648] = ~layer_4[636] | (layer_4[661] & layer_4[636]); 
    assign layer_5[649] = layer_4[661] & ~layer_4[636]; 
    assign layer_5[650] = layer_4[645]; 
    assign layer_5[651] = layer_4[643] | layer_4[638]; 
    assign layer_5[652] = ~layer_4[651] | (layer_4[651] & layer_4[636]); 
    assign layer_5[653] = layer_4[656] | layer_4[639]; 
    assign layer_5[654] = 1'b1; 
    assign layer_5[655] = 1'b0; 
    assign layer_5[656] = ~(layer_4[663] | layer_4[654]); 
    assign layer_5[657] = ~(layer_4[667] | layer_4[670]); 
    assign layer_5[658] = layer_4[647]; 
    assign layer_5[659] = layer_4[655] & ~layer_4[650]; 
    assign layer_5[660] = ~layer_4[662]; 
    assign layer_5[661] = ~(layer_4[652] ^ layer_4[649]); 
    assign layer_5[662] = layer_4[663] ^ layer_4[647]; 
    assign layer_5[663] = ~(layer_4[651] & layer_4[666]); 
    assign layer_5[664] = layer_4[657] & ~layer_4[661]; 
    assign layer_5[665] = ~(layer_4[665] & layer_4[674]); 
    assign layer_5[666] = layer_4[671]; 
    assign layer_5[667] = layer_4[680]; 
    assign layer_5[668] = layer_4[681] ^ layer_4[671]; 
    assign layer_5[669] = layer_4[657] & layer_4[665]; 
    assign layer_5[670] = layer_4[682] & ~layer_4[683]; 
    assign layer_5[671] = ~layer_4[662] | (layer_4[662] & layer_4[671]); 
    assign layer_5[672] = layer_4[668] & layer_4[687]; 
    assign layer_5[673] = ~layer_4[662]; 
    assign layer_5[674] = layer_4[673] ^ layer_4[663]; 
    assign layer_5[675] = ~(layer_4[670] ^ layer_4[684]); 
    assign layer_5[676] = layer_4[686] & ~layer_4[667]; 
    assign layer_5[677] = ~layer_4[666] | (layer_4[682] & layer_4[666]); 
    assign layer_5[678] = ~(layer_4[682] & layer_4[674]); 
    assign layer_5[679] = ~layer_4[667] | (layer_4[679] & layer_4[667]); 
    assign layer_5[680] = ~layer_4[686] | (layer_4[686] & layer_4[673]); 
    assign layer_5[681] = ~layer_4[685]; 
    assign layer_5[682] = ~layer_4[681]; 
    assign layer_5[683] = layer_4[677] | layer_4[673]; 
    assign layer_5[684] = ~layer_4[688]; 
    assign layer_5[685] = ~(layer_4[676] | layer_4[682]); 
    assign layer_5[686] = ~layer_4[696]; 
    assign layer_5[687] = layer_4[694] ^ layer_4[688]; 
    assign layer_5[688] = 1'b1; 
    assign layer_5[689] = layer_4[674] ^ layer_4[672]; 
    assign layer_5[690] = layer_4[691] & ~layer_4[686]; 
    assign layer_5[691] = layer_4[689] & ~layer_4[689]; 
    assign layer_5[692] = ~layer_4[698]; 
    assign layer_5[693] = 1'b1; 
    assign layer_5[694] = ~(layer_4[704] & layer_4[681]); 
    assign layer_5[695] = layer_4[680] & layer_4[689]; 
    assign layer_5[696] = ~(layer_4[695] ^ layer_4[688]); 
    assign layer_5[697] = 1'b0; 
    assign layer_5[698] = ~layer_4[692]; 
    assign layer_5[699] = layer_4[711]; 
    assign layer_5[700] = ~(layer_4[700] & layer_4[696]); 
    assign layer_5[701] = ~layer_4[707]; 
    assign layer_5[702] = ~layer_4[717]; 
    assign layer_5[703] = ~(layer_4[700] & layer_4[697]); 
    assign layer_5[704] = ~layer_4[719]; 
    assign layer_5[705] = ~(layer_4[714] & layer_4[708]); 
    assign layer_5[706] = 1'b0; 
    assign layer_5[707] = layer_4[699] ^ layer_4[695]; 
    assign layer_5[708] = ~layer_4[699]; 
    assign layer_5[709] = ~(layer_4[695] ^ layer_4[704]); 
    assign layer_5[710] = layer_4[724]; 
    assign layer_5[711] = ~(layer_4[698] ^ layer_4[697]); 
    assign layer_5[712] = layer_4[723] & layer_4[719]; 
    assign layer_5[713] = layer_4[698] & ~layer_4[699]; 
    assign layer_5[714] = ~(layer_4[712] | layer_4[717]); 
    assign layer_5[715] = 1'b1; 
    assign layer_5[716] = ~layer_4[703] | (layer_4[717] & layer_4[703]); 
    assign layer_5[717] = layer_4[717] | layer_4[717]; 
    assign layer_5[718] = ~layer_4[728]; 
    assign layer_5[719] = ~layer_4[708]; 
    assign layer_5[720] = ~(layer_4[713] ^ layer_4[727]); 
    assign layer_5[721] = 1'b0; 
    assign layer_5[722] = layer_4[709] ^ layer_4[707]; 
    assign layer_5[723] = layer_4[729]; 
    assign layer_5[724] = layer_4[727] & layer_4[737]; 
    assign layer_5[725] = ~layer_4[737] | (layer_4[737] & layer_4[735]); 
    assign layer_5[726] = 1'b0; 
    assign layer_5[727] = layer_4[715] & ~layer_4[731]; 
    assign layer_5[728] = layer_4[724] ^ layer_4[742]; 
    assign layer_5[729] = layer_4[735]; 
    assign layer_5[730] = 1'b1; 
    assign layer_5[731] = layer_4[722] & ~layer_4[720]; 
    assign layer_5[732] = layer_4[736] | layer_4[733]; 
    assign layer_5[733] = ~(layer_4[742] ^ layer_4[718]); 
    assign layer_5[734] = layer_4[739] ^ layer_4[727]; 
    assign layer_5[735] = layer_4[736] ^ layer_4[746]; 
    assign layer_5[736] = layer_4[730] ^ layer_4[751]; 
    assign layer_5[737] = 1'b0; 
    assign layer_5[738] = ~layer_4[734] | (layer_4[734] & layer_4[728]); 
    assign layer_5[739] = ~layer_4[730] | (layer_4[747] & layer_4[730]); 
    assign layer_5[740] = layer_4[732] | layer_4[748]; 
    assign layer_5[741] = layer_4[755] & ~layer_4[745]; 
    assign layer_5[742] = 1'b0; 
    assign layer_5[743] = layer_4[735] & ~layer_4[730]; 
    assign layer_5[744] = ~(layer_4[736] | layer_4[734]); 
    assign layer_5[745] = ~layer_4[735] | (layer_4[735] & layer_4[735]); 
    assign layer_5[746] = layer_4[745] ^ layer_4[738]; 
    assign layer_5[747] = ~layer_4[740] | (layer_4[740] & layer_4[745]); 
    assign layer_5[748] = ~(layer_4[736] & layer_4[737]); 
    assign layer_5[749] = ~(layer_4[761] ^ layer_4[763]); 
    assign layer_5[750] = layer_4[740] & ~layer_4[743]; 
    assign layer_5[751] = layer_4[735]; 
    assign layer_5[752] = layer_4[746] & ~layer_4[745]; 
    assign layer_5[753] = layer_4[739] & layer_4[744]; 
    assign layer_5[754] = layer_4[750] | layer_4[738]; 
    assign layer_5[755] = layer_4[742] ^ layer_4[760]; 
    assign layer_5[756] = ~layer_4[749] | (layer_4[769] & layer_4[749]); 
    assign layer_5[757] = layer_4[771] | layer_4[746]; 
    assign layer_5[758] = ~layer_4[763] | (layer_4[763] & layer_4[769]); 
    assign layer_5[759] = ~(layer_4[746] | layer_4[773]); 
    assign layer_5[760] = layer_4[746]; 
    assign layer_5[761] = layer_4[757] & layer_4[760]; 
    assign layer_5[762] = ~(layer_4[772] ^ layer_4[769]); 
    assign layer_5[763] = layer_4[761] & ~layer_4[762]; 
    assign layer_5[764] = ~layer_4[751] | (layer_4[762] & layer_4[751]); 
    assign layer_5[765] = ~layer_4[771]; 
    assign layer_5[766] = layer_4[776]; 
    assign layer_5[767] = 1'b0; 
    assign layer_5[768] = ~layer_4[756]; 
    assign layer_5[769] = layer_4[756]; 
    assign layer_5[770] = ~layer_4[784]; 
    assign layer_5[771] = ~layer_4[775]; 
    assign layer_5[772] = ~(layer_4[776] | layer_4[774]); 
    assign layer_5[773] = layer_4[767] & layer_4[771]; 
    assign layer_5[774] = 1'b1; 
    assign layer_5[775] = ~layer_4[759] | (layer_4[782] & layer_4[759]); 
    assign layer_5[776] = layer_4[778] & layer_4[769]; 
    assign layer_5[777] = layer_4[763] ^ layer_4[784]; 
    assign layer_5[778] = ~(layer_4[787] & layer_4[773]); 
    assign layer_5[779] = layer_4[787]; 
    assign layer_5[780] = layer_4[790]; 
    assign layer_5[781] = layer_4[787] & ~layer_4[793]; 
    assign layer_5[782] = ~(layer_4[780] ^ layer_4[779]); 
    assign layer_5[783] = layer_4[769] & ~layer_4[776]; 
    assign layer_5[784] = ~layer_4[783]; 
    assign layer_5[785] = 1'b0; 
    assign layer_5[786] = ~layer_4[771] | (layer_4[771] & layer_4[777]); 
    assign layer_5[787] = layer_4[780] & ~layer_4[801]; 
    assign layer_5[788] = 1'b1; 
    assign layer_5[789] = ~layer_4[800] | (layer_4[803] & layer_4[800]); 
    assign layer_5[790] = 1'b0; 
    assign layer_5[791] = ~(layer_4[807] | layer_4[795]); 
    assign layer_5[792] = layer_4[790] ^ layer_4[781]; 
    assign layer_5[793] = 1'b1; 
    assign layer_5[794] = layer_4[801] & ~layer_4[805]; 
    assign layer_5[795] = layer_4[793] & ~layer_4[780]; 
    assign layer_5[796] = layer_4[796]; 
    assign layer_5[797] = ~(layer_4[786] | layer_4[797]); 
    assign layer_5[798] = 1'b0; 
    assign layer_5[799] = ~(layer_4[788] & layer_4[789]); 
    assign layer_5[800] = layer_4[783]; 
    assign layer_5[801] = 1'b1; 
    assign layer_5[802] = ~layer_4[790]; 
    assign layer_5[803] = layer_4[802] & layer_4[806]; 
    assign layer_5[804] = 1'b0; 
    assign layer_5[805] = 1'b1; 
    assign layer_5[806] = ~layer_4[815] | (layer_4[812] & layer_4[815]); 
    assign layer_5[807] = ~layer_4[799]; 
    assign layer_5[808] = ~(layer_4[796] ^ layer_4[811]); 
    assign layer_5[809] = layer_4[799] ^ layer_4[806]; 
    assign layer_5[810] = ~(layer_4[813] & layer_4[794]); 
    assign layer_5[811] = ~layer_4[805] | (layer_4[805] & layer_4[813]); 
    assign layer_5[812] = ~layer_4[827]; 
    assign layer_5[813] = ~(layer_4[804] | layer_4[811]); 
    assign layer_5[814] = ~layer_4[801] | (layer_4[801] & layer_4[800]); 
    assign layer_5[815] = ~(layer_4[815] & layer_4[812]); 
    assign layer_5[816] = 1'b1; 
    assign layer_5[817] = ~layer_4[813]; 
    assign layer_5[818] = ~(layer_4[812] | layer_4[823]); 
    assign layer_5[819] = layer_4[823] & layer_4[810]; 
    assign layer_5[820] = layer_4[828] | layer_4[820]; 
    assign layer_5[821] = layer_4[816] & ~layer_4[818]; 
    assign layer_5[822] = layer_4[807] & ~layer_4[807]; 
    assign layer_5[823] = layer_4[825] & layer_4[825]; 
    assign layer_5[824] = layer_4[810] & ~layer_4[840]; 
    assign layer_5[825] = ~(layer_4[812] | layer_4[826]); 
    assign layer_5[826] = ~layer_4[835]; 
    assign layer_5[827] = layer_4[829] ^ layer_4[840]; 
    assign layer_5[828] = layer_4[838]; 
    assign layer_5[829] = layer_4[813] & ~layer_4[829]; 
    assign layer_5[830] = ~layer_4[820] | (layer_4[820] & layer_4[813]); 
    assign layer_5[831] = layer_4[822] & layer_4[836]; 
    assign layer_5[832] = layer_4[834] ^ layer_4[821]; 
    assign layer_5[833] = 1'b0; 
    assign layer_5[834] = layer_4[837] & ~layer_4[829]; 
    assign layer_5[835] = layer_4[851] | layer_4[844]; 
    assign layer_5[836] = ~(layer_4[850] & layer_4[849]); 
    assign layer_5[837] = 1'b1; 
    assign layer_5[838] = layer_4[834]; 
    assign layer_5[839] = ~layer_4[835]; 
    assign layer_5[840] = ~(layer_4[841] ^ layer_4[826]); 
    assign layer_5[841] = ~layer_4[835]; 
    assign layer_5[842] = ~layer_4[840] | (layer_4[840] & layer_4[834]); 
    assign layer_5[843] = ~layer_4[844]; 
    assign layer_5[844] = layer_4[837] ^ layer_4[850]; 
    assign layer_5[845] = ~layer_4[849] | (layer_4[858] & layer_4[849]); 
    assign layer_5[846] = layer_4[833] & ~layer_4[847]; 
    assign layer_5[847] = layer_4[859] | layer_4[852]; 
    assign layer_5[848] = layer_4[863] | layer_4[833]; 
    assign layer_5[849] = ~(layer_4[838] ^ layer_4[862]); 
    assign layer_5[850] = ~(layer_4[860] ^ layer_4[848]); 
    assign layer_5[851] = layer_4[860] | layer_4[861]; 
    assign layer_5[852] = layer_4[840] ^ layer_4[837]; 
    assign layer_5[853] = layer_4[848] & ~layer_4[845]; 
    assign layer_5[854] = layer_4[867]; 
    assign layer_5[855] = ~layer_4[852] | (layer_4[852] & layer_4[862]); 
    assign layer_5[856] = layer_4[867] & layer_4[871]; 
    assign layer_5[857] = ~layer_4[863]; 
    assign layer_5[858] = ~(layer_4[860] | layer_4[873]); 
    assign layer_5[859] = 1'b1; 
    assign layer_5[860] = layer_4[868] & layer_4[858]; 
    assign layer_5[861] = layer_4[855] & ~layer_4[876]; 
    assign layer_5[862] = ~(layer_4[867] ^ layer_4[855]); 
    assign layer_5[863] = 1'b0; 
    assign layer_5[864] = ~layer_4[853]; 
    assign layer_5[865] = layer_4[852] & layer_4[861]; 
    assign layer_5[866] = ~layer_4[874]; 
    assign layer_5[867] = 1'b0; 
    assign layer_5[868] = layer_4[873]; 
    assign layer_5[869] = layer_4[882] & ~layer_4[877]; 
    assign layer_5[870] = layer_4[878] & ~layer_4[878]; 
    assign layer_5[871] = ~layer_4[869] | (layer_4[866] & layer_4[869]); 
    assign layer_5[872] = layer_4[872] & ~layer_4[864]; 
    assign layer_5[873] = ~(layer_4[879] ^ layer_4[858]); 
    assign layer_5[874] = ~layer_4[878]; 
    assign layer_5[875] = 1'b0; 
    assign layer_5[876] = layer_4[887] & ~layer_4[873]; 
    assign layer_5[877] = 1'b1; 
    assign layer_5[878] = ~(layer_4[886] & layer_4[887]); 
    assign layer_5[879] = ~layer_4[862]; 
    assign layer_5[880] = layer_4[868]; 
    assign layer_5[881] = ~(layer_4[884] | layer_4[871]); 
    assign layer_5[882] = layer_4[883] | layer_4[871]; 
    assign layer_5[883] = layer_4[896] | layer_4[870]; 
    assign layer_5[884] = ~layer_4[887] | (layer_4[881] & layer_4[887]); 
    assign layer_5[885] = layer_4[891] & ~layer_4[871]; 
    assign layer_5[886] = layer_4[888] | layer_4[896]; 
    assign layer_5[887] = layer_4[899] & layer_4[884]; 
    assign layer_5[888] = ~layer_4[879] | (layer_4[879] & layer_4[872]); 
    assign layer_5[889] = 1'b1; 
    assign layer_5[890] = ~(layer_4[876] ^ layer_4[892]); 
    assign layer_5[891] = layer_4[898] & layer_4[897]; 
    assign layer_5[892] = ~layer_4[881] | (layer_4[908] & layer_4[881]); 
    assign layer_5[893] = layer_4[887] & layer_4[876]; 
    assign layer_5[894] = ~layer_4[883] | (layer_4[892] & layer_4[883]); 
    assign layer_5[895] = ~layer_4[905] | (layer_4[905] & layer_4[905]); 
    assign layer_5[896] = layer_4[897]; 
    assign layer_5[897] = ~layer_4[893] | (layer_4[893] & layer_4[911]); 
    assign layer_5[898] = layer_4[886] | layer_4[885]; 
    assign layer_5[899] = layer_4[894]; 
    assign layer_5[900] = ~layer_4[891] | (layer_4[891] & layer_4[893]); 
    assign layer_5[901] = ~layer_4[899] | (layer_4[904] & layer_4[899]); 
    assign layer_5[902] = ~layer_4[891]; 
    assign layer_5[903] = layer_4[907] | layer_4[886]; 
    assign layer_5[904] = 1'b0; 
    assign layer_5[905] = layer_4[899]; 
    assign layer_5[906] = ~layer_4[898] | (layer_4[898] & layer_4[892]); 
    assign layer_5[907] = ~layer_4[911] | (layer_4[895] & layer_4[911]); 
    assign layer_5[908] = layer_4[901] | layer_4[904]; 
    assign layer_5[909] = ~(layer_4[893] | layer_4[909]); 
    assign layer_5[910] = layer_4[906]; 
    assign layer_5[911] = layer_4[917]; 
    assign layer_5[912] = ~(layer_4[920] | layer_4[900]); 
    assign layer_5[913] = 1'b1; 
    assign layer_5[914] = ~(layer_4[909] & layer_4[903]); 
    assign layer_5[915] = ~layer_4[924] | (layer_4[915] & layer_4[924]); 
    assign layer_5[916] = 1'b0; 
    assign layer_5[917] = layer_4[928] & ~layer_4[930]; 
    assign layer_5[918] = layer_4[932] & ~layer_4[907]; 
    assign layer_5[919] = layer_4[912] & ~layer_4[914]; 
    assign layer_5[920] = ~(layer_4[914] | layer_4[933]); 
    assign layer_5[921] = layer_4[934] ^ layer_4[930]; 
    assign layer_5[922] = layer_4[926] ^ layer_4[919]; 
    assign layer_5[923] = ~(layer_4[915] ^ layer_4[922]); 
    assign layer_5[924] = ~(layer_4[919] | layer_4[936]); 
    assign layer_5[925] = layer_4[935] | layer_4[909]; 
    assign layer_5[926] = ~layer_4[942] | (layer_4[942] & layer_4[923]); 
    assign layer_5[927] = ~layer_4[926] | (layer_4[926] & layer_4[910]); 
    assign layer_5[928] = ~layer_4[943] | (layer_4[943] & layer_4[922]); 
    assign layer_5[929] = layer_4[937] & ~layer_4[931]; 
    assign layer_5[930] = ~layer_4[918] | (layer_4[921] & layer_4[918]); 
    assign layer_5[931] = layer_4[920] & ~layer_4[937]; 
    assign layer_5[932] = layer_4[926] ^ layer_4[926]; 
    assign layer_5[933] = layer_4[941] & ~layer_4[948]; 
    assign layer_5[934] = ~(layer_4[948] ^ layer_4[947]); 
    assign layer_5[935] = ~layer_4[945]; 
    assign layer_5[936] = layer_4[943]; 
    assign layer_5[937] = layer_4[940]; 
    assign layer_5[938] = ~layer_4[929] | (layer_4[953] & layer_4[929]); 
    assign layer_5[939] = ~layer_4[924] | (layer_4[924] & layer_4[950]); 
    assign layer_5[940] = layer_4[952]; 
    assign layer_5[941] = layer_4[953] ^ layer_4[953]; 
    assign layer_5[942] = ~layer_4[936]; 
    assign layer_5[943] = ~layer_4[935] | (layer_4[935] & layer_4[956]); 
    assign layer_5[944] = ~layer_4[956]; 
    assign layer_5[945] = 1'b1; 
    assign layer_5[946] = ~(layer_4[943] | layer_4[940]); 
    assign layer_5[947] = layer_4[935] & layer_4[932]; 
    assign layer_5[948] = ~(layer_4[957] | layer_4[948]); 
    assign layer_5[949] = layer_4[938]; 
    assign layer_5[950] = ~(layer_4[955] ^ layer_4[945]); 
    assign layer_5[951] = ~(layer_4[954] | layer_4[959]); 
    assign layer_5[952] = layer_4[938] & layer_4[935]; 
    assign layer_5[953] = ~(layer_4[958] & layer_4[959]); 
    assign layer_5[954] = layer_4[946] & layer_4[941]; 
    assign layer_5[955] = 1'b1; 
    assign layer_5[956] = ~(layer_4[949] | layer_4[947]); 
    assign layer_5[957] = ~layer_4[965]; 
    assign layer_5[958] = layer_4[945]; 
    assign layer_5[959] = layer_4[958]; 
    assign layer_5[960] = layer_4[951] & ~layer_4[971]; 
    assign layer_5[961] = layer_4[968] ^ layer_4[955]; 
    assign layer_5[962] = ~layer_4[978]; 
    assign layer_5[963] = 1'b1; 
    assign layer_5[964] = layer_4[951] & ~layer_4[954]; 
    assign layer_5[965] = layer_4[954] & ~layer_4[981]; 
    assign layer_5[966] = layer_4[972] & ~layer_4[954]; 
    assign layer_5[967] = layer_4[955]; 
    assign layer_5[968] = layer_4[965] | layer_4[974]; 
    assign layer_5[969] = 1'b0; 
    assign layer_5[970] = layer_4[965] & ~layer_4[959]; 
    assign layer_5[971] = ~layer_4[986]; 
    assign layer_5[972] = ~layer_4[974]; 
    assign layer_5[973] = layer_4[968] | layer_4[956]; 
    assign layer_5[974] = 1'b1; 
    assign layer_5[975] = layer_4[968] | layer_4[976]; 
    assign layer_5[976] = ~layer_4[967] | (layer_4[967] & layer_4[965]); 
    assign layer_5[977] = layer_4[969]; 
    assign layer_5[978] = layer_4[966]; 
    assign layer_5[979] = ~layer_4[983] | (layer_4[964] & layer_4[983]); 
    assign layer_5[980] = layer_4[987] | layer_4[981]; 
    assign layer_5[981] = layer_4[967]; 
    assign layer_5[982] = ~(layer_4[984] & layer_4[968]); 
    assign layer_5[983] = ~(layer_4[978] & layer_4[988]); 
    assign layer_5[984] = ~layer_4[989] | (layer_4[989] & layer_4[972]); 
    assign layer_5[985] = layer_4[969]; 
    assign layer_5[986] = ~(layer_4[998] ^ layer_4[978]); 
    assign layer_5[987] = 1'b1; 
    assign layer_5[988] = layer_4[1002] & ~layer_4[986]; 
    assign layer_5[989] = layer_4[982]; 
    assign layer_5[990] = layer_4[974]; 
    assign layer_5[991] = layer_4[998] | layer_4[995]; 
    assign layer_5[992] = layer_4[977] ^ layer_4[990]; 
    assign layer_5[993] = layer_4[999]; 
    assign layer_5[994] = ~layer_4[1003] | (layer_4[1003] & layer_4[987]); 
    assign layer_5[995] = ~(layer_4[990] | layer_4[1005]); 
    assign layer_5[996] = ~(layer_4[1008] | layer_4[1004]); 
    assign layer_5[997] = ~(layer_4[995] ^ layer_4[1005]); 
    assign layer_5[998] = ~(layer_4[1011] ^ layer_4[985]); 
    assign layer_5[999] = layer_4[1008] | layer_4[990]; 
    assign layer_5[1000] = layer_4[1012] & ~layer_4[996]; 
    assign layer_5[1001] = layer_4[999] & ~layer_4[1017]; 
    assign layer_5[1002] = ~(layer_4[996] | layer_4[1016]); 
    assign layer_5[1003] = ~layer_4[999] | (layer_4[999] & layer_4[999]); 
    assign layer_5[1004] = layer_4[1013] ^ layer_4[987]; 
    assign layer_5[1005] = layer_4[1001] & ~layer_4[1016]; 
    assign layer_5[1006] = ~(layer_4[995] | layer_4[1017]); 
    assign layer_5[1007] = ~layer_4[1004]; 
    assign layer_5[1008] = ~(layer_4[994] ^ layer_4[1006]); 
    assign layer_5[1009] = layer_4[1007] & layer_4[997]; 
    assign layer_5[1010] = ~(layer_4[1023] ^ layer_4[1004]); 
    assign layer_5[1011] = layer_4[1008] & ~layer_4[1014]; 
    assign layer_5[1012] = ~layer_4[996]; 
    assign layer_5[1013] = ~layer_4[1018]; 
    assign layer_5[1014] = ~(layer_4[1022] & layer_4[998]); 
    assign layer_5[1015] = layer_4[1017]; 
    assign layer_5[1016] = layer_4[1016]; 
    assign layer_5[1017] = layer_4[1019] & ~layer_4[1001]; 
    assign layer_5[1018] = layer_4[1023] & ~layer_4[1021]; 
    assign layer_5[1019] = layer_4[1022] & ~layer_4[1021]; 
    assign layer_5[1020] = layer_4[1020] & layer_4[1009]; 
    assign layer_5[1021] = ~layer_4[1020]; 
    assign layer_5[1022] = ~layer_4[1011] | (layer_4[1009] & layer_4[1011]); 
    assign layer_5[1023] = 1'b0; 
    // Layer 6 ============================================================
    assign layer_6[0] = 1'b1; 
    assign layer_6[1] = ~(layer_5[5] ^ layer_5[16]); 
    assign layer_6[2] = ~layer_5[4]; 
    assign layer_6[3] = layer_5[3] ^ layer_5[18]; 
    assign layer_6[4] = layer_5[10]; 
    assign layer_6[5] = layer_5[11]; 
    assign layer_6[6] = layer_5[4] & ~layer_5[9]; 
    assign layer_6[7] = layer_5[11] ^ layer_5[12]; 
    assign layer_6[8] = ~layer_5[11]; 
    assign layer_6[9] = 1'b1; 
    assign layer_6[10] = ~(layer_5[10] ^ layer_5[10]); 
    assign layer_6[11] = layer_5[19] & ~layer_5[8]; 
    assign layer_6[12] = ~(layer_5[22] | layer_5[0]); 
    assign layer_6[13] = layer_5[28] & ~layer_5[12]; 
    assign layer_6[14] = ~(layer_5[1] ^ layer_5[5]); 
    assign layer_6[15] = layer_5[19] & layer_5[21]; 
    assign layer_6[16] = 1'b1; 
    assign layer_6[17] = ~(layer_5[29] ^ layer_5[3]); 
    assign layer_6[18] = 1'b0; 
    assign layer_6[19] = ~layer_5[26] | (layer_5[26] & layer_5[11]); 
    assign layer_6[20] = layer_5[19]; 
    assign layer_6[21] = ~(layer_5[27] | layer_5[15]); 
    assign layer_6[22] = 1'b1; 
    assign layer_6[23] = 1'b0; 
    assign layer_6[24] = ~(layer_5[36] | layer_5[37]); 
    assign layer_6[25] = 1'b1; 
    assign layer_6[26] = ~(layer_5[34] | layer_5[9]); 
    assign layer_6[27] = layer_5[19] & ~layer_5[38]; 
    assign layer_6[28] = layer_5[13]; 
    assign layer_6[29] = layer_5[44] & ~layer_5[29]; 
    assign layer_6[30] = ~layer_5[41] | (layer_5[31] & layer_5[41]); 
    assign layer_6[31] = ~layer_5[37]; 
    assign layer_6[32] = layer_5[23] & ~layer_5[43]; 
    assign layer_6[33] = layer_5[27]; 
    assign layer_6[34] = ~layer_5[34]; 
    assign layer_6[35] = ~(layer_5[49] | layer_5[20]); 
    assign layer_6[36] = ~layer_5[42] | (layer_5[44] & layer_5[42]); 
    assign layer_6[37] = ~layer_5[42]; 
    assign layer_6[38] = ~layer_5[31]; 
    assign layer_6[39] = layer_5[44]; 
    assign layer_6[40] = ~(layer_5[56] & layer_5[32]); 
    assign layer_6[41] = ~layer_5[41] | (layer_5[51] & layer_5[41]); 
    assign layer_6[42] = ~layer_5[43]; 
    assign layer_6[43] = 1'b0; 
    assign layer_6[44] = layer_5[47] | layer_5[45]; 
    assign layer_6[45] = ~(layer_5[35] & layer_5[58]); 
    assign layer_6[46] = layer_5[49]; 
    assign layer_6[47] = layer_5[52] & ~layer_5[54]; 
    assign layer_6[48] = layer_5[59] & layer_5[31]; 
    assign layer_6[49] = layer_5[53] & layer_5[50]; 
    assign layer_6[50] = layer_5[40] ^ layer_5[51]; 
    assign layer_6[51] = ~(layer_5[56] ^ layer_5[34]); 
    assign layer_6[52] = 1'b1; 
    assign layer_6[53] = layer_5[53]; 
    assign layer_6[54] = layer_5[50]; 
    assign layer_6[55] = layer_5[69]; 
    assign layer_6[56] = ~layer_5[54]; 
    assign layer_6[57] = ~layer_5[72] | (layer_5[73] & layer_5[72]); 
    assign layer_6[58] = 1'b0; 
    assign layer_6[59] = ~layer_5[73]; 
    assign layer_6[60] = layer_5[47] & layer_5[70]; 
    assign layer_6[61] = layer_5[51] | layer_5[45]; 
    assign layer_6[62] = ~(layer_5[70] | layer_5[45]); 
    assign layer_6[63] = ~layer_5[74]; 
    assign layer_6[64] = ~layer_5[73] | (layer_5[62] & layer_5[73]); 
    assign layer_6[65] = layer_5[57] | layer_5[72]; 
    assign layer_6[66] = layer_5[57]; 
    assign layer_6[67] = ~layer_5[72]; 
    assign layer_6[68] = 1'b1; 
    assign layer_6[69] = layer_5[56] | layer_5[74]; 
    assign layer_6[70] = layer_5[61] & layer_5[58]; 
    assign layer_6[71] = layer_5[73] ^ layer_5[77]; 
    assign layer_6[72] = layer_5[84] | layer_5[77]; 
    assign layer_6[73] = layer_5[62] & ~layer_5[73]; 
    assign layer_6[74] = ~layer_5[76] | (layer_5[76] & layer_5[65]); 
    assign layer_6[75] = layer_5[84] & ~layer_5[74]; 
    assign layer_6[76] = ~layer_5[60]; 
    assign layer_6[77] = layer_5[79] ^ layer_5[77]; 
    assign layer_6[78] = layer_5[77] & layer_5[69]; 
    assign layer_6[79] = ~layer_5[67] | (layer_5[86] & layer_5[67]); 
    assign layer_6[80] = ~(layer_5[82] & layer_5[89]); 
    assign layer_6[81] = ~layer_5[77]; 
    assign layer_6[82] = layer_5[88] & ~layer_5[97]; 
    assign layer_6[83] = layer_5[89] & layer_5[69]; 
    assign layer_6[84] = layer_5[86] & layer_5[68]; 
    assign layer_6[85] = layer_5[91]; 
    assign layer_6[86] = ~layer_5[85] | (layer_5[85] & layer_5[76]); 
    assign layer_6[87] = ~layer_5[79] | (layer_5[91] & layer_5[79]); 
    assign layer_6[88] = ~(layer_5[87] | layer_5[98]); 
    assign layer_6[89] = layer_5[76] | layer_5[81]; 
    assign layer_6[90] = ~layer_5[88]; 
    assign layer_6[91] = 1'b1; 
    assign layer_6[92] = 1'b0; 
    assign layer_6[93] = 1'b0; 
    assign layer_6[94] = layer_5[107]; 
    assign layer_6[95] = layer_5[91] | layer_5[103]; 
    assign layer_6[96] = ~(layer_5[104] | layer_5[104]); 
    assign layer_6[97] = ~layer_5[98] | (layer_5[98] & layer_5[81]); 
    assign layer_6[98] = layer_5[84]; 
    assign layer_6[99] = layer_5[90]; 
    assign layer_6[100] = 1'b0; 
    assign layer_6[101] = layer_5[107]; 
    assign layer_6[102] = ~layer_5[89] | (layer_5[96] & layer_5[89]); 
    assign layer_6[103] = ~layer_5[94]; 
    assign layer_6[104] = layer_5[109] & layer_5[106]; 
    assign layer_6[105] = ~layer_5[113] | (layer_5[113] & layer_5[101]); 
    assign layer_6[106] = layer_5[103] & layer_5[108]; 
    assign layer_6[107] = ~(layer_5[95] | layer_5[101]); 
    assign layer_6[108] = ~(layer_5[104] ^ layer_5[111]); 
    assign layer_6[109] = layer_5[113] & layer_5[118]; 
    assign layer_6[110] = layer_5[114] ^ layer_5[106]; 
    assign layer_6[111] = layer_5[127]; 
    assign layer_6[112] = ~(layer_5[111] | layer_5[123]); 
    assign layer_6[113] = ~layer_5[127] | (layer_5[117] & layer_5[127]); 
    assign layer_6[114] = layer_5[126] & layer_5[114]; 
    assign layer_6[115] = layer_5[98]; 
    assign layer_6[116] = layer_5[121] & layer_5[117]; 
    assign layer_6[117] = 1'b1; 
    assign layer_6[118] = ~layer_5[107] | (layer_5[107] & layer_5[122]); 
    assign layer_6[119] = layer_5[105] & ~layer_5[134]; 
    assign layer_6[120] = ~(layer_5[136] ^ layer_5[119]); 
    assign layer_6[121] = ~(layer_5[116] ^ layer_5[121]); 
    assign layer_6[122] = ~layer_5[135]; 
    assign layer_6[123] = ~(layer_5[139] ^ layer_5[129]); 
    assign layer_6[124] = ~(layer_5[135] ^ layer_5[111]); 
    assign layer_6[125] = ~(layer_5[128] ^ layer_5[139]); 
    assign layer_6[126] = layer_5[110]; 
    assign layer_6[127] = ~layer_5[114] | (layer_5[135] & layer_5[114]); 
    assign layer_6[128] = ~layer_5[114]; 
    assign layer_6[129] = layer_5[131]; 
    assign layer_6[130] = layer_5[125] & layer_5[126]; 
    assign layer_6[131] = layer_5[141] & layer_5[116]; 
    assign layer_6[132] = 1'b1; 
    assign layer_6[133] = 1'b1; 
    assign layer_6[134] = layer_5[119]; 
    assign layer_6[135] = ~(layer_5[148] ^ layer_5[123]); 
    assign layer_6[136] = ~layer_5[130]; 
    assign layer_6[137] = layer_5[129] & ~layer_5[129]; 
    assign layer_6[138] = ~layer_5[154]; 
    assign layer_6[139] = ~(layer_5[125] | layer_5[122]); 
    assign layer_6[140] = 1'b0; 
    assign layer_6[141] = layer_5[125] ^ layer_5[131]; 
    assign layer_6[142] = ~layer_5[132] | (layer_5[132] & layer_5[148]); 
    assign layer_6[143] = layer_5[154] ^ layer_5[133]; 
    assign layer_6[144] = 1'b0; 
    assign layer_6[145] = ~(layer_5[138] | layer_5[152]); 
    assign layer_6[146] = 1'b0; 
    assign layer_6[147] = layer_5[138] & ~layer_5[148]; 
    assign layer_6[148] = layer_5[146] ^ layer_5[137]; 
    assign layer_6[149] = layer_5[151] | layer_5[161]; 
    assign layer_6[150] = 1'b1; 
    assign layer_6[151] = layer_5[152]; 
    assign layer_6[152] = layer_5[166] ^ layer_5[159]; 
    assign layer_6[153] = layer_5[145]; 
    assign layer_6[154] = layer_5[164]; 
    assign layer_6[155] = 1'b0; 
    assign layer_6[156] = ~(layer_5[141] | layer_5[158]); 
    assign layer_6[157] = layer_5[151]; 
    assign layer_6[158] = 1'b0; 
    assign layer_6[159] = layer_5[146] & ~layer_5[165]; 
    assign layer_6[160] = ~(layer_5[152] ^ layer_5[152]); 
    assign layer_6[161] = 1'b0; 
    assign layer_6[162] = ~layer_5[153] | (layer_5[158] & layer_5[153]); 
    assign layer_6[163] = 1'b1; 
    assign layer_6[164] = ~layer_5[177] | (layer_5[177] & layer_5[149]); 
    assign layer_6[165] = ~layer_5[172]; 
    assign layer_6[166] = ~(layer_5[168] ^ layer_5[159]); 
    assign layer_6[167] = 1'b1; 
    assign layer_6[168] = ~(layer_5[160] & layer_5[162]); 
    assign layer_6[169] = layer_5[160] & ~layer_5[155]; 
    assign layer_6[170] = layer_5[155] & ~layer_5[162]; 
    assign layer_6[171] = ~(layer_5[181] ^ layer_5[176]); 
    assign layer_6[172] = layer_5[178]; 
    assign layer_6[173] = ~layer_5[188] | (layer_5[170] & layer_5[188]); 
    assign layer_6[174] = ~(layer_5[168] | layer_5[160]); 
    assign layer_6[175] = ~layer_5[176] | (layer_5[164] & layer_5[176]); 
    assign layer_6[176] = ~layer_5[189]; 
    assign layer_6[177] = ~(layer_5[178] | layer_5[177]); 
    assign layer_6[178] = ~layer_5[182]; 
    assign layer_6[179] = layer_5[166]; 
    assign layer_6[180] = layer_5[166]; 
    assign layer_6[181] = ~layer_5[168] | (layer_5[180] & layer_5[168]); 
    assign layer_6[182] = ~layer_5[175]; 
    assign layer_6[183] = layer_5[188]; 
    assign layer_6[184] = layer_5[198] & ~layer_5[176]; 
    assign layer_6[185] = layer_5[195]; 
    assign layer_6[186] = ~layer_5[198] | (layer_5[198] & layer_5[187]); 
    assign layer_6[187] = layer_5[179] ^ layer_5[184]; 
    assign layer_6[188] = layer_5[177] ^ layer_5[176]; 
    assign layer_6[189] = ~(layer_5[205] ^ layer_5[176]); 
    assign layer_6[190] = layer_5[177] | layer_5[203]; 
    assign layer_6[191] = ~(layer_5[207] ^ layer_5[200]); 
    assign layer_6[192] = ~(layer_5[180] & layer_5[194]); 
    assign layer_6[193] = ~(layer_5[204] | layer_5[180]); 
    assign layer_6[194] = ~(layer_5[181] ^ layer_5[193]); 
    assign layer_6[195] = layer_5[179]; 
    assign layer_6[196] = ~(layer_5[195] & layer_5[206]); 
    assign layer_6[197] = ~(layer_5[212] & layer_5[193]); 
    assign layer_6[198] = ~(layer_5[205] | layer_5[184]); 
    assign layer_6[199] = layer_5[191]; 
    assign layer_6[200] = 1'b1; 
    assign layer_6[201] = layer_5[213]; 
    assign layer_6[202] = ~(layer_5[212] ^ layer_5[189]); 
    assign layer_6[203] = layer_5[196] ^ layer_5[201]; 
    assign layer_6[204] = ~layer_5[189]; 
    assign layer_6[205] = layer_5[196] & ~layer_5[214]; 
    assign layer_6[206] = layer_5[211] & ~layer_5[212]; 
    assign layer_6[207] = layer_5[203] & layer_5[197]; 
    assign layer_6[208] = ~layer_5[192]; 
    assign layer_6[209] = 1'b1; 
    assign layer_6[210] = layer_5[222] & ~layer_5[208]; 
    assign layer_6[211] = ~(layer_5[204] ^ layer_5[223]); 
    assign layer_6[212] = ~layer_5[226]; 
    assign layer_6[213] = ~layer_5[226]; 
    assign layer_6[214] = ~(layer_5[223] | layer_5[225]); 
    assign layer_6[215] = layer_5[227] ^ layer_5[210]; 
    assign layer_6[216] = ~(layer_5[220] ^ layer_5[210]); 
    assign layer_6[217] = layer_5[210]; 
    assign layer_6[218] = layer_5[228] & layer_5[207]; 
    assign layer_6[219] = 1'b1; 
    assign layer_6[220] = ~(layer_5[221] & layer_5[226]); 
    assign layer_6[221] = ~layer_5[228] | (layer_5[228] & layer_5[213]); 
    assign layer_6[222] = layer_5[227] & ~layer_5[211]; 
    assign layer_6[223] = layer_5[225]; 
    assign layer_6[224] = layer_5[232] & ~layer_5[229]; 
    assign layer_6[225] = 1'b0; 
    assign layer_6[226] = ~(layer_5[241] | layer_5[213]); 
    assign layer_6[227] = ~layer_5[215]; 
    assign layer_6[228] = layer_5[239] ^ layer_5[235]; 
    assign layer_6[229] = layer_5[218] & ~layer_5[222]; 
    assign layer_6[230] = layer_5[233] | layer_5[232]; 
    assign layer_6[231] = ~(layer_5[218] ^ layer_5[218]); 
    assign layer_6[232] = ~layer_5[242]; 
    assign layer_6[233] = layer_5[226] & ~layer_5[233]; 
    assign layer_6[234] = layer_5[240] & ~layer_5[248]; 
    assign layer_6[235] = layer_5[236] & ~layer_5[233]; 
    assign layer_6[236] = layer_5[229] & ~layer_5[232]; 
    assign layer_6[237] = ~(layer_5[227] ^ layer_5[251]); 
    assign layer_6[238] = layer_5[233]; 
    assign layer_6[239] = layer_5[225]; 
    assign layer_6[240] = layer_5[232] ^ layer_5[225]; 
    assign layer_6[241] = layer_5[252]; 
    assign layer_6[242] = layer_5[235] & ~layer_5[248]; 
    assign layer_6[243] = layer_5[243]; 
    assign layer_6[244] = ~(layer_5[249] & layer_5[244]); 
    assign layer_6[245] = ~layer_5[240] | (layer_5[240] & layer_5[255]); 
    assign layer_6[246] = ~layer_5[258] | (layer_5[247] & layer_5[258]); 
    assign layer_6[247] = layer_5[240]; 
    assign layer_6[248] = layer_5[254] & ~layer_5[245]; 
    assign layer_6[249] = layer_5[240] & ~layer_5[240]; 
    assign layer_6[250] = ~(layer_5[252] & layer_5[258]); 
    assign layer_6[251] = ~(layer_5[261] ^ layer_5[251]); 
    assign layer_6[252] = layer_5[242] ^ layer_5[253]; 
    assign layer_6[253] = layer_5[237] & ~layer_5[252]; 
    assign layer_6[254] = layer_5[247] & ~layer_5[242]; 
    assign layer_6[255] = 1'b0; 
    assign layer_6[256] = layer_5[263] ^ layer_5[259]; 
    assign layer_6[257] = 1'b1; 
    assign layer_6[258] = 1'b1; 
    assign layer_6[259] = 1'b0; 
    assign layer_6[260] = layer_5[257]; 
    assign layer_6[261] = layer_5[256] | layer_5[251]; 
    assign layer_6[262] = ~layer_5[261]; 
    assign layer_6[263] = layer_5[265]; 
    assign layer_6[264] = ~layer_5[259] | (layer_5[259] & layer_5[265]); 
    assign layer_6[265] = layer_5[264] ^ layer_5[249]; 
    assign layer_6[266] = layer_5[281] & ~layer_5[255]; 
    assign layer_6[267] = layer_5[269]; 
    assign layer_6[268] = ~layer_5[272] | (layer_5[272] & layer_5[282]); 
    assign layer_6[269] = 1'b1; 
    assign layer_6[270] = 1'b0; 
    assign layer_6[271] = layer_5[261]; 
    assign layer_6[272] = 1'b0; 
    assign layer_6[273] = ~(layer_5[276] | layer_5[284]); 
    assign layer_6[274] = layer_5[273] & layer_5[268]; 
    assign layer_6[275] = layer_5[283] | layer_5[279]; 
    assign layer_6[276] = 1'b1; 
    assign layer_6[277] = ~layer_5[267] | (layer_5[292] & layer_5[267]); 
    assign layer_6[278] = ~layer_5[283] | (layer_5[283] & layer_5[291]); 
    assign layer_6[279] = ~(layer_5[287] ^ layer_5[282]); 
    assign layer_6[280] = ~layer_5[265] | (layer_5[270] & layer_5[265]); 
    assign layer_6[281] = layer_5[290]; 
    assign layer_6[282] = ~layer_5[295] | (layer_5[295] & layer_5[273]); 
    assign layer_6[283] = ~layer_5[276]; 
    assign layer_6[284] = layer_5[291]; 
    assign layer_6[285] = 1'b1; 
    assign layer_6[286] = ~layer_5[270] | (layer_5[288] & layer_5[270]); 
    assign layer_6[287] = layer_5[289] & layer_5[285]; 
    assign layer_6[288] = ~layer_5[279]; 
    assign layer_6[289] = layer_5[287]; 
    assign layer_6[290] = 1'b1; 
    assign layer_6[291] = ~layer_5[301] | (layer_5[301] & layer_5[282]); 
    assign layer_6[292] = ~(layer_5[281] & layer_5[290]); 
    assign layer_6[293] = ~(layer_5[296] ^ layer_5[290]); 
    assign layer_6[294] = layer_5[307]; 
    assign layer_6[295] = layer_5[286] & ~layer_5[286]; 
    assign layer_6[296] = layer_5[294] ^ layer_5[294]; 
    assign layer_6[297] = ~layer_5[287]; 
    assign layer_6[298] = ~layer_5[285] | (layer_5[285] & layer_5[286]); 
    assign layer_6[299] = ~layer_5[309] | (layer_5[306] & layer_5[309]); 
    assign layer_6[300] = layer_5[294] & ~layer_5[299]; 
    assign layer_6[301] = ~layer_5[294] | (layer_5[294] & layer_5[294]); 
    assign layer_6[302] = layer_5[301] & ~layer_5[290]; 
    assign layer_6[303] = layer_5[293] & ~layer_5[293]; 
    assign layer_6[304] = ~(layer_5[299] & layer_5[311]); 
    assign layer_6[305] = 1'b0; 
    assign layer_6[306] = layer_5[322]; 
    assign layer_6[307] = ~(layer_5[312] | layer_5[302]); 
    assign layer_6[308] = layer_5[312] | layer_5[294]; 
    assign layer_6[309] = ~(layer_5[309] & layer_5[296]); 
    assign layer_6[310] = layer_5[316] ^ layer_5[309]; 
    assign layer_6[311] = ~layer_5[327] | (layer_5[327] & layer_5[325]); 
    assign layer_6[312] = ~layer_5[313] | (layer_5[325] & layer_5[313]); 
    assign layer_6[313] = layer_5[315] | layer_5[316]; 
    assign layer_6[314] = layer_5[304] ^ layer_5[324]; 
    assign layer_6[315] = ~layer_5[327] | (layer_5[325] & layer_5[327]); 
    assign layer_6[316] = layer_5[323]; 
    assign layer_6[317] = layer_5[300]; 
    assign layer_6[318] = layer_5[302] & ~layer_5[303]; 
    assign layer_6[319] = layer_5[311] & ~layer_5[322]; 
    assign layer_6[320] = 1'b0; 
    assign layer_6[321] = ~layer_5[327] | (layer_5[329] & layer_5[327]); 
    assign layer_6[322] = ~layer_5[326]; 
    assign layer_6[323] = layer_5[313] | layer_5[315]; 
    assign layer_6[324] = ~layer_5[339] | (layer_5[339] & layer_5[316]); 
    assign layer_6[325] = layer_5[337] & ~layer_5[334]; 
    assign layer_6[326] = 1'b1; 
    assign layer_6[327] = layer_5[336]; 
    assign layer_6[328] = ~(layer_5[327] | layer_5[314]); 
    assign layer_6[329] = 1'b0; 
    assign layer_6[330] = layer_5[324]; 
    assign layer_6[331] = ~layer_5[331] | (layer_5[331] & layer_5[338]); 
    assign layer_6[332] = ~layer_5[342]; 
    assign layer_6[333] = ~layer_5[346] | (layer_5[335] & layer_5[346]); 
    assign layer_6[334] = ~layer_5[323]; 
    assign layer_6[335] = layer_5[329] ^ layer_5[320]; 
    assign layer_6[336] = layer_5[339]; 
    assign layer_6[337] = 1'b0; 
    assign layer_6[338] = layer_5[324] & ~layer_5[321]; 
    assign layer_6[339] = ~(layer_5[329] ^ layer_5[326]); 
    assign layer_6[340] = layer_5[354]; 
    assign layer_6[341] = ~(layer_5[325] | layer_5[350]); 
    assign layer_6[342] = layer_5[328]; 
    assign layer_6[343] = layer_5[330] | layer_5[356]; 
    assign layer_6[344] = 1'b1; 
    assign layer_6[345] = ~(layer_5[347] | layer_5[342]); 
    assign layer_6[346] = ~layer_5[356] | (layer_5[349] & layer_5[356]); 
    assign layer_6[347] = layer_5[340] & ~layer_5[362]; 
    assign layer_6[348] = layer_5[360]; 
    assign layer_6[349] = layer_5[360] & ~layer_5[339]; 
    assign layer_6[350] = ~(layer_5[336] | layer_5[342]); 
    assign layer_6[351] = ~layer_5[363]; 
    assign layer_6[352] = layer_5[344] | layer_5[344]; 
    assign layer_6[353] = layer_5[338] ^ layer_5[337]; 
    assign layer_6[354] = ~(layer_5[369] ^ layer_5[347]); 
    assign layer_6[355] = ~layer_5[361] | (layer_5[361] & layer_5[350]); 
    assign layer_6[356] = layer_5[362] ^ layer_5[344]; 
    assign layer_6[357] = layer_5[372]; 
    assign layer_6[358] = ~layer_5[352] | (layer_5[365] & layer_5[352]); 
    assign layer_6[359] = ~layer_5[371] | (layer_5[347] & layer_5[371]); 
    assign layer_6[360] = 1'b0; 
    assign layer_6[361] = ~layer_5[357] | (layer_5[357] & layer_5[348]); 
    assign layer_6[362] = ~layer_5[362]; 
    assign layer_6[363] = 1'b1; 
    assign layer_6[364] = layer_5[364] | layer_5[377]; 
    assign layer_6[365] = layer_5[359] & layer_5[351]; 
    assign layer_6[366] = ~layer_5[367]; 
    assign layer_6[367] = 1'b1; 
    assign layer_6[368] = 1'b0; 
    assign layer_6[369] = layer_5[362] & ~layer_5[359]; 
    assign layer_6[370] = layer_5[386] & layer_5[358]; 
    assign layer_6[371] = ~(layer_5[387] | layer_5[365]); 
    assign layer_6[372] = 1'b1; 
    assign layer_6[373] = layer_5[361]; 
    assign layer_6[374] = layer_5[371] & ~layer_5[372]; 
    assign layer_6[375] = layer_5[383] ^ layer_5[381]; 
    assign layer_6[376] = ~(layer_5[373] | layer_5[362]); 
    assign layer_6[377] = ~(layer_5[383] | layer_5[375]); 
    assign layer_6[378] = ~layer_5[374] | (layer_5[363] & layer_5[374]); 
    assign layer_6[379] = 1'b0; 
    assign layer_6[380] = ~(layer_5[378] ^ layer_5[367]); 
    assign layer_6[381] = layer_5[383] & ~layer_5[384]; 
    assign layer_6[382] = ~(layer_5[390] | layer_5[394]); 
    assign layer_6[383] = ~layer_5[367]; 
    assign layer_6[384] = layer_5[377] | layer_5[374]; 
    assign layer_6[385] = ~layer_5[372]; 
    assign layer_6[386] = ~layer_5[384] | (layer_5[384] & layer_5[385]); 
    assign layer_6[387] = ~(layer_5[386] | layer_5[373]); 
    assign layer_6[388] = layer_5[388]; 
    assign layer_6[389] = layer_5[404] & ~layer_5[393]; 
    assign layer_6[390] = ~layer_5[376]; 
    assign layer_6[391] = layer_5[402] | layer_5[381]; 
    assign layer_6[392] = layer_5[396] & ~layer_5[392]; 
    assign layer_6[393] = ~layer_5[387]; 
    assign layer_6[394] = layer_5[398]; 
    assign layer_6[395] = layer_5[382]; 
    assign layer_6[396] = ~layer_5[386]; 
    assign layer_6[397] = layer_5[383]; 
    assign layer_6[398] = ~(layer_5[403] & layer_5[388]); 
    assign layer_6[399] = 1'b1; 
    assign layer_6[400] = layer_5[405]; 
    assign layer_6[401] = 1'b1; 
    assign layer_6[402] = ~layer_5[415]; 
    assign layer_6[403] = ~layer_5[393] | (layer_5[393] & layer_5[416]); 
    assign layer_6[404] = ~layer_5[409]; 
    assign layer_6[405] = ~layer_5[414] | (layer_5[414] & layer_5[416]); 
    assign layer_6[406] = 1'b1; 
    assign layer_6[407] = layer_5[397]; 
    assign layer_6[408] = ~layer_5[408] | (layer_5[408] & layer_5[392]); 
    assign layer_6[409] = ~layer_5[410] | (layer_5[410] & layer_5[394]); 
    assign layer_6[410] = 1'b0; 
    assign layer_6[411] = layer_5[422]; 
    assign layer_6[412] = ~(layer_5[426] & layer_5[404]); 
    assign layer_6[413] = ~(layer_5[420] & layer_5[409]); 
    assign layer_6[414] = layer_5[399] & layer_5[401]; 
    assign layer_6[415] = layer_5[420] & ~layer_5[410]; 
    assign layer_6[416] = layer_5[402] & ~layer_5[410]; 
    assign layer_6[417] = layer_5[427] | layer_5[407]; 
    assign layer_6[418] = layer_5[408] & ~layer_5[430]; 
    assign layer_6[419] = ~layer_5[406] | (layer_5[423] & layer_5[406]); 
    assign layer_6[420] = ~(layer_5[426] ^ layer_5[416]); 
    assign layer_6[421] = layer_5[432]; 
    assign layer_6[422] = ~layer_5[437]; 
    assign layer_6[423] = ~(layer_5[434] & layer_5[438]); 
    assign layer_6[424] = layer_5[423] & ~layer_5[408]; 
    assign layer_6[425] = 1'b1; 
    assign layer_6[426] = layer_5[425] ^ layer_5[421]; 
    assign layer_6[427] = layer_5[424]; 
    assign layer_6[428] = 1'b0; 
    assign layer_6[429] = layer_5[431] & layer_5[426]; 
    assign layer_6[430] = ~layer_5[439] | (layer_5[439] & layer_5[421]); 
    assign layer_6[431] = layer_5[427] | layer_5[431]; 
    assign layer_6[432] = layer_5[448] ^ layer_5[422]; 
    assign layer_6[433] = layer_5[441]; 
    assign layer_6[434] = ~layer_5[436] | (layer_5[433] & layer_5[436]); 
    assign layer_6[435] = ~(layer_5[439] & layer_5[431]); 
    assign layer_6[436] = ~layer_5[432] | (layer_5[432] & layer_5[431]); 
    assign layer_6[437] = layer_5[449] & ~layer_5[441]; 
    assign layer_6[438] = layer_5[443] & ~layer_5[425]; 
    assign layer_6[439] = layer_5[427] & ~layer_5[451]; 
    assign layer_6[440] = layer_5[434] & ~layer_5[450]; 
    assign layer_6[441] = layer_5[455] & layer_5[433]; 
    assign layer_6[442] = layer_5[451] ^ layer_5[427]; 
    assign layer_6[443] = ~(layer_5[429] & layer_5[435]); 
    assign layer_6[444] = 1'b1; 
    assign layer_6[445] = ~layer_5[456] | (layer_5[435] & layer_5[456]); 
    assign layer_6[446] = 1'b0; 
    assign layer_6[447] = layer_5[446] | layer_5[433]; 
    assign layer_6[448] = ~layer_5[451] | (layer_5[449] & layer_5[451]); 
    assign layer_6[449] = ~layer_5[435] | (layer_5[435] & layer_5[436]); 
    assign layer_6[450] = layer_5[435] ^ layer_5[436]; 
    assign layer_6[451] = ~layer_5[447]; 
    assign layer_6[452] = ~layer_5[437] | (layer_5[437] & layer_5[457]); 
    assign layer_6[453] = layer_5[448] & layer_5[466]; 
    assign layer_6[454] = 1'b0; 
    assign layer_6[455] = ~layer_5[439] | (layer_5[439] & layer_5[446]); 
    assign layer_6[456] = ~layer_5[466] | (layer_5[466] & layer_5[463]); 
    assign layer_6[457] = layer_5[456] & layer_5[447]; 
    assign layer_6[458] = 1'b0; 
    assign layer_6[459] = 1'b1; 
    assign layer_6[460] = 1'b0; 
    assign layer_6[461] = 1'b1; 
    assign layer_6[462] = ~layer_5[462] | (layer_5[476] & layer_5[462]); 
    assign layer_6[463] = ~layer_5[464]; 
    assign layer_6[464] = layer_5[476] ^ layer_5[475]; 
    assign layer_6[465] = ~layer_5[480] | (layer_5[480] & layer_5[474]); 
    assign layer_6[466] = layer_5[457] & ~layer_5[468]; 
    assign layer_6[467] = ~layer_5[461]; 
    assign layer_6[468] = ~layer_5[466] | (layer_5[466] & layer_5[453]); 
    assign layer_6[469] = layer_5[468]; 
    assign layer_6[470] = ~(layer_5[459] ^ layer_5[468]); 
    assign layer_6[471] = layer_5[460]; 
    assign layer_6[472] = layer_5[457] & ~layer_5[455]; 
    assign layer_6[473] = ~layer_5[471]; 
    assign layer_6[474] = ~layer_5[458] | (layer_5[475] & layer_5[458]); 
    assign layer_6[475] = ~layer_5[479] | (layer_5[491] & layer_5[479]); 
    assign layer_6[476] = 1'b1; 
    assign layer_6[477] = ~layer_5[479] | (layer_5[487] & layer_5[479]); 
    assign layer_6[478] = 1'b0; 
    assign layer_6[479] = layer_5[480] & layer_5[478]; 
    assign layer_6[480] = ~(layer_5[492] & layer_5[469]); 
    assign layer_6[481] = layer_5[482] & ~layer_5[470]; 
    assign layer_6[482] = ~layer_5[478] | (layer_5[478] & layer_5[488]); 
    assign layer_6[483] = layer_5[469]; 
    assign layer_6[484] = layer_5[496]; 
    assign layer_6[485] = 1'b1; 
    assign layer_6[486] = layer_5[471] ^ layer_5[501]; 
    assign layer_6[487] = ~(layer_5[493] & layer_5[473]); 
    assign layer_6[488] = ~(layer_5[475] ^ layer_5[502]); 
    assign layer_6[489] = 1'b1; 
    assign layer_6[490] = 1'b0; 
    assign layer_6[491] = layer_5[503]; 
    assign layer_6[492] = ~layer_5[499]; 
    assign layer_6[493] = ~(layer_5[485] & layer_5[498]); 
    assign layer_6[494] = ~(layer_5[478] | layer_5[499]); 
    assign layer_6[495] = 1'b1; 
    assign layer_6[496] = layer_5[491]; 
    assign layer_6[497] = layer_5[490] ^ layer_5[510]; 
    assign layer_6[498] = ~layer_5[499] | (layer_5[484] & layer_5[499]); 
    assign layer_6[499] = layer_5[507]; 
    assign layer_6[500] = 1'b0; 
    assign layer_6[501] = layer_5[492] | layer_5[512]; 
    assign layer_6[502] = layer_5[517] | layer_5[511]; 
    assign layer_6[503] = layer_5[512]; 
    assign layer_6[504] = layer_5[495]; 
    assign layer_6[505] = ~(layer_5[494] | layer_5[508]); 
    assign layer_6[506] = ~(layer_5[498] | layer_5[512]); 
    assign layer_6[507] = layer_5[507] & ~layer_5[516]; 
    assign layer_6[508] = layer_5[513] ^ layer_5[515]; 
    assign layer_6[509] = ~layer_5[519] | (layer_5[496] & layer_5[519]); 
    assign layer_6[510] = layer_5[519]; 
    assign layer_6[511] = ~layer_5[511] | (layer_5[511] & layer_5[516]); 
    assign layer_6[512] = ~(layer_5[510] ^ layer_5[516]); 
    assign layer_6[513] = ~(layer_5[512] & layer_5[521]); 
    assign layer_6[514] = layer_5[529] | layer_5[510]; 
    assign layer_6[515] = ~(layer_5[499] | layer_5[503]); 
    assign layer_6[516] = ~(layer_5[513] | layer_5[523]); 
    assign layer_6[517] = ~(layer_5[517] ^ layer_5[526]); 
    assign layer_6[518] = layer_5[506] & layer_5[519]; 
    assign layer_6[519] = 1'b0; 
    assign layer_6[520] = layer_5[516] & ~layer_5[504]; 
    assign layer_6[521] = 1'b1; 
    assign layer_6[522] = ~layer_5[523]; 
    assign layer_6[523] = 1'b0; 
    assign layer_6[524] = layer_5[524] | layer_5[539]; 
    assign layer_6[525] = ~(layer_5[531] | layer_5[512]); 
    assign layer_6[526] = 1'b1; 
    assign layer_6[527] = ~layer_5[526]; 
    assign layer_6[528] = layer_5[523] & ~layer_5[517]; 
    assign layer_6[529] = ~layer_5[535]; 
    assign layer_6[530] = ~(layer_5[535] ^ layer_5[533]); 
    assign layer_6[531] = layer_5[531] & ~layer_5[515]; 
    assign layer_6[532] = ~layer_5[517]; 
    assign layer_6[533] = layer_5[533] & layer_5[547]; 
    assign layer_6[534] = layer_5[535] & ~layer_5[530]; 
    assign layer_6[535] = layer_5[537]; 
    assign layer_6[536] = ~(layer_5[549] ^ layer_5[527]); 
    assign layer_6[537] = 1'b1; 
    assign layer_6[538] = ~layer_5[543] | (layer_5[534] & layer_5[543]); 
    assign layer_6[539] = ~(layer_5[541] & layer_5[532]); 
    assign layer_6[540] = layer_5[550]; 
    assign layer_6[541] = layer_5[541] & layer_5[540]; 
    assign layer_6[542] = ~layer_5[543]; 
    assign layer_6[543] = ~layer_5[530] | (layer_5[530] & layer_5[554]); 
    assign layer_6[544] = layer_5[548] ^ layer_5[533]; 
    assign layer_6[545] = layer_5[558] | layer_5[554]; 
    assign layer_6[546] = ~(layer_5[561] | layer_5[543]); 
    assign layer_6[547] = layer_5[549] & ~layer_5[543]; 
    assign layer_6[548] = ~(layer_5[559] ^ layer_5[550]); 
    assign layer_6[549] = 1'b1; 
    assign layer_6[550] = layer_5[565] & ~layer_5[538]; 
    assign layer_6[551] = layer_5[537] & ~layer_5[561]; 
    assign layer_6[552] = layer_5[567] & ~layer_5[553]; 
    assign layer_6[553] = layer_5[546]; 
    assign layer_6[554] = layer_5[563]; 
    assign layer_6[555] = layer_5[555]; 
    assign layer_6[556] = ~layer_5[570] | (layer_5[557] & layer_5[570]); 
    assign layer_6[557] = ~layer_5[563]; 
    assign layer_6[558] = layer_5[563]; 
    assign layer_6[559] = ~layer_5[571] | (layer_5[571] & layer_5[557]); 
    assign layer_6[560] = 1'b0; 
    assign layer_6[561] = ~layer_5[553]; 
    assign layer_6[562] = ~(layer_5[564] ^ layer_5[577]); 
    assign layer_6[563] = layer_5[557] & ~layer_5[568]; 
    assign layer_6[564] = layer_5[551] ^ layer_5[559]; 
    assign layer_6[565] = layer_5[579]; 
    assign layer_6[566] = layer_5[552] & layer_5[575]; 
    assign layer_6[567] = layer_5[565] & layer_5[560]; 
    assign layer_6[568] = 1'b0; 
    assign layer_6[569] = layer_5[564] ^ layer_5[569]; 
    assign layer_6[570] = ~layer_5[579] | (layer_5[579] & layer_5[555]); 
    assign layer_6[571] = ~(layer_5[586] ^ layer_5[581]); 
    assign layer_6[572] = ~layer_5[570] | (layer_5[570] & layer_5[565]); 
    assign layer_6[573] = layer_5[558]; 
    assign layer_6[574] = layer_5[583] & layer_5[559]; 
    assign layer_6[575] = layer_5[575]; 
    assign layer_6[576] = layer_5[576]; 
    assign layer_6[577] = layer_5[570] ^ layer_5[560]; 
    assign layer_6[578] = 1'b1; 
    assign layer_6[579] = layer_5[588]; 
    assign layer_6[580] = ~layer_5[563]; 
    assign layer_6[581] = 1'b1; 
    assign layer_6[582] = layer_5[592] & layer_5[590]; 
    assign layer_6[583] = layer_5[571]; 
    assign layer_6[584] = layer_5[595]; 
    assign layer_6[585] = ~(layer_5[576] & layer_5[568]); 
    assign layer_6[586] = ~layer_5[589] | (layer_5[589] & layer_5[574]); 
    assign layer_6[587] = ~(layer_5[583] | layer_5[576]); 
    assign layer_6[588] = layer_5[593] & ~layer_5[577]; 
    assign layer_6[589] = ~(layer_5[598] ^ layer_5[584]); 
    assign layer_6[590] = layer_5[595] | layer_5[596]; 
    assign layer_6[591] = layer_5[580] & ~layer_5[596]; 
    assign layer_6[592] = ~layer_5[591]; 
    assign layer_6[593] = layer_5[589]; 
    assign layer_6[594] = layer_5[581] & ~layer_5[596]; 
    assign layer_6[595] = ~layer_5[580]; 
    assign layer_6[596] = layer_5[608] | layer_5[597]; 
    assign layer_6[597] = 1'b1; 
    assign layer_6[598] = ~layer_5[586]; 
    assign layer_6[599] = layer_5[609]; 
    assign layer_6[600] = 1'b0; 
    assign layer_6[601] = layer_5[590]; 
    assign layer_6[602] = ~layer_5[613]; 
    assign layer_6[603] = ~(layer_5[592] ^ layer_5[601]); 
    assign layer_6[604] = ~(layer_5[588] ^ layer_5[611]); 
    assign layer_6[605] = ~layer_5[602]; 
    assign layer_6[606] = ~layer_5[610] | (layer_5[612] & layer_5[610]); 
    assign layer_6[607] = layer_5[612] & ~layer_5[592]; 
    assign layer_6[608] = ~layer_5[608] | (layer_5[608] & layer_5[600]); 
    assign layer_6[609] = ~layer_5[615]; 
    assign layer_6[610] = layer_5[594]; 
    assign layer_6[611] = layer_5[601] & ~layer_5[599]; 
    assign layer_6[612] = layer_5[617] & ~layer_5[618]; 
    assign layer_6[613] = ~layer_5[605]; 
    assign layer_6[614] = 1'b0; 
    assign layer_6[615] = 1'b0; 
    assign layer_6[616] = ~layer_5[603] | (layer_5[603] & layer_5[624]); 
    assign layer_6[617] = ~layer_5[611] | (layer_5[611] & layer_5[605]); 
    assign layer_6[618] = layer_5[611] | layer_5[609]; 
    assign layer_6[619] = ~layer_5[614]; 
    assign layer_6[620] = layer_5[616] & layer_5[603]; 
    assign layer_6[621] = ~(layer_5[616] ^ layer_5[633]); 
    assign layer_6[622] = layer_5[621]; 
    assign layer_6[623] = ~(layer_5[617] & layer_5[611]); 
    assign layer_6[624] = 1'b0; 
    assign layer_6[625] = ~layer_5[636]; 
    assign layer_6[626] = layer_5[620] | layer_5[619]; 
    assign layer_6[627] = ~layer_5[619] | (layer_5[619] & layer_5[621]); 
    assign layer_6[628] = layer_5[617]; 
    assign layer_6[629] = 1'b0; 
    assign layer_6[630] = layer_5[626] | layer_5[617]; 
    assign layer_6[631] = ~layer_5[644]; 
    assign layer_6[632] = layer_5[626] | layer_5[640]; 
    assign layer_6[633] = ~layer_5[649] | (layer_5[649] & layer_5[632]); 
    assign layer_6[634] = layer_5[627]; 
    assign layer_6[635] = layer_5[633] | layer_5[629]; 
    assign layer_6[636] = layer_5[628]; 
    assign layer_6[637] = ~(layer_5[639] | layer_5[650]); 
    assign layer_6[638] = layer_5[626] & ~layer_5[640]; 
    assign layer_6[639] = ~(layer_5[628] | layer_5[648]); 
    assign layer_6[640] = layer_5[655] & ~layer_5[647]; 
    assign layer_6[641] = ~layer_5[639] | (layer_5[639] & layer_5[636]); 
    assign layer_6[642] = ~layer_5[637]; 
    assign layer_6[643] = ~layer_5[627]; 
    assign layer_6[644] = layer_5[632] & layer_5[627]; 
    assign layer_6[645] = ~layer_5[649]; 
    assign layer_6[646] = layer_5[637] ^ layer_5[640]; 
    assign layer_6[647] = ~layer_5[631] | (layer_5[636] & layer_5[631]); 
    assign layer_6[648] = ~layer_5[641]; 
    assign layer_6[649] = layer_5[653]; 
    assign layer_6[650] = layer_5[666]; 
    assign layer_6[651] = layer_5[664]; 
    assign layer_6[652] = layer_5[662]; 
    assign layer_6[653] = ~layer_5[646]; 
    assign layer_6[654] = 1'b0; 
    assign layer_6[655] = layer_5[662] & ~layer_5[653]; 
    assign layer_6[656] = layer_5[643]; 
    assign layer_6[657] = ~layer_5[645]; 
    assign layer_6[658] = layer_5[648] & layer_5[672]; 
    assign layer_6[659] = layer_5[670] & ~layer_5[667]; 
    assign layer_6[660] = ~layer_5[672] | (layer_5[672] & layer_5[648]); 
    assign layer_6[661] = ~(layer_5[660] ^ layer_5[649]); 
    assign layer_6[662] = layer_5[668]; 
    assign layer_6[663] = ~(layer_5[664] & layer_5[648]); 
    assign layer_6[664] = ~layer_5[664] | (layer_5[679] & layer_5[664]); 
    assign layer_6[665] = layer_5[670] ^ layer_5[671]; 
    assign layer_6[666] = ~(layer_5[667] | layer_5[657]); 
    assign layer_6[667] = layer_5[664] & ~layer_5[673]; 
    assign layer_6[668] = layer_5[669] & ~layer_5[670]; 
    assign layer_6[669] = layer_5[666] & layer_5[671]; 
    assign layer_6[670] = layer_5[674] & ~layer_5[679]; 
    assign layer_6[671] = ~(layer_5[685] | layer_5[667]); 
    assign layer_6[672] = 1'b1; 
    assign layer_6[673] = 1'b0; 
    assign layer_6[674] = 1'b1; 
    assign layer_6[675] = layer_5[687] | layer_5[677]; 
    assign layer_6[676] = layer_5[660] & layer_5[684]; 
    assign layer_6[677] = layer_5[678] ^ layer_5[667]; 
    assign layer_6[678] = ~layer_5[669]; 
    assign layer_6[679] = ~layer_5[662] | (layer_5[675] & layer_5[662]); 
    assign layer_6[680] = layer_5[665] & ~layer_5[670]; 
    assign layer_6[681] = layer_5[686] & layer_5[696]; 
    assign layer_6[682] = ~layer_5[692]; 
    assign layer_6[683] = layer_5[693] ^ layer_5[670]; 
    assign layer_6[684] = ~layer_5[687] | (layer_5[687] & layer_5[693]); 
    assign layer_6[685] = layer_5[697] | layer_5[675]; 
    assign layer_6[686] = ~layer_5[685]; 
    assign layer_6[687] = ~layer_5[688] | (layer_5[688] & layer_5[688]); 
    assign layer_6[688] = ~(layer_5[674] | layer_5[700]); 
    assign layer_6[689] = ~(layer_5[698] | layer_5[672]); 
    assign layer_6[690] = ~layer_5[680] | (layer_5[685] & layer_5[680]); 
    assign layer_6[691] = ~(layer_5[701] & layer_5[692]); 
    assign layer_6[692] = layer_5[681]; 
    assign layer_6[693] = ~layer_5[707] | (layer_5[696] & layer_5[707]); 
    assign layer_6[694] = 1'b0; 
    assign layer_6[695] = ~layer_5[691]; 
    assign layer_6[696] = ~(layer_5[696] ^ layer_5[683]); 
    assign layer_6[697] = ~layer_5[682]; 
    assign layer_6[698] = ~(layer_5[697] ^ layer_5[689]); 
    assign layer_6[699] = 1'b0; 
    assign layer_6[700] = ~(layer_5[705] & layer_5[693]); 
    assign layer_6[701] = 1'b0; 
    assign layer_6[702] = 1'b0; 
    assign layer_6[703] = layer_5[709] | layer_5[686]; 
    assign layer_6[704] = ~(layer_5[716] ^ layer_5[702]); 
    assign layer_6[705] = layer_5[714]; 
    assign layer_6[706] = layer_5[702] | layer_5[703]; 
    assign layer_6[707] = layer_5[713] ^ layer_5[704]; 
    assign layer_6[708] = layer_5[705] & layer_5[707]; 
    assign layer_6[709] = ~(layer_5[709] ^ layer_5[719]); 
    assign layer_6[710] = layer_5[712] ^ layer_5[725]; 
    assign layer_6[711] = 1'b0; 
    assign layer_6[712] = layer_5[698] | layer_5[701]; 
    assign layer_6[713] = layer_5[717] | layer_5[698]; 
    assign layer_6[714] = layer_5[706] | layer_5[709]; 
    assign layer_6[715] = 1'b1; 
    assign layer_6[716] = ~(layer_5[706] | layer_5[702]); 
    assign layer_6[717] = layer_5[715]; 
    assign layer_6[718] = layer_5[715] | layer_5[709]; 
    assign layer_6[719] = ~(layer_5[724] ^ layer_5[726]); 
    assign layer_6[720] = layer_5[713] & ~layer_5[725]; 
    assign layer_6[721] = 1'b1; 
    assign layer_6[722] = layer_5[713] ^ layer_5[713]; 
    assign layer_6[723] = 1'b0; 
    assign layer_6[724] = layer_5[725]; 
    assign layer_6[725] = layer_5[732] ^ layer_5[713]; 
    assign layer_6[726] = layer_5[715]; 
    assign layer_6[727] = ~layer_5[731]; 
    assign layer_6[728] = ~layer_5[738] | (layer_5[726] & layer_5[738]); 
    assign layer_6[729] = 1'b0; 
    assign layer_6[730] = layer_5[714] | layer_5[713]; 
    assign layer_6[731] = layer_5[727]; 
    assign layer_6[732] = layer_5[737] ^ layer_5[737]; 
    assign layer_6[733] = ~(layer_5[747] & layer_5[719]); 
    assign layer_6[734] = layer_5[746] | layer_5[747]; 
    assign layer_6[735] = layer_5[746] ^ layer_5[744]; 
    assign layer_6[736] = layer_5[727] ^ layer_5[722]; 
    assign layer_6[737] = ~layer_5[750] | (layer_5[723] & layer_5[750]); 
    assign layer_6[738] = layer_5[743] & ~layer_5[734]; 
    assign layer_6[739] = layer_5[741]; 
    assign layer_6[740] = layer_5[725] & ~layer_5[725]; 
    assign layer_6[741] = ~layer_5[748] | (layer_5[733] & layer_5[748]); 
    assign layer_6[742] = layer_5[757] ^ layer_5[754]; 
    assign layer_6[743] = 1'b0; 
    assign layer_6[744] = layer_5[754] & layer_5[735]; 
    assign layer_6[745] = layer_5[758]; 
    assign layer_6[746] = 1'b1; 
    assign layer_6[747] = 1'b1; 
    assign layer_6[748] = layer_5[759]; 
    assign layer_6[749] = ~(layer_5[764] & layer_5[743]); 
    assign layer_6[750] = layer_5[737]; 
    assign layer_6[751] = ~layer_5[760]; 
    assign layer_6[752] = ~layer_5[742] | (layer_5[742] & layer_5[739]); 
    assign layer_6[753] = ~layer_5[756] | (layer_5[756] & layer_5[750]); 
    assign layer_6[754] = ~(layer_5[742] | layer_5[755]); 
    assign layer_6[755] = layer_5[746] & ~layer_5[755]; 
    assign layer_6[756] = ~(layer_5[751] ^ layer_5[765]); 
    assign layer_6[757] = ~layer_5[742]; 
    assign layer_6[758] = ~layer_5[769]; 
    assign layer_6[759] = layer_5[757] ^ layer_5[773]; 
    assign layer_6[760] = layer_5[757] & ~layer_5[775]; 
    assign layer_6[761] = ~(layer_5[763] ^ layer_5[763]); 
    assign layer_6[762] = ~(layer_5[770] ^ layer_5[769]); 
    assign layer_6[763] = layer_5[777] & ~layer_5[766]; 
    assign layer_6[764] = layer_5[774] & ~layer_5[774]; 
    assign layer_6[765] = layer_5[772] & ~layer_5[766]; 
    assign layer_6[766] = 1'b0; 
    assign layer_6[767] = ~(layer_5[765] ^ layer_5[763]); 
    assign layer_6[768] = ~layer_5[762] | (layer_5[762] & layer_5[768]); 
    assign layer_6[769] = layer_5[759]; 
    assign layer_6[770] = layer_5[778]; 
    assign layer_6[771] = 1'b1; 
    assign layer_6[772] = layer_5[775]; 
    assign layer_6[773] = layer_5[767]; 
    assign layer_6[774] = ~(layer_5[772] | layer_5[766]); 
    assign layer_6[775] = layer_5[771] | layer_5[773]; 
    assign layer_6[776] = layer_5[776] & layer_5[791]; 
    assign layer_6[777] = layer_5[768] | layer_5[772]; 
    assign layer_6[778] = ~(layer_5[764] & layer_5[762]); 
    assign layer_6[779] = layer_5[771] & ~layer_5[793]; 
    assign layer_6[780] = layer_5[763]; 
    assign layer_6[781] = ~(layer_5[792] ^ layer_5[786]); 
    assign layer_6[782] = 1'b1; 
    assign layer_6[783] = 1'b0; 
    assign layer_6[784] = layer_5[771] & layer_5[789]; 
    assign layer_6[785] = layer_5[771] & ~layer_5[790]; 
    assign layer_6[786] = ~(layer_5[796] & layer_5[789]); 
    assign layer_6[787] = layer_5[775] & ~layer_5[771]; 
    assign layer_6[788] = layer_5[797] & ~layer_5[798]; 
    assign layer_6[789] = ~layer_5[780]; 
    assign layer_6[790] = ~(layer_5[785] & layer_5[773]); 
    assign layer_6[791] = ~(layer_5[784] & layer_5[778]); 
    assign layer_6[792] = layer_5[798] ^ layer_5[787]; 
    assign layer_6[793] = 1'b1; 
    assign layer_6[794] = ~layer_5[800] | (layer_5[804] & layer_5[800]); 
    assign layer_6[795] = layer_5[790]; 
    assign layer_6[796] = ~layer_5[788] | (layer_5[796] & layer_5[788]); 
    assign layer_6[797] = layer_5[812] ^ layer_5[804]; 
    assign layer_6[798] = ~layer_5[813]; 
    assign layer_6[799] = ~(layer_5[802] | layer_5[795]); 
    assign layer_6[800] = layer_5[808] & ~layer_5[815]; 
    assign layer_6[801] = ~(layer_5[795] & layer_5[784]); 
    assign layer_6[802] = ~(layer_5[812] | layer_5[801]); 
    assign layer_6[803] = 1'b1; 
    assign layer_6[804] = ~layer_5[809]; 
    assign layer_6[805] = ~layer_5[807]; 
    assign layer_6[806] = 1'b1; 
    assign layer_6[807] = ~(layer_5[798] & layer_5[806]); 
    assign layer_6[808] = layer_5[823]; 
    assign layer_6[809] = layer_5[805] ^ layer_5[818]; 
    assign layer_6[810] = 1'b0; 
    assign layer_6[811] = 1'b1; 
    assign layer_6[812] = layer_5[813]; 
    assign layer_6[813] = layer_5[803]; 
    assign layer_6[814] = layer_5[807] | layer_5[814]; 
    assign layer_6[815] = ~(layer_5[800] ^ layer_5[815]); 
    assign layer_6[816] = ~layer_5[823] | (layer_5[823] & layer_5[801]); 
    assign layer_6[817] = layer_5[808]; 
    assign layer_6[818] = layer_5[823] | layer_5[823]; 
    assign layer_6[819] = layer_5[808]; 
    assign layer_6[820] = ~(layer_5[812] & layer_5[819]); 
    assign layer_6[821] = ~(layer_5[828] & layer_5[804]); 
    assign layer_6[822] = ~(layer_5[807] ^ layer_5[824]); 
    assign layer_6[823] = layer_5[839] ^ layer_5[807]; 
    assign layer_6[824] = layer_5[814]; 
    assign layer_6[825] = ~(layer_5[828] | layer_5[813]); 
    assign layer_6[826] = layer_5[829]; 
    assign layer_6[827] = layer_5[816] | layer_5[833]; 
    assign layer_6[828] = ~layer_5[813] | (layer_5[840] & layer_5[813]); 
    assign layer_6[829] = 1'b0; 
    assign layer_6[830] = layer_5[846] & ~layer_5[837]; 
    assign layer_6[831] = 1'b1; 
    assign layer_6[832] = layer_5[819]; 
    assign layer_6[833] = layer_5[841] ^ layer_5[825]; 
    assign layer_6[834] = layer_5[829] & layer_5[839]; 
    assign layer_6[835] = 1'b1; 
    assign layer_6[836] = layer_5[828]; 
    assign layer_6[837] = layer_5[832]; 
    assign layer_6[838] = ~layer_5[828] | (layer_5[846] & layer_5[828]); 
    assign layer_6[839] = ~layer_5[837]; 
    assign layer_6[840] = 1'b0; 
    assign layer_6[841] = 1'b1; 
    assign layer_6[842] = layer_5[839] & ~layer_5[835]; 
    assign layer_6[843] = layer_5[851] & ~layer_5[858]; 
    assign layer_6[844] = ~layer_5[841] | (layer_5[841] & layer_5[842]); 
    assign layer_6[845] = layer_5[861] & layer_5[854]; 
    assign layer_6[846] = layer_5[854] & ~layer_5[848]; 
    assign layer_6[847] = 1'b1; 
    assign layer_6[848] = ~(layer_5[839] | layer_5[849]); 
    assign layer_6[849] = ~layer_5[847]; 
    assign layer_6[850] = ~layer_5[836]; 
    assign layer_6[851] = layer_5[850] & ~layer_5[846]; 
    assign layer_6[852] = ~(layer_5[864] & layer_5[859]); 
    assign layer_6[853] = ~layer_5[839] | (layer_5[839] & layer_5[857]); 
    assign layer_6[854] = 1'b0; 
    assign layer_6[855] = ~(layer_5[866] ^ layer_5[854]); 
    assign layer_6[856] = 1'b0; 
    assign layer_6[857] = ~(layer_5[846] | layer_5[862]); 
    assign layer_6[858] = ~(layer_5[865] & layer_5[855]); 
    assign layer_6[859] = layer_5[856] & ~layer_5[855]; 
    assign layer_6[860] = layer_5[862] ^ layer_5[862]; 
    assign layer_6[861] = layer_5[865] | layer_5[860]; 
    assign layer_6[862] = layer_5[869] & layer_5[865]; 
    assign layer_6[863] = layer_5[876] & ~layer_5[847]; 
    assign layer_6[864] = ~layer_5[847] | (layer_5[869] & layer_5[847]); 
    assign layer_6[865] = ~layer_5[875] | (layer_5[875] & layer_5[875]); 
    assign layer_6[866] = layer_5[872] ^ layer_5[881]; 
    assign layer_6[867] = layer_5[868]; 
    assign layer_6[868] = 1'b0; 
    assign layer_6[869] = 1'b0; 
    assign layer_6[870] = layer_5[878] & layer_5[868]; 
    assign layer_6[871] = layer_5[863] & ~layer_5[861]; 
    assign layer_6[872] = 1'b0; 
    assign layer_6[873] = layer_5[858] & layer_5[870]; 
    assign layer_6[874] = ~layer_5[867]; 
    assign layer_6[875] = layer_5[890] & ~layer_5[862]; 
    assign layer_6[876] = ~(layer_5[888] & layer_5[879]); 
    assign layer_6[877] = ~layer_5[879] | (layer_5[869] & layer_5[879]); 
    assign layer_6[878] = ~(layer_5[874] ^ layer_5[886]); 
    assign layer_6[879] = 1'b0; 
    assign layer_6[880] = layer_5[872] & ~layer_5[881]; 
    assign layer_6[881] = ~layer_5[864] | (layer_5[872] & layer_5[864]); 
    assign layer_6[882] = ~layer_5[897]; 
    assign layer_6[883] = layer_5[885] ^ layer_5[893]; 
    assign layer_6[884] = layer_5[875] & ~layer_5[886]; 
    assign layer_6[885] = ~layer_5[871] | (layer_5[893] & layer_5[871]); 
    assign layer_6[886] = layer_5[887] | layer_5[893]; 
    assign layer_6[887] = ~(layer_5[878] ^ layer_5[896]); 
    assign layer_6[888] = ~layer_5[878]; 
    assign layer_6[889] = ~(layer_5[882] | layer_5[882]); 
    assign layer_6[890] = layer_5[880]; 
    assign layer_6[891] = 1'b1; 
    assign layer_6[892] = layer_5[908]; 
    assign layer_6[893] = ~(layer_5[883] & layer_5[893]); 
    assign layer_6[894] = ~(layer_5[904] & layer_5[904]); 
    assign layer_6[895] = ~(layer_5[888] | layer_5[886]); 
    assign layer_6[896] = layer_5[881] | layer_5[910]; 
    assign layer_6[897] = ~(layer_5[905] & layer_5[902]); 
    assign layer_6[898] = layer_5[901] & ~layer_5[914]; 
    assign layer_6[899] = 1'b1; 
    assign layer_6[900] = ~(layer_5[896] | layer_5[902]); 
    assign layer_6[901] = layer_5[901]; 
    assign layer_6[902] = 1'b1; 
    assign layer_6[903] = ~(layer_5[901] ^ layer_5[899]); 
    assign layer_6[904] = layer_5[902] | layer_5[916]; 
    assign layer_6[905] = layer_5[911] & ~layer_5[917]; 
    assign layer_6[906] = layer_5[919] & layer_5[893]; 
    assign layer_6[907] = layer_5[894] & layer_5[897]; 
    assign layer_6[908] = ~layer_5[923]; 
    assign layer_6[909] = layer_5[895] & ~layer_5[897]; 
    assign layer_6[910] = ~layer_5[901] | (layer_5[901] & layer_5[907]); 
    assign layer_6[911] = layer_5[903] ^ layer_5[915]; 
    assign layer_6[912] = layer_5[898] & ~layer_5[918]; 
    assign layer_6[913] = layer_5[923] & ~layer_5[926]; 
    assign layer_6[914] = ~layer_5[909]; 
    assign layer_6[915] = layer_5[905] & layer_5[913]; 
    assign layer_6[916] = layer_5[909] | layer_5[923]; 
    assign layer_6[917] = 1'b1; 
    assign layer_6[918] = layer_5[922] & ~layer_5[926]; 
    assign layer_6[919] = layer_5[914] & layer_5[913]; 
    assign layer_6[920] = ~layer_5[909]; 
    assign layer_6[921] = layer_5[908] & layer_5[912]; 
    assign layer_6[922] = layer_5[935] ^ layer_5[924]; 
    assign layer_6[923] = ~layer_5[908] | (layer_5[907] & layer_5[908]); 
    assign layer_6[924] = layer_5[938]; 
    assign layer_6[925] = 1'b0; 
    assign layer_6[926] = layer_5[929]; 
    assign layer_6[927] = layer_5[942]; 
    assign layer_6[928] = ~layer_5[913] | (layer_5[919] & layer_5[913]); 
    assign layer_6[929] = ~(layer_5[931] & layer_5[943]); 
    assign layer_6[930] = 1'b0; 
    assign layer_6[931] = layer_5[918]; 
    assign layer_6[932] = ~layer_5[923]; 
    assign layer_6[933] = layer_5[937] | layer_5[939]; 
    assign layer_6[934] = layer_5[940]; 
    assign layer_6[935] = layer_5[947] & ~layer_5[946]; 
    assign layer_6[936] = layer_5[947] & ~layer_5[928]; 
    assign layer_6[937] = layer_5[946]; 
    assign layer_6[938] = ~(layer_5[953] | layer_5[949]); 
    assign layer_6[939] = layer_5[953] & ~layer_5[936]; 
    assign layer_6[940] = layer_5[924]; 
    assign layer_6[941] = ~layer_5[952]; 
    assign layer_6[942] = layer_5[930] | layer_5[946]; 
    assign layer_6[943] = ~(layer_5[959] | layer_5[928]); 
    assign layer_6[944] = 1'b1; 
    assign layer_6[945] = ~layer_5[941] | (layer_5[935] & layer_5[941]); 
    assign layer_6[946] = 1'b1; 
    assign layer_6[947] = layer_5[931] & layer_5[930]; 
    assign layer_6[948] = ~(layer_5[934] & layer_5[940]); 
    assign layer_6[949] = 1'b0; 
    assign layer_6[950] = layer_5[950]; 
    assign layer_6[951] = ~(layer_5[938] & layer_5[949]); 
    assign layer_6[952] = ~layer_5[968]; 
    assign layer_6[953] = layer_5[957] & ~layer_5[944]; 
    assign layer_6[954] = layer_5[944] & layer_5[948]; 
    assign layer_6[955] = 1'b1; 
    assign layer_6[956] = ~(layer_5[945] & layer_5[946]); 
    assign layer_6[957] = layer_5[970] | layer_5[955]; 
    assign layer_6[958] = layer_5[972] | layer_5[952]; 
    assign layer_6[959] = ~(layer_5[957] ^ layer_5[957]); 
    assign layer_6[960] = 1'b1; 
    assign layer_6[961] = ~(layer_5[954] ^ layer_5[955]); 
    assign layer_6[962] = layer_5[975] & ~layer_5[968]; 
    assign layer_6[963] = ~layer_5[966]; 
    assign layer_6[964] = 1'b0; 
    assign layer_6[965] = 1'b0; 
    assign layer_6[966] = ~layer_5[970]; 
    assign layer_6[967] = layer_5[968] | layer_5[961]; 
    assign layer_6[968] = layer_5[962] ^ layer_5[970]; 
    assign layer_6[969] = layer_5[983] & ~layer_5[953]; 
    assign layer_6[970] = layer_5[962] & ~layer_5[958]; 
    assign layer_6[971] = ~(layer_5[956] ^ layer_5[963]); 
    assign layer_6[972] = 1'b1; 
    assign layer_6[973] = 1'b1; 
    assign layer_6[974] = ~layer_5[970]; 
    assign layer_6[975] = layer_5[966] | layer_5[990]; 
    assign layer_6[976] = layer_5[984] & ~layer_5[988]; 
    assign layer_6[977] = ~layer_5[986] | (layer_5[986] & layer_5[962]); 
    assign layer_6[978] = layer_5[981]; 
    assign layer_6[979] = ~layer_5[967] | (layer_5[976] & layer_5[967]); 
    assign layer_6[980] = layer_5[970]; 
    assign layer_6[981] = ~layer_5[972]; 
    assign layer_6[982] = 1'b0; 
    assign layer_6[983] = ~layer_5[987] | (layer_5[971] & layer_5[987]); 
    assign layer_6[984] = ~(layer_5[995] | layer_5[977]); 
    assign layer_6[985] = layer_5[985] & layer_5[1000]; 
    assign layer_6[986] = ~(layer_5[1002] & layer_5[990]); 
    assign layer_6[987] = ~layer_5[983] | (layer_5[983] & layer_5[972]); 
    assign layer_6[988] = ~layer_5[1002] | (layer_5[1002] & layer_5[976]); 
    assign layer_6[989] = layer_5[990]; 
    assign layer_6[990] = ~(layer_5[981] & layer_5[1002]); 
    assign layer_6[991] = layer_5[982]; 
    assign layer_6[992] = layer_5[986] & layer_5[983]; 
    assign layer_6[993] = layer_5[989]; 
    assign layer_6[994] = layer_5[1003] & ~layer_5[1001]; 
    assign layer_6[995] = ~(layer_5[980] ^ layer_5[979]); 
    assign layer_6[996] = ~(layer_5[984] & layer_5[979]); 
    assign layer_6[997] = ~layer_5[991]; 
    assign layer_6[998] = ~layer_5[986] | (layer_5[994] & layer_5[986]); 
    assign layer_6[999] = layer_5[990] | layer_5[1004]; 
    assign layer_6[1000] = layer_5[1011]; 
    assign layer_6[1001] = ~(layer_5[1011] ^ layer_5[984]); 
    assign layer_6[1002] = layer_5[1003] | layer_5[998]; 
    assign layer_6[1003] = ~(layer_5[988] | layer_5[1012]); 
    assign layer_6[1004] = ~(layer_5[1019] & layer_5[1008]); 
    assign layer_6[1005] = layer_5[993] & layer_5[1018]; 
    assign layer_6[1006] = ~layer_5[1014] | (layer_5[1014] & layer_5[998]); 
    assign layer_6[1007] = 1'b1; 
    assign layer_6[1008] = ~layer_5[1022]; 
    assign layer_6[1009] = ~(layer_5[1022] | layer_5[1022]); 
    assign layer_6[1010] = ~(layer_5[1014] | layer_5[1018]); 
    assign layer_6[1011] = ~layer_5[995] | (layer_5[995] & layer_5[1006]); 
    assign layer_6[1012] = layer_5[1018] ^ layer_5[999]; 
    assign layer_6[1013] = layer_5[1002] & layer_5[1002]; 
    assign layer_6[1014] = layer_5[1008]; 
    assign layer_6[1015] = layer_5[1019] | layer_5[1017]; 
    assign layer_6[1016] = 1'b0; 
    assign layer_6[1017] = layer_5[1020]; 
    assign layer_6[1018] = ~layer_5[1017] | (layer_5[1017] & layer_5[1018]); 
    assign layer_6[1019] = ~(layer_5[1006] & layer_5[1019]); 
    assign layer_6[1020] = ~layer_5[1006]; 
    assign layer_6[1021] = layer_5[1011] | layer_5[1023]; 
    assign layer_6[1022] = layer_5[1019]; 
    assign layer_6[1023] = ~layer_5[1019]; 
    // Layer 7 ============================================================
    assign out[0] = layer_6[13] | layer_6[16]; 
    assign out[1] = ~layer_6[15] | (layer_6[7] & layer_6[15]); 
    assign out[2] = ~(layer_6[4] ^ layer_6[1]); 
    assign out[3] = layer_6[6]; 
    assign out[4] = layer_6[10] & ~layer_6[1]; 
    assign out[5] = ~layer_6[20]; 
    assign out[6] = ~(layer_6[3] & layer_6[5]); 
    assign out[7] = layer_6[6] & ~layer_6[10]; 
    assign out[8] = layer_6[2] & layer_6[1]; 
    assign out[9] = layer_6[22] ^ layer_6[5]; 
    assign out[10] = ~layer_6[2]; 
    assign out[11] = layer_6[21] & layer_6[15]; 
    assign out[12] = layer_6[22] ^ layer_6[1]; 
    assign out[13] = ~layer_6[1] | (layer_6[12] & layer_6[1]); 
    assign out[14] = ~(layer_6[0] | layer_6[18]); 
    assign out[15] = ~layer_6[16] | (layer_6[9] & layer_6[16]); 
    assign out[16] = ~layer_6[3]; 
    assign out[17] = ~layer_6[14]; 
    assign out[18] = ~layer_6[34]; 
    assign out[19] = layer_6[24] ^ layer_6[8]; 
    assign out[20] = layer_6[29]; 
    assign out[21] = ~layer_6[18] | (layer_6[18] & layer_6[10]); 
    assign out[22] = layer_6[36] | layer_6[9]; 
    assign out[23] = layer_6[34] & ~layer_6[21]; 
    assign out[24] = ~(layer_6[11] | layer_6[23]); 
    assign out[25] = 1'b1; 
    assign out[26] = layer_6[25] & ~layer_6[19]; 
    assign out[27] = layer_6[11] & ~layer_6[11]; 
    assign out[28] = 1'b0; 
    assign out[29] = layer_6[21] & ~layer_6[33]; 
    assign out[30] = layer_6[15] & ~layer_6[14]; 
    assign out[31] = ~layer_6[23] | (layer_6[23] & layer_6[20]); 
    assign out[32] = layer_6[34]; 
    assign out[33] = ~(layer_6[35] & layer_6[41]); 
    assign out[34] = layer_6[48]; 
    assign out[35] = layer_6[43] ^ layer_6[43]; 
    assign out[36] = ~(layer_6[21] ^ layer_6[32]); 
    assign out[37] = ~(layer_6[40] & layer_6[22]); 
    assign out[38] = 1'b1; 
    assign out[39] = layer_6[49] & layer_6[47]; 
    assign out[40] = layer_6[30] ^ layer_6[35]; 
    assign out[41] = ~layer_6[28]; 
    assign out[42] = ~layer_6[37] | (layer_6[37] & layer_6[53]); 
    assign out[43] = ~layer_6[42]; 
    assign out[44] = layer_6[37]; 
    assign out[45] = layer_6[61] ^ layer_6[44]; 
    assign out[46] = ~(layer_6[59] | layer_6[57]); 
    assign out[47] = ~layer_6[33] | (layer_6[40] & layer_6[33]); 
    assign out[48] = layer_6[36]; 
    assign out[49] = layer_6[48] & layer_6[42]; 
    assign out[50] = layer_6[52] | layer_6[55]; 
    assign out[51] = ~(layer_6[56] ^ layer_6[40]); 
    assign out[52] = layer_6[65] & ~layer_6[47]; 
    assign out[53] = ~(layer_6[41] & layer_6[41]); 
    assign out[54] = ~layer_6[48] | (layer_6[39] & layer_6[48]); 
    assign out[55] = ~(layer_6[53] | layer_6[54]); 
    assign out[56] = ~layer_6[56]; 
    assign out[57] = ~(layer_6[47] ^ layer_6[54]); 
    assign out[58] = ~(layer_6[42] & layer_6[55]); 
    assign out[59] = ~layer_6[70]; 
    assign out[60] = layer_6[65]; 
    assign out[61] = ~(layer_6[51] & layer_6[74]); 
    assign out[62] = ~layer_6[74] | (layer_6[74] & layer_6[46]); 
    assign out[63] = layer_6[68]; 
    assign out[64] = ~(layer_6[68] ^ layer_6[71]); 
    assign out[65] = layer_6[50] | layer_6[58]; 
    assign out[66] = layer_6[62] | layer_6[60]; 
    assign out[67] = ~layer_6[55]; 
    assign out[68] = layer_6[67] ^ layer_6[64]; 
    assign out[69] = layer_6[83]; 
    assign out[70] = layer_6[70]; 
    assign out[71] = ~(layer_6[70] | layer_6[73]); 
    assign out[72] = 1'b0; 
    assign out[73] = ~layer_6[60]; 
    assign out[74] = layer_6[77] ^ layer_6[69]; 
    assign out[75] = layer_6[64] ^ layer_6[74]; 
    assign out[76] = ~(layer_6[78] & layer_6[61]); 
    assign out[77] = layer_6[64]; 
    assign out[78] = ~layer_6[71] | (layer_6[71] & layer_6[71]); 
    assign out[79] = layer_6[89] & ~layer_6[92]; 
    assign out[80] = ~layer_6[82] | (layer_6[82] & layer_6[63]); 
    assign out[81] = layer_6[95] ^ layer_6[86]; 
    assign out[82] = ~(layer_6[93] | layer_6[75]); 
    assign out[83] = ~layer_6[87]; 
    assign out[84] = ~(layer_6[94] & layer_6[96]); 
    assign out[85] = layer_6[99] & layer_6[87]; 
    assign out[86] = layer_6[71] ^ layer_6[84]; 
    assign out[87] = layer_6[88]; 
    assign out[88] = 1'b1; 
    assign out[89] = layer_6[103]; 
    assign out[90] = 1'b0; 
    assign out[91] = ~layer_6[86]; 
    assign out[92] = ~(layer_6[86] & layer_6[75]); 
    assign out[93] = 1'b1; 
    assign out[94] = ~(layer_6[78] | layer_6[83]); 
    assign out[95] = layer_6[80]; 
    assign out[96] = ~(layer_6[99] & layer_6[100]); 
    assign out[97] = layer_6[101] & ~layer_6[113]; 
    assign out[98] = layer_6[102] & ~layer_6[86]; 
    assign out[99] = layer_6[111]; 
    assign out[100] = ~(layer_6[114] ^ layer_6[86]); 
    assign out[101] = 1'b0; 
    assign out[102] = layer_6[95] ^ layer_6[100]; 
    assign out[103] = layer_6[117] ^ layer_6[87]; 
    assign out[104] = layer_6[113]; 
    assign out[105] = ~(layer_6[91] ^ layer_6[91]); 
    assign out[106] = 1'b1; 
    assign out[107] = layer_6[111] ^ layer_6[99]; 
    assign out[108] = ~(layer_6[107] ^ layer_6[106]); 
    assign out[109] = layer_6[112]; 
    assign out[110] = layer_6[119] & ~layer_6[114]; 
    assign out[111] = layer_6[119]; 
    assign out[112] = ~layer_6[116]; 
    assign out[113] = 1'b0; 
    assign out[114] = layer_6[124] & ~layer_6[129]; 
    assign out[115] = layer_6[113] | layer_6[125]; 
    assign out[116] = 1'b1; 
    assign out[117] = ~(layer_6[128] & layer_6[106]); 
    assign out[118] = layer_6[110] ^ layer_6[111]; 
    assign out[119] = ~layer_6[105] | (layer_6[129] & layer_6[105]); 
    assign out[120] = 1'b0; 
    assign out[121] = layer_6[122]; 
    assign out[122] = layer_6[121] & ~layer_6[123]; 
    assign out[123] = ~(layer_6[120] & layer_6[125]); 
    assign out[124] = layer_6[114] & ~layer_6[124]; 
    assign out[125] = ~(layer_6[116] & layer_6[130]); 
    assign out[126] = layer_6[142] | layer_6[109]; 
    assign out[127] = layer_6[131] | layer_6[127]; 
    assign out[128] = ~layer_6[114] | (layer_6[114] & layer_6[129]); 
    assign out[129] = ~(layer_6[144] | layer_6[138]); 
    assign out[130] = layer_6[140] | layer_6[121]; 
    assign out[131] = 1'b1; 
    assign out[132] = 1'b0; 
    assign out[133] = layer_6[140] & layer_6[118]; 
    assign out[134] = ~layer_6[131] | (layer_6[137] & layer_6[131]); 
    assign out[135] = ~layer_6[127]; 
    assign out[136] = ~layer_6[148] | (layer_6[148] & layer_6[145]); 
    assign out[137] = ~(layer_6[131] & layer_6[152]); 
    assign out[138] = layer_6[144] ^ layer_6[151]; 
    assign out[139] = layer_6[141] ^ layer_6[131]; 
    assign out[140] = layer_6[134]; 
    assign out[141] = layer_6[150] | layer_6[144]; 
    assign out[142] = layer_6[143]; 
    assign out[143] = 1'b0; 
    assign out[144] = layer_6[156]; 
    assign out[145] = layer_6[134]; 
    assign out[146] = 1'b0; 
    assign out[147] = 1'b0; 
    assign out[148] = layer_6[138]; 
    assign out[149] = layer_6[152]; 
    assign out[150] = 1'b0; 
    assign out[151] = ~layer_6[163]; 
    assign out[152] = layer_6[165]; 
    assign out[153] = 1'b1; 
    assign out[154] = 1'b0; 
    assign out[155] = layer_6[171] ^ layer_6[144]; 
    assign out[156] = ~layer_6[163]; 
    assign out[157] = ~layer_6[154] | (layer_6[154] & layer_6[162]); 
    assign out[158] = ~(layer_6[155] ^ layer_6[166]); 
    assign out[159] = ~layer_6[157] | (layer_6[164] & layer_6[157]); 
    assign out[160] = layer_6[176] | layer_6[172]; 
    assign out[161] = 1'b0; 
    assign out[162] = ~layer_6[159] | (layer_6[167] & layer_6[159]); 
    assign out[163] = layer_6[173] ^ layer_6[154]; 
    assign out[164] = layer_6[157] & layer_6[153]; 
    assign out[165] = layer_6[164] | layer_6[164]; 
    assign out[166] = ~(layer_6[171] & layer_6[168]); 
    assign out[167] = layer_6[155] ^ layer_6[156]; 
    assign out[168] = layer_6[181] | layer_6[180]; 
    assign out[169] = ~layer_6[156]; 
    assign out[170] = 1'b1; 
    assign out[171] = ~(layer_6[163] | layer_6[174]); 
    assign out[172] = ~(layer_6[187] | layer_6[168]); 
    assign out[173] = ~layer_6[165]; 
    assign out[174] = 1'b1; 
    assign out[175] = layer_6[177] | layer_6[177]; 
    assign out[176] = ~(layer_6[168] | layer_6[180]); 
    assign out[177] = layer_6[182] & ~layer_6[181]; 
    assign out[178] = ~layer_6[171] | (layer_6[180] & layer_6[171]); 
    assign out[179] = layer_6[178] & ~layer_6[189]; 
    assign out[180] = layer_6[178]; 
    assign out[181] = ~layer_6[169] | (layer_6[180] & layer_6[169]); 
    assign out[182] = layer_6[181]; 
    assign out[183] = layer_6[182] | layer_6[190]; 
    assign out[184] = ~layer_6[169]; 
    assign out[185] = layer_6[199]; 
    assign out[186] = ~(layer_6[198] ^ layer_6[182]); 
    assign out[187] = layer_6[189] ^ layer_6[172]; 
    assign out[188] = layer_6[175] & ~layer_6[197]; 
    assign out[189] = ~(layer_6[181] ^ layer_6[180]); 
    assign out[190] = ~layer_6[204]; 
    assign out[191] = ~(layer_6[188] | layer_6[205]); 
    assign out[192] = ~(layer_6[187] & layer_6[180]); 
    assign out[193] = layer_6[207] & ~layer_6[205]; 
    assign out[194] = ~(layer_6[178] & layer_6[183]); 
    assign out[195] = ~layer_6[191]; 
    assign out[196] = ~layer_6[206]; 
    assign out[197] = ~(layer_6[208] ^ layer_6[209]); 
    assign out[198] = ~layer_6[186]; 
    assign out[199] = ~(layer_6[190] ^ layer_6[187]); 
    assign out[200] = ~layer_6[208]; 
    assign out[201] = ~layer_6[186]; 
    assign out[202] = layer_6[198] | layer_6[189]; 
    assign out[203] = layer_6[198] & layer_6[198]; 
    assign out[204] = layer_6[216] ^ layer_6[190]; 
    assign out[205] = layer_6[207] & ~layer_6[209]; 
    assign out[206] = layer_6[202] & ~layer_6[205]; 
    assign out[207] = ~layer_6[214] | (layer_6[216] & layer_6[214]); 
    assign out[208] = 1'b1; 
    assign out[209] = ~(layer_6[206] | layer_6[196]); 
    assign out[210] = ~layer_6[212]; 
    assign out[211] = ~layer_6[221] | (layer_6[223] & layer_6[221]); 
    assign out[212] = ~(layer_6[215] | layer_6[222]); 
    assign out[213] = layer_6[216]; 
    assign out[214] = ~layer_6[216] | (layer_6[224] & layer_6[216]); 
    assign out[215] = ~layer_6[202]; 
    assign out[216] = 1'b1; 
    assign out[217] = layer_6[215] & layer_6[208]; 
    assign out[218] = layer_6[208] ^ layer_6[204]; 
    assign out[219] = layer_6[215] | layer_6[234]; 
    assign out[220] = ~layer_6[220] | (layer_6[220] & layer_6[230]); 
    assign out[221] = ~(layer_6[211] | layer_6[204]); 
    assign out[222] = ~layer_6[235] | (layer_6[223] & layer_6[235]); 
    assign out[223] = 1'b1; 
    assign out[224] = ~layer_6[224]; 
    assign out[225] = ~layer_6[237] | (layer_6[237] & layer_6[224]); 
    assign out[226] = layer_6[223] & ~layer_6[239]; 
    assign out[227] = layer_6[212] & ~layer_6[225]; 
    assign out[228] = 1'b1; 
    assign out[229] = ~layer_6[220]; 
    assign out[230] = ~layer_6[214] | (layer_6[214] & layer_6[233]); 
    assign out[231] = layer_6[220] ^ layer_6[215]; 
    assign out[232] = ~(layer_6[233] | layer_6[223]); 
    assign out[233] = layer_6[217] & ~layer_6[221]; 
    assign out[234] = layer_6[218] & ~layer_6[232]; 
    assign out[235] = layer_6[251] & ~layer_6[223]; 
    assign out[236] = ~layer_6[241] | (layer_6[241] & layer_6[226]); 
    assign out[237] = ~(layer_6[234] | layer_6[221]); 
    assign out[238] = ~(layer_6[246] | layer_6[228]); 
    assign out[239] = ~(layer_6[225] ^ layer_6[223]); 
    assign out[240] = ~layer_6[244] | (layer_6[244] & layer_6[243]); 
    assign out[241] = ~layer_6[247] | (layer_6[243] & layer_6[247]); 
    assign out[242] = ~layer_6[253]; 
    assign out[243] = ~(layer_6[250] & layer_6[231]); 
    assign out[244] = ~layer_6[232]; 
    assign out[245] = ~layer_6[236] | (layer_6[236] & layer_6[245]); 
    assign out[246] = 1'b1; 
    assign out[247] = ~layer_6[241]; 
    assign out[248] = layer_6[255]; 
    assign out[249] = layer_6[245] ^ layer_6[261]; 
    assign out[250] = ~(layer_6[234] ^ layer_6[247]); 
    assign out[251] = ~(layer_6[249] ^ layer_6[265]); 
    assign out[252] = layer_6[257]; 
    assign out[253] = ~layer_6[243] | (layer_6[250] & layer_6[243]); 
    assign out[254] = layer_6[246]; 
    assign out[255] = ~layer_6[250]; 
    assign out[256] = layer_6[265] & ~layer_6[259]; 
    assign out[257] = ~layer_6[267]; 
    assign out[258] = ~layer_6[256]; 
    assign out[259] = ~(layer_6[253] | layer_6[248]); 
    assign out[260] = ~layer_6[275]; 
    assign out[261] = layer_6[263] ^ layer_6[244]; 
    assign out[262] = layer_6[268] & layer_6[277]; 
    assign out[263] = layer_6[277]; 
    assign out[264] = layer_6[252]; 
    assign out[265] = layer_6[270]; 
    assign out[266] = ~layer_6[264]; 
    assign out[267] = layer_6[254] ^ layer_6[277]; 
    assign out[268] = ~(layer_6[264] | layer_6[275]); 
    assign out[269] = ~layer_6[262]; 
    assign out[270] = ~(layer_6[284] ^ layer_6[261]); 
    assign out[271] = layer_6[269] & ~layer_6[278]; 
    assign out[272] = layer_6[261] & ~layer_6[288]; 
    assign out[273] = ~(layer_6[289] ^ layer_6[269]); 
    assign out[274] = layer_6[260] & ~layer_6[276]; 
    assign out[275] = layer_6[274]; 
    assign out[276] = layer_6[278] & ~layer_6[287]; 
    assign out[277] = layer_6[270] & ~layer_6[292]; 
    assign out[278] = 1'b0; 
    assign out[279] = 1'b0; 
    assign out[280] = layer_6[271] & ~layer_6[284]; 
    assign out[281] = ~layer_6[269] | (layer_6[297] & layer_6[269]); 
    assign out[282] = layer_6[287] & layer_6[291]; 
    assign out[283] = layer_6[286] | layer_6[281]; 
    assign out[284] = 1'b0; 
    assign out[285] = ~layer_6[285]; 
    assign out[286] = ~layer_6[296]; 
    assign out[287] = layer_6[296] | layer_6[292]; 
    assign out[288] = ~(layer_6[288] & layer_6[280]); 
    assign out[289] = ~layer_6[276]; 
    assign out[290] = ~(layer_6[304] & layer_6[302]); 
    assign out[291] = 1'b1; 
    assign out[292] = ~layer_6[291] | (layer_6[299] & layer_6[291]); 
    assign out[293] = layer_6[304] ^ layer_6[292]; 
    assign out[294] = layer_6[288]; 
    assign out[295] = 1'b1; 
    assign out[296] = layer_6[280]; 
    assign out[297] = layer_6[290] | layer_6[283]; 
    assign out[298] = layer_6[297] & ~layer_6[306]; 
    assign out[299] = layer_6[299] | layer_6[306]; 
    assign out[300] = ~(layer_6[311] ^ layer_6[290]); 
    assign out[301] = layer_6[296] & ~layer_6[292]; 
    assign out[302] = ~(layer_6[288] & layer_6[316]); 
    assign out[303] = 1'b0; 
    assign out[304] = layer_6[305] | layer_6[291]; 
    assign out[305] = layer_6[318]; 
    assign out[306] = ~layer_6[312] | (layer_6[312] & layer_6[306]); 
    assign out[307] = layer_6[311] | layer_6[321]; 
    assign out[308] = layer_6[294] | layer_6[306]; 
    assign out[309] = layer_6[324]; 
    assign out[310] = ~layer_6[320]; 
    assign out[311] = ~layer_6[300] | (layer_6[300] & layer_6[318]); 
    assign out[312] = layer_6[319] & layer_6[312]; 
    assign out[313] = ~layer_6[308]; 
    assign out[314] = 1'b0; 
    assign out[315] = layer_6[299] | layer_6[322]; 
    assign out[316] = ~(layer_6[312] | layer_6[301]); 
    assign out[317] = ~layer_6[327]; 
    assign out[318] = layer_6[317] & layer_6[306]; 
    assign out[319] = layer_6[317] | layer_6[327]; 
    assign out[320] = layer_6[305] & ~layer_6[321]; 
    assign out[321] = layer_6[308] & ~layer_6[335]; 
    assign out[322] = ~layer_6[311]; 
    assign out[323] = ~(layer_6[322] ^ layer_6[335]); 
    assign out[324] = ~(layer_6[321] ^ layer_6[311]); 
    assign out[325] = ~(layer_6[336] & layer_6[338]); 
    assign out[326] = 1'b0; 
    assign out[327] = layer_6[326] ^ layer_6[317]; 
    assign out[328] = layer_6[335] & ~layer_6[330]; 
    assign out[329] = ~layer_6[326]; 
    assign out[330] = layer_6[318] | layer_6[340]; 
    assign out[331] = ~(layer_6[323] & layer_6[319]); 
    assign out[332] = ~layer_6[343] | (layer_6[342] & layer_6[343]); 
    assign out[333] = 1'b0; 
    assign out[334] = ~layer_6[325] | (layer_6[325] & layer_6[335]); 
    assign out[335] = ~(layer_6[339] | layer_6[339]); 
    assign out[336] = ~layer_6[343]; 
    assign out[337] = layer_6[331] ^ layer_6[326]; 
    assign out[338] = ~layer_6[346]; 
    assign out[339] = layer_6[355] ^ layer_6[334]; 
    assign out[340] = layer_6[334]; 
    assign out[341] = ~layer_6[338]; 
    assign out[342] = ~(layer_6[348] & layer_6[347]); 
    assign out[343] = layer_6[329] | layer_6[341]; 
    assign out[344] = layer_6[350] ^ layer_6[332]; 
    assign out[345] = layer_6[360] | layer_6[359]; 
    assign out[346] = layer_6[349] & layer_6[338]; 
    assign out[347] = layer_6[358]; 
    assign out[348] = ~layer_6[332] | (layer_6[342] & layer_6[332]); 
    assign out[349] = 1'b0; 
    assign out[350] = 1'b1; 
    assign out[351] = ~(layer_6[345] ^ layer_6[365]); 
    assign out[352] = ~(layer_6[368] ^ layer_6[338]); 
    assign out[353] = ~layer_6[343]; 
    assign out[354] = ~layer_6[348]; 
    assign out[355] = ~layer_6[347] | (layer_6[340] & layer_6[347]); 
    assign out[356] = ~(layer_6[349] | layer_6[358]); 
    assign out[357] = ~(layer_6[369] | layer_6[362]); 
    assign out[358] = layer_6[346]; 
    assign out[359] = ~(layer_6[375] & layer_6[353]); 
    assign out[360] = layer_6[356] | layer_6[357]; 
    assign out[361] = ~(layer_6[346] ^ layer_6[373]); 
    assign out[362] = layer_6[359] ^ layer_6[371]; 
    assign out[363] = layer_6[356] & ~layer_6[358]; 
    assign out[364] = ~layer_6[360]; 
    assign out[365] = 1'b0; 
    assign out[366] = layer_6[377]; 
    assign out[367] = ~layer_6[360]; 
    assign out[368] = layer_6[379] & ~layer_6[366]; 
    assign out[369] = ~layer_6[362]; 
    assign out[370] = layer_6[357] | layer_6[384]; 
    assign out[371] = ~(layer_6[365] | layer_6[358]); 
    assign out[372] = layer_6[374] | layer_6[387]; 
    assign out[373] = ~(layer_6[389] | layer_6[362]); 
    assign out[374] = layer_6[377] | layer_6[360]; 
    assign out[375] = layer_6[367] ^ layer_6[389]; 
    assign out[376] = ~layer_6[360]; 
    assign out[377] = layer_6[385]; 
    assign out[378] = ~(layer_6[369] ^ layer_6[392]); 
    assign out[379] = ~layer_6[392]; 
    assign out[380] = ~layer_6[381] | (layer_6[370] & layer_6[381]); 
    assign out[381] = layer_6[390] | layer_6[373]; 
    assign out[382] = ~(layer_6[386] | layer_6[389]); 
    assign out[383] = ~layer_6[378] | (layer_6[378] & layer_6[371]); 
    assign out[384] = layer_6[370] & ~layer_6[393]; 
    assign out[385] = ~(layer_6[389] ^ layer_6[374]); 
    assign out[386] = ~layer_6[383]; 
    assign out[387] = ~(layer_6[373] | layer_6[391]); 
    assign out[388] = layer_6[393] & ~layer_6[391]; 
    assign out[389] = layer_6[385] | layer_6[385]; 
    assign out[390] = layer_6[398] ^ layer_6[404]; 
    assign out[391] = ~(layer_6[402] ^ layer_6[377]); 
    assign out[392] = ~(layer_6[408] & layer_6[388]); 
    assign out[393] = layer_6[377] ^ layer_6[407]; 
    assign out[394] = ~layer_6[385]; 
    assign out[395] = ~(layer_6[402] & layer_6[381]); 
    assign out[396] = layer_6[407]; 
    assign out[397] = ~layer_6[394] | (layer_6[391] & layer_6[394]); 
    assign out[398] = ~(layer_6[393] ^ layer_6[385]); 
    assign out[399] = 1'b0; 
    assign out[400] = ~(layer_6[398] ^ layer_6[389]); 
    assign out[401] = ~layer_6[389] | (layer_6[389] & layer_6[389]); 
    assign out[402] = layer_6[391] & ~layer_6[414]; 
    assign out[403] = layer_6[405] & ~layer_6[410]; 
    assign out[404] = ~layer_6[406] | (layer_6[397] & layer_6[406]); 
    assign out[405] = ~(layer_6[416] ^ layer_6[420]); 
    assign out[406] = ~layer_6[415] | (layer_6[411] & layer_6[415]); 
    assign out[407] = layer_6[404] & ~layer_6[405]; 
    assign out[408] = ~(layer_6[423] ^ layer_6[414]); 
    assign out[409] = layer_6[417] & layer_6[412]; 
    assign out[410] = layer_6[425] | layer_6[396]; 
    assign out[411] = 1'b1; 
    assign out[412] = ~layer_6[412] | (layer_6[406] & layer_6[412]); 
    assign out[413] = layer_6[403] & ~layer_6[408]; 
    assign out[414] = ~layer_6[400]; 
    assign out[415] = layer_6[416] & layer_6[411]; 
    assign out[416] = layer_6[418] & layer_6[416]; 
    assign out[417] = 1'b1; 
    assign out[418] = layer_6[419] ^ layer_6[401]; 
    assign out[419] = ~(layer_6[417] & layer_6[433]); 
    assign out[420] = ~(layer_6[413] ^ layer_6[403]); 
    assign out[421] = ~layer_6[418]; 
    assign out[422] = layer_6[431] & ~layer_6[415]; 
    assign out[423] = ~layer_6[416]; 
    assign out[424] = layer_6[421] & layer_6[420]; 
    assign out[425] = ~layer_6[420] | (layer_6[413] & layer_6[420]); 
    assign out[426] = ~(layer_6[441] | layer_6[435]); 
    assign out[427] = ~layer_6[416] | (layer_6[416] & layer_6[416]); 
    assign out[428] = ~layer_6[423] | (layer_6[423] & layer_6[440]); 
    assign out[429] = layer_6[429] & ~layer_6[438]; 
    assign out[430] = 1'b0; 
    assign out[431] = layer_6[439] | layer_6[431]; 
    assign out[432] = ~layer_6[431]; 
    assign out[433] = ~layer_6[439] | (layer_6[439] & layer_6[424]); 
    assign out[434] = ~(layer_6[441] ^ layer_6[420]); 
    assign out[435] = ~layer_6[426]; 
    assign out[436] = layer_6[428]; 
    assign out[437] = 1'b0; 
    assign out[438] = layer_6[426] | layer_6[437]; 
    assign out[439] = ~(layer_6[443] & layer_6[449]); 
    assign out[440] = layer_6[448] ^ layer_6[433]; 
    assign out[441] = ~layer_6[454]; 
    assign out[442] = layer_6[432] | layer_6[457]; 
    assign out[443] = layer_6[429] ^ layer_6[441]; 
    assign out[444] = layer_6[436] & layer_6[459]; 
    assign out[445] = 1'b0; 
    assign out[446] = ~layer_6[457]; 
    assign out[447] = 1'b0; 
    assign out[448] = ~layer_6[433] | (layer_6[433] & layer_6[451]); 
    assign out[449] = layer_6[433]; 
    assign out[450] = layer_6[456] ^ layer_6[457]; 
    assign out[451] = layer_6[465] ^ layer_6[438]; 
    assign out[452] = layer_6[458] & layer_6[464]; 
    assign out[453] = ~layer_6[457] | (layer_6[457] & layer_6[452]); 
    assign out[454] = layer_6[461] | layer_6[460]; 
    assign out[455] = layer_6[468]; 
    assign out[456] = 1'b0; 
    assign out[457] = ~layer_6[452] | (layer_6[452] & layer_6[442]); 
    assign out[458] = layer_6[452] & ~layer_6[447]; 
    assign out[459] = 1'b1; 
    assign out[460] = layer_6[457] & ~layer_6[472]; 
    assign out[461] = layer_6[452]; 
    assign out[462] = ~layer_6[450]; 
    assign out[463] = ~(layer_6[476] ^ layer_6[467]); 
    assign out[464] = ~layer_6[450]; 
    assign out[465] = ~layer_6[466]; 
    assign out[466] = ~(layer_6[475] | layer_6[479]); 
    assign out[467] = layer_6[459] | layer_6[467]; 
    assign out[468] = ~layer_6[481] | (layer_6[481] & layer_6[477]); 
    assign out[469] = ~layer_6[478]; 
    assign out[470] = ~layer_6[469]; 
    assign out[471] = layer_6[481]; 
    assign out[472] = layer_6[471] & ~layer_6[472]; 
    assign out[473] = layer_6[480]; 
    assign out[474] = layer_6[480] & ~layer_6[462]; 
    assign out[475] = layer_6[473] ^ layer_6[485]; 
    assign out[476] = 1'b0; 
    assign out[477] = ~(layer_6[462] & layer_6[460]); 
    assign out[478] = 1'b1; 
    assign out[479] = layer_6[472] ^ layer_6[486]; 
    assign out[480] = ~layer_6[494] | (layer_6[494] & layer_6[472]); 
    assign out[481] = ~layer_6[480]; 
    assign out[482] = ~(layer_6[475] ^ layer_6[472]); 
    assign out[483] = 1'b0; 
    assign out[484] = ~layer_6[489]; 
    assign out[485] = layer_6[498] ^ layer_6[469]; 
    assign out[486] = ~layer_6[476] | (layer_6[482] & layer_6[476]); 
    assign out[487] = ~(layer_6[490] ^ layer_6[489]); 
    assign out[488] = ~(layer_6[502] ^ layer_6[493]); 
    assign out[489] = ~(layer_6[484] & layer_6[476]); 
    assign out[490] = layer_6[482]; 
    assign out[491] = layer_6[488]; 
    assign out[492] = layer_6[484] & ~layer_6[483]; 
    assign out[493] = ~layer_6[502] | (layer_6[502] & layer_6[479]); 
    assign out[494] = ~layer_6[504]; 
    assign out[495] = ~(layer_6[503] ^ layer_6[501]); 
    assign out[496] = ~layer_6[504] | (layer_6[504] & layer_6[510]); 
    assign out[497] = layer_6[503] & ~layer_6[510]; 
    assign out[498] = layer_6[483] & layer_6[509]; 
    assign out[499] = layer_6[494] & ~layer_6[488]; 
    assign out[500] = ~(layer_6[510] | layer_6[497]); 
    assign out[501] = layer_6[507] & layer_6[488]; 
    assign out[502] = ~layer_6[504] | (layer_6[504] & layer_6[501]); 
    assign out[503] = layer_6[507]; 
    assign out[504] = ~(layer_6[516] & layer_6[491]); 
    assign out[505] = layer_6[514] & ~layer_6[500]; 
    assign out[506] = ~(layer_6[501] | layer_6[515]); 
    assign out[507] = ~layer_6[496]; 
    assign out[508] = layer_6[522]; 
    assign out[509] = ~(layer_6[511] ^ layer_6[520]); 
    assign out[510] = layer_6[506]; 
    assign out[511] = layer_6[497] ^ layer_6[516]; 
    assign out[512] = layer_6[504]; 
    assign out[513] = ~layer_6[507]; 
    assign out[514] = layer_6[518] ^ layer_6[500]; 
    assign out[515] = 1'b1; 
    assign out[516] = layer_6[521]; 
    assign out[517] = layer_6[530] | layer_6[523]; 
    assign out[518] = layer_6[509]; 
    assign out[519] = 1'b0; 
    assign out[520] = layer_6[534] | layer_6[523]; 
    assign out[521] = 1'b0; 
    assign out[522] = ~layer_6[520]; 
    assign out[523] = layer_6[510] & ~layer_6[506]; 
    assign out[524] = layer_6[539] ^ layer_6[537]; 
    assign out[525] = ~(layer_6[537] | layer_6[530]); 
    assign out[526] = layer_6[537] & layer_6[512]; 
    assign out[527] = ~(layer_6[543] & layer_6[513]); 
    assign out[528] = layer_6[535]; 
    assign out[529] = ~(layer_6[542] | layer_6[524]); 
    assign out[530] = ~(layer_6[526] | layer_6[532]); 
    assign out[531] = layer_6[528] & ~layer_6[531]; 
    assign out[532] = layer_6[541] & ~layer_6[533]; 
    assign out[533] = layer_6[548] ^ layer_6[527]; 
    assign out[534] = ~layer_6[540]; 
    assign out[535] = ~(layer_6[543] ^ layer_6[534]); 
    assign out[536] = layer_6[527]; 
    assign out[537] = 1'b0; 
    assign out[538] = ~layer_6[552] | (layer_6[527] & layer_6[552]); 
    assign out[539] = ~layer_6[529] | (layer_6[529] & layer_6[537]); 
    assign out[540] = layer_6[540]; 
    assign out[541] = ~(layer_6[552] | layer_6[528]); 
    assign out[542] = ~layer_6[536] | (layer_6[536] & layer_6[527]); 
    assign out[543] = layer_6[531] | layer_6[553]; 
    assign out[544] = 1'b0; 
    assign out[545] = ~(layer_6[543] | layer_6[532]); 
    assign out[546] = layer_6[534] | layer_6[544]; 
    assign out[547] = ~(layer_6[537] | layer_6[558]); 
    assign out[548] = ~(layer_6[557] & layer_6[552]); 
    assign out[549] = ~(layer_6[555] & layer_6[538]); 
    assign out[550] = layer_6[541] | layer_6[547]; 
    assign out[551] = layer_6[551] & ~layer_6[546]; 
    assign out[552] = ~layer_6[564] | (layer_6[564] & layer_6[553]); 
    assign out[553] = layer_6[557] | layer_6[537]; 
    assign out[554] = ~layer_6[554]; 
    assign out[555] = layer_6[550]; 
    assign out[556] = layer_6[562]; 
    assign out[557] = ~layer_6[560] | (layer_6[559] & layer_6[560]); 
    assign out[558] = layer_6[562]; 
    assign out[559] = layer_6[543] & ~layer_6[542]; 
    assign out[560] = ~(layer_6[560] ^ layer_6[547]); 
    assign out[561] = layer_6[570] & ~layer_6[573]; 
    assign out[562] = layer_6[575] ^ layer_6[548]; 
    assign out[563] = layer_6[562] | layer_6[551]; 
    assign out[564] = layer_6[566]; 
    assign out[565] = layer_6[567] | layer_6[571]; 
    assign out[566] = layer_6[560] & layer_6[576]; 
    assign out[567] = layer_6[555] ^ layer_6[579]; 
    assign out[568] = ~(layer_6[553] & layer_6[574]); 
    assign out[569] = ~layer_6[560] | (layer_6[566] & layer_6[560]); 
    assign out[570] = layer_6[586]; 
    assign out[571] = layer_6[559]; 
    assign out[572] = ~(layer_6[567] | layer_6[572]); 
    assign out[573] = 1'b1; 
    assign out[574] = layer_6[579] | layer_6[574]; 
    assign out[575] = ~layer_6[578] | (layer_6[578] & layer_6[562]); 
    assign out[576] = layer_6[583] ^ layer_6[568]; 
    assign out[577] = ~layer_6[568]; 
    assign out[578] = layer_6[590]; 
    assign out[579] = layer_6[583] & ~layer_6[592]; 
    assign out[580] = layer_6[574] | layer_6[569]; 
    assign out[581] = ~(layer_6[570] ^ layer_6[581]); 
    assign out[582] = layer_6[583]; 
    assign out[583] = layer_6[567] & ~layer_6[595]; 
    assign out[584] = layer_6[584]; 
    assign out[585] = ~(layer_6[586] & layer_6[575]); 
    assign out[586] = layer_6[573] | layer_6[596]; 
    assign out[587] = ~(layer_6[598] & layer_6[591]); 
    assign out[588] = ~(layer_6[573] ^ layer_6[583]); 
    assign out[589] = ~layer_6[584] | (layer_6[604] & layer_6[584]); 
    assign out[590] = ~layer_6[581] | (layer_6[590] & layer_6[581]); 
    assign out[591] = layer_6[605] & layer_6[599]; 
    assign out[592] = ~(layer_6[591] ^ layer_6[576]); 
    assign out[593] = layer_6[579] ^ layer_6[594]; 
    assign out[594] = layer_6[593]; 
    assign out[595] = layer_6[594]; 
    assign out[596] = ~(layer_6[592] & layer_6[595]); 
    assign out[597] = layer_6[611] | layer_6[586]; 
    assign out[598] = layer_6[597] & ~layer_6[588]; 
    assign out[599] = 1'b1; 
    assign out[600] = layer_6[612] & ~layer_6[605]; 
    assign out[601] = layer_6[594] & ~layer_6[599]; 
    assign out[602] = ~(layer_6[612] ^ layer_6[592]); 
    assign out[603] = ~layer_6[617]; 
    assign out[604] = ~(layer_6[590] ^ layer_6[606]); 
    assign out[605] = ~layer_6[603] | (layer_6[610] & layer_6[603]); 
    assign out[606] = ~layer_6[609]; 
    assign out[607] = layer_6[598] | layer_6[592]; 
    assign out[608] = ~layer_6[595]; 
    assign out[609] = ~layer_6[622]; 
    assign out[610] = 1'b1; 
    assign out[611] = layer_6[616] | layer_6[621]; 
    assign out[612] = 1'b1; 
    assign out[613] = layer_6[625] & ~layer_6[600]; 
    assign out[614] = ~layer_6[619] | (layer_6[615] & layer_6[619]); 
    assign out[615] = ~layer_6[611] | (layer_6[607] & layer_6[611]); 
    assign out[616] = layer_6[625] | layer_6[611]; 
    assign out[617] = layer_6[607] | layer_6[610]; 
    assign out[618] = ~(layer_6[617] ^ layer_6[625]); 
    assign out[619] = ~layer_6[632] | (layer_6[632] & layer_6[611]); 
    assign out[620] = 1'b0; 
    assign out[621] = ~layer_6[613] | (layer_6[613] & layer_6[604]); 
    assign out[622] = ~layer_6[632]; 
    assign out[623] = ~layer_6[633] | (layer_6[627] & layer_6[633]); 
    assign out[624] = ~(layer_6[640] | layer_6[622]); 
    assign out[625] = 1'b0; 
    assign out[626] = layer_6[629] & layer_6[631]; 
    assign out[627] = ~(layer_6[611] & layer_6[612]); 
    assign out[628] = layer_6[624] ^ layer_6[637]; 
    assign out[629] = layer_6[642] ^ layer_6[621]; 
    assign out[630] = ~(layer_6[638] ^ layer_6[632]); 
    assign out[631] = ~(layer_6[639] | layer_6[615]); 
    assign out[632] = layer_6[642] & ~layer_6[622]; 
    assign out[633] = ~(layer_6[646] & layer_6[637]); 
    assign out[634] = layer_6[620] & ~layer_6[624]; 
    assign out[635] = ~layer_6[647] | (layer_6[620] & layer_6[647]); 
    assign out[636] = ~(layer_6[624] ^ layer_6[637]); 
    assign out[637] = 1'b0; 
    assign out[638] = layer_6[639] & ~layer_6[644]; 
    assign out[639] = 1'b0; 
    assign out[640] = layer_6[635]; 
    assign out[641] = ~layer_6[645] | (layer_6[645] & layer_6[627]); 
    assign out[642] = ~layer_6[655] | (layer_6[655] & layer_6[631]); 
    assign out[643] = ~layer_6[655]; 
    assign out[644] = 1'b1; 
    assign out[645] = ~layer_6[648]; 
    assign out[646] = layer_6[654] & ~layer_6[658]; 
    assign out[647] = layer_6[651]; 
    assign out[648] = ~layer_6[636] | (layer_6[636] & layer_6[663]); 
    assign out[649] = 1'b1; 
    assign out[650] = ~layer_6[658] | (layer_6[658] & layer_6[635]); 
    assign out[651] = ~(layer_6[654] | layer_6[639]); 
    assign out[652] = layer_6[646] | layer_6[648]; 
    assign out[653] = ~layer_6[649] | (layer_6[663] & layer_6[649]); 
    assign out[654] = layer_6[667]; 
    assign out[655] = layer_6[664] | layer_6[640]; 
    assign out[656] = layer_6[661] & ~layer_6[649]; 
    assign out[657] = ~(layer_6[649] ^ layer_6[653]); 
    assign out[658] = layer_6[651] | layer_6[643]; 
    assign out[659] = layer_6[655] | layer_6[663]; 
    assign out[660] = 1'b0; 
    assign out[661] = ~(layer_6[652] ^ layer_6[671]); 
    assign out[662] = ~layer_6[645] | (layer_6[647] & layer_6[645]); 
    assign out[663] = layer_6[660] & ~layer_6[656]; 
    assign out[664] = layer_6[671] ^ layer_6[651]; 
    assign out[665] = ~layer_6[659]; 
    assign out[666] = layer_6[664] & ~layer_6[661]; 
    assign out[667] = ~(layer_6[681] & layer_6[671]); 
    assign out[668] = layer_6[652] | layer_6[661]; 
    assign out[669] = 1'b0; 
    assign out[670] = ~layer_6[674] | (layer_6[678] & layer_6[674]); 
    assign out[671] = layer_6[657] & ~layer_6[655]; 
    assign out[672] = layer_6[666] ^ layer_6[687]; 
    assign out[673] = ~(layer_6[688] | layer_6[668]); 
    assign out[674] = ~(layer_6[660] ^ layer_6[674]); 
    assign out[675] = layer_6[667] & ~layer_6[660]; 
    assign out[676] = layer_6[659] & ~layer_6[661]; 
    assign out[677] = layer_6[660] & ~layer_6[690]; 
    assign out[678] = ~layer_6[661]; 
    assign out[679] = ~(layer_6[681] ^ layer_6[676]); 
    assign out[680] = ~layer_6[667] | (layer_6[667] & layer_6[667]); 
    assign out[681] = layer_6[688] | layer_6[681]; 
    assign out[682] = layer_6[685] & ~layer_6[688]; 
    assign out[683] = layer_6[686]; 
    assign out[684] = 1'b0; 
    assign out[685] = layer_6[675] & layer_6[670]; 
    assign out[686] = layer_6[696] & ~layer_6[684]; 
    assign out[687] = ~(layer_6[677] & layer_6[677]); 
    assign out[688] = ~(layer_6[704] ^ layer_6[695]); 
    assign out[689] = ~(layer_6[696] | layer_6[684]); 
    assign out[690] = layer_6[706] & layer_6[700]; 
    assign out[691] = layer_6[696]; 
    assign out[692] = layer_6[690] ^ layer_6[685]; 
    assign out[693] = ~(layer_6[692] & layer_6[677]); 
    assign out[694] = layer_6[680] | layer_6[703]; 
    assign out[695] = layer_6[704]; 
    assign out[696] = layer_6[699]; 
    assign out[697] = ~(layer_6[706] ^ layer_6[683]); 
    assign out[698] = layer_6[699] & ~layer_6[706]; 
    assign out[699] = layer_6[688] & layer_6[687]; 
    assign out[700] = ~layer_6[684] | (layer_6[690] & layer_6[684]); 
    assign out[701] = layer_6[715]; 
    assign out[702] = layer_6[710] | layer_6[698]; 
    assign out[703] = ~layer_6[708]; 
    assign out[704] = layer_6[690] & ~layer_6[718]; 
    assign out[705] = layer_6[691] & layer_6[706]; 
    assign out[706] = ~(layer_6[721] ^ layer_6[720]); 
    assign out[707] = ~(layer_6[697] ^ layer_6[714]); 
    assign out[708] = layer_6[706]; 
    assign out[709] = layer_6[695] & layer_6[700]; 
    assign out[710] = 1'b1; 
    assign out[711] = layer_6[697] ^ layer_6[705]; 
    assign out[712] = ~layer_6[695]; 
    assign out[713] = ~(layer_6[707] ^ layer_6[717]); 
    assign out[714] = ~(layer_6[705] ^ layer_6[728]); 
    assign out[715] = layer_6[708] & ~layer_6[725]; 
    assign out[716] = ~layer_6[726] | (layer_6[715] & layer_6[726]); 
    assign out[717] = layer_6[711] ^ layer_6[721]; 
    assign out[718] = layer_6[709] & ~layer_6[712]; 
    assign out[719] = ~(layer_6[713] ^ layer_6[717]); 
    assign out[720] = layer_6[711] ^ layer_6[733]; 
    assign out[721] = ~(layer_6[729] | layer_6[731]); 
    assign out[722] = 1'b1; 
    assign out[723] = layer_6[718]; 
    assign out[724] = layer_6[718] | layer_6[733]; 
    assign out[725] = ~(layer_6[730] | layer_6[720]); 
    assign out[726] = ~(layer_6[739] & layer_6[726]); 
    assign out[727] = 1'b0; 
    assign out[728] = layer_6[726] & layer_6[712]; 
    assign out[729] = layer_6[741] & ~layer_6[723]; 
    assign out[730] = layer_6[726] ^ layer_6[718]; 
    assign out[731] = layer_6[743] ^ layer_6[728]; 
    assign out[732] = layer_6[735] ^ layer_6[747]; 
    assign out[733] = ~(layer_6[739] | layer_6[742]); 
    assign out[734] = layer_6[739]; 
    assign out[735] = layer_6[736] | layer_6[742]; 
    assign out[736] = layer_6[737] & ~layer_6[720]; 
    assign out[737] = ~(layer_6[731] ^ layer_6[728]); 
    assign out[738] = layer_6[732] & ~layer_6[752]; 
    assign out[739] = layer_6[752] & layer_6[752]; 
    assign out[740] = ~(layer_6[749] | layer_6[743]); 
    assign out[741] = 1'b0; 
    assign out[742] = 1'b0; 
    assign out[743] = layer_6[759] & layer_6[735]; 
    assign out[744] = ~layer_6[743] | (layer_6[728] & layer_6[743]); 
    assign out[745] = layer_6[743] & layer_6[752]; 
    assign out[746] = ~(layer_6[751] & layer_6[736]); 
    assign out[747] = ~layer_6[734]; 
    assign out[748] = layer_6[759] & layer_6[753]; 
    assign out[749] = layer_6[746] & layer_6[748]; 
    assign out[750] = layer_6[760] | layer_6[741]; 
    assign out[751] = layer_6[766] & ~layer_6[755]; 
    assign out[752] = layer_6[749] & layer_6[757]; 
    assign out[753] = layer_6[764] | layer_6[736]; 
    assign out[754] = layer_6[740]; 
    assign out[755] = layer_6[770]; 
    assign out[756] = ~(layer_6[767] ^ layer_6[744]); 
    assign out[757] = ~(layer_6[771] & layer_6[740]); 
    assign out[758] = ~layer_6[758]; 
    assign out[759] = layer_6[758] | layer_6[766]; 
    assign out[760] = ~(layer_6[745] & layer_6[767]); 
    assign out[761] = 1'b0; 
    assign out[762] = ~(layer_6[766] ^ layer_6[750]); 
    assign out[763] = 1'b1; 
    assign out[764] = 1'b0; 
    assign out[765] = ~(layer_6[754] & layer_6[750]); 
    assign out[766] = ~layer_6[761] | (layer_6[761] & layer_6[764]); 
    assign out[767] = layer_6[768] | layer_6[758]; 
    assign out[768] = layer_6[758]; 
    assign out[769] = layer_6[766] & ~layer_6[763]; 
    assign out[770] = layer_6[774]; 
    assign out[771] = ~(layer_6[760] ^ layer_6[782]); 
    assign out[772] = 1'b0; 
    assign out[773] = ~(layer_6[780] ^ layer_6[760]); 
    assign out[774] = layer_6[771]; 
    assign out[775] = layer_6[776] & ~layer_6[779]; 
    assign out[776] = layer_6[788] & ~layer_6[789]; 
    assign out[777] = ~(layer_6[788] & layer_6[760]); 
    assign out[778] = layer_6[775] | layer_6[778]; 
    assign out[779] = layer_6[781] & ~layer_6[766]; 
    assign out[780] = 1'b1; 
    assign out[781] = ~(layer_6[771] ^ layer_6[772]); 
    assign out[782] = layer_6[780] & ~layer_6[798]; 
    assign out[783] = ~layer_6[794]; 
    assign out[784] = layer_6[779] & ~layer_6[773]; 
    assign out[785] = ~(layer_6[797] | layer_6[780]); 
    assign out[786] = layer_6[792]; 
    assign out[787] = layer_6[782] | layer_6[780]; 
    assign out[788] = 1'b0; 
    assign out[789] = ~layer_6[797] | (layer_6[797] & layer_6[791]); 
    assign out[790] = 1'b1; 
    assign out[791] = 1'b0; 
    assign out[792] = 1'b0; 
    assign out[793] = layer_6[808] ^ layer_6[789]; 
    assign out[794] = 1'b1; 
    assign out[795] = layer_6[782]; 
    assign out[796] = 1'b0; 
    assign out[797] = layer_6[810] | layer_6[811]; 
    assign out[798] = layer_6[787]; 
    assign out[799] = layer_6[810] & ~layer_6[814]; 
    assign out[800] = layer_6[788] & ~layer_6[814]; 
    assign out[801] = ~(layer_6[804] | layer_6[800]); 
    assign out[802] = ~(layer_6[802] & layer_6[817]); 
    assign out[803] = layer_6[789] | layer_6[788]; 
    assign out[804] = 1'b1; 
    assign out[805] = ~layer_6[818] | (layer_6[818] & layer_6[807]); 
    assign out[806] = layer_6[817] ^ layer_6[818]; 
    assign out[807] = layer_6[797] | layer_6[795]; 
    assign out[808] = 1'b0; 
    assign out[809] = layer_6[820] ^ layer_6[810]; 
    assign out[810] = ~(layer_6[823] | layer_6[814]); 
    assign out[811] = 1'b0; 
    assign out[812] = 1'b1; 
    assign out[813] = ~(layer_6[800] | layer_6[827]); 
    assign out[814] = layer_6[814]; 
    assign out[815] = layer_6[828] & layer_6[824]; 
    assign out[816] = layer_6[805]; 
    assign out[817] = layer_6[830] & layer_6[829]; 
    assign out[818] = ~layer_6[802] | (layer_6[802] & layer_6[832]); 
    assign out[819] = ~layer_6[834]; 
    assign out[820] = ~layer_6[823]; 
    assign out[821] = layer_6[809] ^ layer_6[822]; 
    assign out[822] = ~(layer_6[831] ^ layer_6[817]); 
    assign out[823] = layer_6[813] & layer_6[807]; 
    assign out[824] = layer_6[807] & ~layer_6[838]; 
    assign out[825] = 1'b0; 
    assign out[826] = 1'b0; 
    assign out[827] = layer_6[812] | layer_6[831]; 
    assign out[828] = ~(layer_6[843] | layer_6[812]); 
    assign out[829] = 1'b0; 
    assign out[830] = layer_6[821] ^ layer_6[818]; 
    assign out[831] = ~layer_6[823] | (layer_6[823] & layer_6[837]); 
    assign out[832] = layer_6[837] | layer_6[820]; 
    assign out[833] = ~(layer_6[841] | layer_6[825]); 
    assign out[834] = 1'b1; 
    assign out[835] = layer_6[849] & ~layer_6[832]; 
    assign out[836] = ~layer_6[849] | (layer_6[849] & layer_6[832]); 
    assign out[837] = layer_6[837] & ~layer_6[829]; 
    assign out[838] = ~layer_6[848] | (layer_6[848] & layer_6[827]); 
    assign out[839] = ~(layer_6[836] | layer_6[852]); 
    assign out[840] = layer_6[843] | layer_6[841]; 
    assign out[841] = layer_6[833] & ~layer_6[830]; 
    assign out[842] = layer_6[831] & layer_6[844]; 
    assign out[843] = layer_6[830] & ~layer_6[836]; 
    assign out[844] = layer_6[860] ^ layer_6[850]; 
    assign out[845] = 1'b1; 
    assign out[846] = layer_6[851] ^ layer_6[857]; 
    assign out[847] = layer_6[837]; 
    assign out[848] = 1'b1; 
    assign out[849] = layer_6[841] & ~layer_6[854]; 
    assign out[850] = layer_6[853] & ~layer_6[857]; 
    assign out[851] = ~layer_6[848] | (layer_6[860] & layer_6[848]); 
    assign out[852] = 1'b0; 
    assign out[853] = ~(layer_6[863] | layer_6[857]); 
    assign out[854] = ~layer_6[855]; 
    assign out[855] = layer_6[865]; 
    assign out[856] = ~layer_6[852] | (layer_6[852] & layer_6[844]); 
    assign out[857] = layer_6[842]; 
    assign out[858] = ~layer_6[871]; 
    assign out[859] = ~(layer_6[843] ^ layer_6[869]); 
    assign out[860] = ~layer_6[853]; 
    assign out[861] = layer_6[864] ^ layer_6[847]; 
    assign out[862] = ~(layer_6[861] | layer_6[857]); 
    assign out[863] = 1'b1; 
    assign out[864] = 1'b0; 
    assign out[865] = layer_6[877] & layer_6[867]; 
    assign out[866] = ~(layer_6[866] & layer_6[859]); 
    assign out[867] = layer_6[865] & layer_6[874]; 
    assign out[868] = ~layer_6[858] | (layer_6[858] & layer_6[865]); 
    assign out[869] = layer_6[880] ^ layer_6[869]; 
    assign out[870] = layer_6[859] & ~layer_6[871]; 
    assign out[871] = layer_6[873]; 
    assign out[872] = layer_6[877]; 
    assign out[873] = ~(layer_6[882] | layer_6[865]); 
    assign out[874] = layer_6[876]; 
    assign out[875] = layer_6[862] & layer_6[871]; 
    assign out[876] = layer_6[875] ^ layer_6[875]; 
    assign out[877] = ~(layer_6[888] ^ layer_6[873]); 
    assign out[878] = layer_6[875] & ~layer_6[877]; 
    assign out[879] = ~layer_6[876] | (layer_6[876] & layer_6[870]); 
    assign out[880] = layer_6[867] | layer_6[863]; 
    assign out[881] = layer_6[887] & layer_6[865]; 
    assign out[882] = ~layer_6[868] | (layer_6[888] & layer_6[868]); 
    assign out[883] = ~(layer_6[884] | layer_6[885]); 
    assign out[884] = layer_6[896]; 
    assign out[885] = layer_6[887] & ~layer_6[877]; 
    assign out[886] = ~layer_6[876]; 
    assign out[887] = ~(layer_6[881] & layer_6[895]); 
    assign out[888] = ~layer_6[890]; 
    assign out[889] = layer_6[879]; 
    assign out[890] = layer_6[880]; 
    assign out[891] = ~layer_6[894]; 
    assign out[892] = layer_6[881]; 
    assign out[893] = layer_6[884] & ~layer_6[896]; 
    assign out[894] = 1'b1; 
    assign out[895] = layer_6[890] & ~layer_6[881]; 
    assign out[896] = 1'b1; 
    assign out[897] = layer_6[882] | layer_6[897]; 
    assign out[898] = ~(layer_6[884] ^ layer_6[884]); 
    assign out[899] = ~(layer_6[884] ^ layer_6[902]); 
    assign out[900] = layer_6[889]; 
    assign out[901] = layer_6[916] & ~layer_6[901]; 
    assign out[902] = layer_6[895] & ~layer_6[913]; 
    assign out[903] = ~layer_6[912]; 
    assign out[904] = layer_6[893]; 
    assign out[905] = ~(layer_6[910] | layer_6[904]); 
    assign out[906] = layer_6[894] ^ layer_6[898]; 
    assign out[907] = layer_6[911]; 
    assign out[908] = 1'b1; 
    assign out[909] = layer_6[922] & ~layer_6[918]; 
    assign out[910] = 1'b0; 
    assign out[911] = ~(layer_6[924] ^ layer_6[914]); 
    assign out[912] = layer_6[919] & ~layer_6[923]; 
    assign out[913] = layer_6[898]; 
    assign out[914] = 1'b1; 
    assign out[915] = layer_6[904] ^ layer_6[910]; 
    assign out[916] = ~layer_6[923]; 
    assign out[917] = layer_6[914] & ~layer_6[902]; 
    assign out[918] = layer_6[914] | layer_6[925]; 
    assign out[919] = ~layer_6[903]; 
    assign out[920] = layer_6[921] & layer_6[919]; 
    assign out[921] = 1'b1; 
    assign out[922] = layer_6[929] | layer_6[920]; 
    assign out[923] = layer_6[909] ^ layer_6[933]; 
    assign out[924] = 1'b1; 
    assign out[925] = ~layer_6[926]; 
    assign out[926] = ~layer_6[919] | (layer_6[919] & layer_6[932]); 
    assign out[927] = layer_6[911] & layer_6[934]; 
    assign out[928] = layer_6[927] | layer_6[940]; 
    assign out[929] = ~(layer_6[913] | layer_6[929]); 
    assign out[930] = ~layer_6[940] | (layer_6[943] & layer_6[940]); 
    assign out[931] = ~(layer_6[939] & layer_6[920]); 
    assign out[932] = layer_6[930]; 
    assign out[933] = layer_6[931] ^ layer_6[918]; 
    assign out[934] = 1'b1; 
    assign out[935] = layer_6[935] & layer_6[927]; 
    assign out[936] = layer_6[949] & ~layer_6[926]; 
    assign out[937] = ~(layer_6[944] ^ layer_6[951]); 
    assign out[938] = layer_6[943] ^ layer_6[945]; 
    assign out[939] = layer_6[950] | layer_6[925]; 
    assign out[940] = ~layer_6[950]; 
    assign out[941] = layer_6[927] ^ layer_6[924]; 
    assign out[942] = layer_6[957] ^ layer_6[945]; 
    assign out[943] = ~layer_6[939]; 
    assign out[944] = ~layer_6[958] | (layer_6[958] & layer_6[956]); 
    assign out[945] = layer_6[948] & ~layer_6[928]; 
    assign out[946] = ~layer_6[962]; 
    assign out[947] = layer_6[946] & ~layer_6[937]; 
    assign out[948] = layer_6[932]; 
    assign out[949] = ~layer_6[949] | (layer_6[951] & layer_6[949]); 
    assign out[950] = layer_6[933] & ~layer_6[956]; 
    assign out[951] = 1'b1; 
    assign out[952] = layer_6[943]; 
    assign out[953] = ~layer_6[948] | (layer_6[948] & layer_6[939]); 
    assign out[954] = layer_6[964] ^ layer_6[966]; 
    assign out[955] = 1'b1; 
    assign out[956] = ~(layer_6[971] | layer_6[946]); 
    assign out[957] = layer_6[958]; 
    assign out[958] = ~layer_6[966] | (layer_6[966] & layer_6[971]); 
    assign out[959] = ~layer_6[966] | (layer_6[973] & layer_6[966]); 
    assign out[960] = ~(layer_6[970] ^ layer_6[974]); 
    assign out[961] = ~layer_6[965] | (layer_6[965] & layer_6[966]); 
    assign out[962] = ~(layer_6[963] ^ layer_6[969]); 
    assign out[963] = 1'b0; 
    assign out[964] = layer_6[956] | layer_6[958]; 
    assign out[965] = layer_6[951] ^ layer_6[960]; 
    assign out[966] = layer_6[967] | layer_6[955]; 
    assign out[967] = 1'b1; 
    assign out[968] = ~(layer_6[971] & layer_6[976]); 
    assign out[969] = ~layer_6[971]; 
    assign out[970] = layer_6[983] & ~layer_6[958]; 
    assign out[971] = layer_6[964] & ~layer_6[959]; 
    assign out[972] = ~(layer_6[983] | layer_6[968]); 
    assign out[973] = layer_6[958] ^ layer_6[960]; 
    assign out[974] = ~layer_6[970]; 
    assign out[975] = ~(layer_6[975] ^ layer_6[970]); 
    assign out[976] = ~layer_6[963] | (layer_6[963] & layer_6[981]); 
    assign out[977] = ~(layer_6[975] ^ layer_6[990]); 
    assign out[978] = layer_6[984] ^ layer_6[962]; 
    assign out[979] = layer_6[971] | layer_6[983]; 
    assign out[980] = layer_6[993] & ~layer_6[973]; 
    assign out[981] = ~layer_6[993]; 
    assign out[982] = layer_6[982] ^ layer_6[973]; 
    assign out[983] = ~(layer_6[988] | layer_6[995]); 
    assign out[984] = ~(layer_6[1000] & layer_6[974]); 
    assign out[985] = layer_6[971] ^ layer_6[972]; 
    assign out[986] = layer_6[1000] & layer_6[977]; 
    assign out[987] = 1'b0; 
    assign out[988] = ~(layer_6[994] ^ layer_6[997]); 
    assign out[989] = layer_6[980] | layer_6[1004]; 
    assign out[990] = layer_6[988]; 
    assign out[991] = layer_6[988] ^ layer_6[1001]; 
    assign out[992] = layer_6[998] & layer_6[1004]; 
    assign out[993] = layer_6[981]; 
    assign out[994] = ~layer_6[1000]; 
    assign out[995] = ~(layer_6[996] ^ layer_6[979]); 
    assign out[996] = ~layer_6[1000]; 
    assign out[997] = ~(layer_6[983] & layer_6[1005]); 
    assign out[998] = ~(layer_6[997] & layer_6[997]); 
    assign out[999] = layer_6[1010]; 
    assign out[1000] = layer_6[999]; 
    assign out[1001] = layer_6[989] | layer_6[1010]; 
    assign out[1002] = ~layer_6[1016]; 
    assign out[1003] = layer_6[995] & ~layer_6[990]; 
    assign out[1004] = ~(layer_6[1009] ^ layer_6[1016]); 
    assign out[1005] = layer_6[1012]; 
    assign out[1006] = layer_6[993] & ~layer_6[1009]; 
    assign out[1007] = ~layer_6[991]; 
    assign out[1008] = ~(layer_6[1022] ^ layer_6[997]); 
    assign out[1009] = layer_6[998]; 
    assign out[1010] = layer_6[1023] | layer_6[1013]; 
    assign out[1011] = layer_6[1021] | layer_6[1021]; 
    assign out[1012] = ~layer_6[1021]; 
    assign out[1013] = ~(layer_6[1014] & layer_6[1008]); 
    assign out[1014] = ~layer_6[1014]; 
    assign out[1015] = layer_6[1005]; 
    assign out[1016] = ~(layer_6[1019] & layer_6[1003]); 
    assign out[1017] = layer_6[1020] & layer_6[1003]; 
    assign out[1018] = layer_6[1009] ^ layer_6[1022]; 
    assign out[1019] = ~(layer_6[1012] ^ layer_6[1015]); 
    assign out[1020] = layer_6[1013]; 
    assign out[1021] = layer_6[1013]; 
    assign out[1022] = ~layer_6[1008]; 
    assign out[1023] = ~layer_6[1017] | (layer_6[1017] & layer_6[1013]); 

endmodule
