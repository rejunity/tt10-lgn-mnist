// Generated from: barabasi_20250115-080837_acc7913_seed176567_epochs100_dispersion128_1020-1020-1020-1020-1020-1020-1020-1020.npz
`ifdef SIM
module sky130_fd_sc_hd__inv_1 (
    input wire A,
    output wire Y
);
    assign Y = ~A;
endmodule
`endif
module relay_conn (
    input wire in,
    output wire out
);
    wire tmp;
    /* verilator lint_off PINMISSING */
    // https://skywater-pdk.readthedocs.io/en/main/contents/libraries/sky130_fd_sc_hd/cells/inv/README.html
    (* keep = "true" *) sky130_fd_sc_hd__inv_1 inv_a ( .Y(tmp), .A(in)  );
    (* keep = "true" *) sky130_fd_sc_hd__inv_1 inv_b ( .Y(out), .A(tmp) );
    /* verilator lint_on PINMISSING */
endmodule 
module net (
    input wire  [255:0] in,
    output wire [1019:0] out
);
    wire [1020:0] layer_0;
    wire [1020:0] layer_1;
    wire [1020:0] layer_2;
    wire [1020:0] layer_3;
    wire [1020:0] layer_4;
    wire [1020:0] layer_5;
    wire [1020:0] layer_6;

    // Layer 0 ============================================================
    wire [1:0] far_0_0_0;    relay_conn far_0_0_0_a(.in(in[99]), .out(far_0_0_0[0]));    relay_conn far_0_0_0_b(.in(in[19]), .out(far_0_0_0[1]));
    wire [1:0] far_0_0_1;    relay_conn far_0_0_1_a(.in(far_0_0_0[0]), .out(far_0_0_1[0]));    relay_conn far_0_0_1_b(.in(far_0_0_0[1]), .out(far_0_0_1[1]));
    assign layer_0[0] = ~far_0_0_1[1]; 
    wire [1:0] far_0_1_0;    relay_conn far_0_1_0_a(.in(in[102]), .out(far_0_1_0[0]));    relay_conn far_0_1_0_b(.in(in[172]), .out(far_0_1_0[1]));
    wire [1:0] far_0_1_1;    relay_conn far_0_1_1_a(.in(far_0_1_0[0]), .out(far_0_1_1[0]));    relay_conn far_0_1_1_b(.in(far_0_1_0[1]), .out(far_0_1_1[1]));
    assign layer_0[1] = far_0_1_1[1] & ~far_0_1_1[0]; 
    assign layer_0[2] = in[22] ^ in[15]; 
    wire [1:0] far_0_3_0;    relay_conn far_0_3_0_a(.in(in[148]), .out(far_0_3_0[0]));    relay_conn far_0_3_0_b(.in(in[240]), .out(far_0_3_0[1]));
    wire [1:0] far_0_3_1;    relay_conn far_0_3_1_a(.in(far_0_3_0[0]), .out(far_0_3_1[0]));    relay_conn far_0_3_1_b(.in(far_0_3_0[1]), .out(far_0_3_1[1]));
    assign layer_0[3] = far_0_3_1[0] & far_0_3_1[1]; 
    wire [1:0] far_0_4_0;    relay_conn far_0_4_0_a(.in(in[157]), .out(far_0_4_0[0]));    relay_conn far_0_4_0_b(.in(in[117]), .out(far_0_4_0[1]));
    assign layer_0[4] = far_0_4_0[0] & ~far_0_4_0[1]; 
    assign layer_0[5] = ~in[211] | (in[211] & in[201]); 
    wire [1:0] far_0_6_0;    relay_conn far_0_6_0_a(.in(in[175]), .out(far_0_6_0[0]));    relay_conn far_0_6_0_b(.in(in[239]), .out(far_0_6_0[1]));
    wire [1:0] far_0_6_1;    relay_conn far_0_6_1_a(.in(far_0_6_0[0]), .out(far_0_6_1[0]));    relay_conn far_0_6_1_b(.in(far_0_6_0[1]), .out(far_0_6_1[1]));
    assign layer_0[6] = ~far_0_6_1[1] | (far_0_6_1[0] & far_0_6_1[1]); 
    assign layer_0[7] = ~in[175]; 
    wire [1:0] far_0_8_0;    relay_conn far_0_8_0_a(.in(in[173]), .out(far_0_8_0[0]));    relay_conn far_0_8_0_b(.in(in[215]), .out(far_0_8_0[1]));
    assign layer_0[8] = ~far_0_8_0[1] | (far_0_8_0[0] & far_0_8_0[1]); 
    assign layer_0[9] = ~in[211] | (in[211] & in[225]); 
    wire [1:0] far_0_10_0;    relay_conn far_0_10_0_a(.in(in[188]), .out(far_0_10_0[0]));    relay_conn far_0_10_0_b(.in(in[109]), .out(far_0_10_0[1]));
    wire [1:0] far_0_10_1;    relay_conn far_0_10_1_a(.in(far_0_10_0[0]), .out(far_0_10_1[0]));    relay_conn far_0_10_1_b(.in(far_0_10_0[1]), .out(far_0_10_1[1]));
    assign layer_0[10] = far_0_10_1[0] & far_0_10_1[1]; 
    wire [1:0] far_0_11_0;    relay_conn far_0_11_0_a(.in(in[177]), .out(far_0_11_0[0]));    relay_conn far_0_11_0_b(.in(in[225]), .out(far_0_11_0[1]));
    assign layer_0[11] = far_0_11_0[0] & far_0_11_0[1]; 
    assign layer_0[12] = ~(in[197] & in[199]); 
    wire [1:0] far_0_13_0;    relay_conn far_0_13_0_a(.in(in[174]), .out(far_0_13_0[0]));    relay_conn far_0_13_0_b(.in(in[99]), .out(far_0_13_0[1]));
    wire [1:0] far_0_13_1;    relay_conn far_0_13_1_a(.in(far_0_13_0[0]), .out(far_0_13_1[0]));    relay_conn far_0_13_1_b(.in(far_0_13_0[1]), .out(far_0_13_1[1]));
    assign layer_0[13] = far_0_13_1[0] & ~far_0_13_1[1]; 
    wire [1:0] far_0_14_0;    relay_conn far_0_14_0_a(.in(in[254]), .out(far_0_14_0[0]));    relay_conn far_0_14_0_b(.in(in[137]), .out(far_0_14_0[1]));
    wire [1:0] far_0_14_1;    relay_conn far_0_14_1_a(.in(far_0_14_0[0]), .out(far_0_14_1[0]));    relay_conn far_0_14_1_b(.in(far_0_14_0[1]), .out(far_0_14_1[1]));
    wire [1:0] far_0_14_2;    relay_conn far_0_14_2_a(.in(far_0_14_1[0]), .out(far_0_14_2[0]));    relay_conn far_0_14_2_b(.in(far_0_14_1[1]), .out(far_0_14_2[1]));
    assign layer_0[14] = far_0_14_2[0]; 
    assign layer_0[15] = ~in[71] | (in[71] & in[59]); 
    assign layer_0[16] = in[157] & ~in[165]; 
    assign layer_0[17] = ~in[221]; 
    wire [1:0] far_0_18_0;    relay_conn far_0_18_0_a(.in(in[88]), .out(far_0_18_0[0]));    relay_conn far_0_18_0_b(.in(in[179]), .out(far_0_18_0[1]));
    wire [1:0] far_0_18_1;    relay_conn far_0_18_1_a(.in(far_0_18_0[0]), .out(far_0_18_1[0]));    relay_conn far_0_18_1_b(.in(far_0_18_0[1]), .out(far_0_18_1[1]));
    assign layer_0[18] = ~far_0_18_1[1]; 
    wire [1:0] far_0_19_0;    relay_conn far_0_19_0_a(.in(in[73]), .out(far_0_19_0[0]));    relay_conn far_0_19_0_b(.in(in[117]), .out(far_0_19_0[1]));
    assign layer_0[19] = far_0_19_0[0] & ~far_0_19_0[1]; 
    wire [1:0] far_0_20_0;    relay_conn far_0_20_0_a(.in(in[186]), .out(far_0_20_0[0]));    relay_conn far_0_20_0_b(.in(in[127]), .out(far_0_20_0[1]));
    assign layer_0[20] = far_0_20_0[1] & ~far_0_20_0[0]; 
    wire [1:0] far_0_21_0;    relay_conn far_0_21_0_a(.in(in[15]), .out(far_0_21_0[0]));    relay_conn far_0_21_0_b(.in(in[82]), .out(far_0_21_0[1]));
    wire [1:0] far_0_21_1;    relay_conn far_0_21_1_a(.in(far_0_21_0[0]), .out(far_0_21_1[0]));    relay_conn far_0_21_1_b(.in(far_0_21_0[1]), .out(far_0_21_1[1]));
    assign layer_0[21] = ~far_0_21_1[0] | (far_0_21_1[0] & far_0_21_1[1]); 
    wire [1:0] far_0_22_0;    relay_conn far_0_22_0_a(.in(in[165]), .out(far_0_22_0[0]));    relay_conn far_0_22_0_b(.in(in[197]), .out(far_0_22_0[1]));
    assign layer_0[22] = ~far_0_22_0[0] | (far_0_22_0[0] & far_0_22_0[1]); 
    wire [1:0] far_0_23_0;    relay_conn far_0_23_0_a(.in(in[176]), .out(far_0_23_0[0]));    relay_conn far_0_23_0_b(.in(in[139]), .out(far_0_23_0[1]));
    assign layer_0[23] = far_0_23_0[0] | far_0_23_0[1]; 
    assign layer_0[24] = in[186] & ~in[191]; 
    wire [1:0] far_0_25_0;    relay_conn far_0_25_0_a(.in(in[113]), .out(far_0_25_0[0]));    relay_conn far_0_25_0_b(.in(in[204]), .out(far_0_25_0[1]));
    wire [1:0] far_0_25_1;    relay_conn far_0_25_1_a(.in(far_0_25_0[0]), .out(far_0_25_1[0]));    relay_conn far_0_25_1_b(.in(far_0_25_0[1]), .out(far_0_25_1[1]));
    assign layer_0[25] = ~far_0_25_1[1] | (far_0_25_1[0] & far_0_25_1[1]); 
    assign layer_0[26] = ~in[160] | (in[186] & in[160]); 
    wire [1:0] far_0_27_0;    relay_conn far_0_27_0_a(.in(in[92]), .out(far_0_27_0[0]));    relay_conn far_0_27_0_b(.in(in[211]), .out(far_0_27_0[1]));
    wire [1:0] far_0_27_1;    relay_conn far_0_27_1_a(.in(far_0_27_0[0]), .out(far_0_27_1[0]));    relay_conn far_0_27_1_b(.in(far_0_27_0[1]), .out(far_0_27_1[1]));
    wire [1:0] far_0_27_2;    relay_conn far_0_27_2_a(.in(far_0_27_1[0]), .out(far_0_27_2[0]));    relay_conn far_0_27_2_b(.in(far_0_27_1[1]), .out(far_0_27_2[1]));
    assign layer_0[27] = far_0_27_2[0]; 
    wire [1:0] far_0_28_0;    relay_conn far_0_28_0_a(.in(in[151]), .out(far_0_28_0[0]));    relay_conn far_0_28_0_b(.in(in[48]), .out(far_0_28_0[1]));
    wire [1:0] far_0_28_1;    relay_conn far_0_28_1_a(.in(far_0_28_0[0]), .out(far_0_28_1[0]));    relay_conn far_0_28_1_b(.in(far_0_28_0[1]), .out(far_0_28_1[1]));
    wire [1:0] far_0_28_2;    relay_conn far_0_28_2_a(.in(far_0_28_1[0]), .out(far_0_28_2[0]));    relay_conn far_0_28_2_b(.in(far_0_28_1[1]), .out(far_0_28_2[1]));
    assign layer_0[28] = far_0_28_2[0] & ~far_0_28_2[1]; 
    assign layer_0[29] = in[199] & ~in[179]; 
    wire [1:0] far_0_30_0;    relay_conn far_0_30_0_a(.in(in[130]), .out(far_0_30_0[0]));    relay_conn far_0_30_0_b(.in(in[5]), .out(far_0_30_0[1]));
    wire [1:0] far_0_30_1;    relay_conn far_0_30_1_a(.in(far_0_30_0[0]), .out(far_0_30_1[0]));    relay_conn far_0_30_1_b(.in(far_0_30_0[1]), .out(far_0_30_1[1]));
    wire [1:0] far_0_30_2;    relay_conn far_0_30_2_a(.in(far_0_30_1[0]), .out(far_0_30_2[0]));    relay_conn far_0_30_2_b(.in(far_0_30_1[1]), .out(far_0_30_2[1]));
    assign layer_0[30] = ~far_0_30_2[1]; 
    wire [1:0] far_0_31_0;    relay_conn far_0_31_0_a(.in(in[221]), .out(far_0_31_0[0]));    relay_conn far_0_31_0_b(.in(in[125]), .out(far_0_31_0[1]));
    wire [1:0] far_0_31_1;    relay_conn far_0_31_1_a(.in(far_0_31_0[0]), .out(far_0_31_1[0]));    relay_conn far_0_31_1_b(.in(far_0_31_0[1]), .out(far_0_31_1[1]));
    wire [1:0] far_0_31_2;    relay_conn far_0_31_2_a(.in(far_0_31_1[0]), .out(far_0_31_2[0]));    relay_conn far_0_31_2_b(.in(far_0_31_1[1]), .out(far_0_31_2[1]));
    assign layer_0[31] = far_0_31_2[0] ^ far_0_31_2[1]; 
    wire [1:0] far_0_32_0;    relay_conn far_0_32_0_a(.in(in[64]), .out(far_0_32_0[0]));    relay_conn far_0_32_0_b(.in(in[101]), .out(far_0_32_0[1]));
    assign layer_0[32] = ~(far_0_32_0[0] ^ far_0_32_0[1]); 
    wire [1:0] far_0_33_0;    relay_conn far_0_33_0_a(.in(in[225]), .out(far_0_33_0[0]));    relay_conn far_0_33_0_b(.in(in[99]), .out(far_0_33_0[1]));
    wire [1:0] far_0_33_1;    relay_conn far_0_33_1_a(.in(far_0_33_0[0]), .out(far_0_33_1[0]));    relay_conn far_0_33_1_b(.in(far_0_33_0[1]), .out(far_0_33_1[1]));
    wire [1:0] far_0_33_2;    relay_conn far_0_33_2_a(.in(far_0_33_1[0]), .out(far_0_33_2[0]));    relay_conn far_0_33_2_b(.in(far_0_33_1[1]), .out(far_0_33_2[1]));
    assign layer_0[33] = ~far_0_33_2[1]; 
    wire [1:0] far_0_34_0;    relay_conn far_0_34_0_a(.in(in[238]), .out(far_0_34_0[0]));    relay_conn far_0_34_0_b(.in(in[151]), .out(far_0_34_0[1]));
    wire [1:0] far_0_34_1;    relay_conn far_0_34_1_a(.in(far_0_34_0[0]), .out(far_0_34_1[0]));    relay_conn far_0_34_1_b(.in(far_0_34_0[1]), .out(far_0_34_1[1]));
    assign layer_0[34] = ~(far_0_34_1[0] | far_0_34_1[1]); 
    assign layer_0[35] = ~in[81]; 
    assign layer_0[36] = in[202]; 
    wire [1:0] far_0_37_0;    relay_conn far_0_37_0_a(.in(in[136]), .out(far_0_37_0[0]));    relay_conn far_0_37_0_b(.in(in[66]), .out(far_0_37_0[1]));
    wire [1:0] far_0_37_1;    relay_conn far_0_37_1_a(.in(far_0_37_0[0]), .out(far_0_37_1[0]));    relay_conn far_0_37_1_b(.in(far_0_37_0[1]), .out(far_0_37_1[1]));
    assign layer_0[37] = far_0_37_1[0] | far_0_37_1[1]; 
    wire [1:0] far_0_38_0;    relay_conn far_0_38_0_a(.in(in[79]), .out(far_0_38_0[0]));    relay_conn far_0_38_0_b(.in(in[17]), .out(far_0_38_0[1]));
    assign layer_0[38] = ~(far_0_38_0[0] | far_0_38_0[1]); 
    assign layer_0[39] = ~in[188] | (in[173] & in[188]); 
    assign layer_0[40] = in[186] & ~in[188]; 
    wire [1:0] far_0_41_0;    relay_conn far_0_41_0_a(.in(in[113]), .out(far_0_41_0[0]));    relay_conn far_0_41_0_b(.in(in[186]), .out(far_0_41_0[1]));
    wire [1:0] far_0_41_1;    relay_conn far_0_41_1_a(.in(far_0_41_0[0]), .out(far_0_41_1[0]));    relay_conn far_0_41_1_b(.in(far_0_41_0[1]), .out(far_0_41_1[1]));
    assign layer_0[41] = far_0_41_1[0] ^ far_0_41_1[1]; 
    assign layer_0[42] = ~in[236] | (in[236] & in[205]); 
    wire [1:0] far_0_43_0;    relay_conn far_0_43_0_a(.in(in[240]), .out(far_0_43_0[0]));    relay_conn far_0_43_0_b(.in(in[202]), .out(far_0_43_0[1]));
    assign layer_0[43] = far_0_43_0[0] & far_0_43_0[1]; 
    wire [1:0] far_0_44_0;    relay_conn far_0_44_0_a(.in(in[38]), .out(far_0_44_0[0]));    relay_conn far_0_44_0_b(.in(in[151]), .out(far_0_44_0[1]));
    wire [1:0] far_0_44_1;    relay_conn far_0_44_1_a(.in(far_0_44_0[0]), .out(far_0_44_1[0]));    relay_conn far_0_44_1_b(.in(far_0_44_0[1]), .out(far_0_44_1[1]));
    wire [1:0] far_0_44_2;    relay_conn far_0_44_2_a(.in(far_0_44_1[0]), .out(far_0_44_2[0]));    relay_conn far_0_44_2_b(.in(far_0_44_1[1]), .out(far_0_44_2[1]));
    assign layer_0[44] = far_0_44_2[1] & ~far_0_44_2[0]; 
    wire [1:0] far_0_45_0;    relay_conn far_0_45_0_a(.in(in[220]), .out(far_0_45_0[0]));    relay_conn far_0_45_0_b(.in(in[164]), .out(far_0_45_0[1]));
    assign layer_0[45] = far_0_45_0[0] & ~far_0_45_0[1]; 
    wire [1:0] far_0_46_0;    relay_conn far_0_46_0_a(.in(in[48]), .out(far_0_46_0[0]));    relay_conn far_0_46_0_b(.in(in[6]), .out(far_0_46_0[1]));
    assign layer_0[46] = ~far_0_46_0[0]; 
    wire [1:0] far_0_47_0;    relay_conn far_0_47_0_a(.in(in[66]), .out(far_0_47_0[0]));    relay_conn far_0_47_0_b(.in(in[113]), .out(far_0_47_0[1]));
    assign layer_0[47] = ~(far_0_47_0[0] & far_0_47_0[1]); 
    assign layer_0[48] = in[98] | in[109]; 
    assign layer_0[49] = in[240] | in[226]; 
    assign layer_0[50] = ~in[165] | (in[134] & in[165]); 
    assign layer_0[51] = in[239] & ~in[219]; 
    wire [1:0] far_0_52_0;    relay_conn far_0_52_0_a(.in(in[133]), .out(far_0_52_0[0]));    relay_conn far_0_52_0_b(.in(in[247]), .out(far_0_52_0[1]));
    wire [1:0] far_0_52_1;    relay_conn far_0_52_1_a(.in(far_0_52_0[0]), .out(far_0_52_1[0]));    relay_conn far_0_52_1_b(.in(far_0_52_0[1]), .out(far_0_52_1[1]));
    wire [1:0] far_0_52_2;    relay_conn far_0_52_2_a(.in(far_0_52_1[0]), .out(far_0_52_2[0]));    relay_conn far_0_52_2_b(.in(far_0_52_1[1]), .out(far_0_52_2[1]));
    assign layer_0[52] = far_0_52_2[0] | far_0_52_2[1]; 
    wire [1:0] far_0_53_0;    relay_conn far_0_53_0_a(.in(in[199]), .out(far_0_53_0[0]));    relay_conn far_0_53_0_b(.in(in[74]), .out(far_0_53_0[1]));
    wire [1:0] far_0_53_1;    relay_conn far_0_53_1_a(.in(far_0_53_0[0]), .out(far_0_53_1[0]));    relay_conn far_0_53_1_b(.in(far_0_53_0[1]), .out(far_0_53_1[1]));
    wire [1:0] far_0_53_2;    relay_conn far_0_53_2_a(.in(far_0_53_1[0]), .out(far_0_53_2[0]));    relay_conn far_0_53_2_b(.in(far_0_53_1[1]), .out(far_0_53_2[1]));
    assign layer_0[53] = far_0_53_2[1]; 
    wire [1:0] far_0_54_0;    relay_conn far_0_54_0_a(.in(in[193]), .out(far_0_54_0[0]));    relay_conn far_0_54_0_b(.in(in[119]), .out(far_0_54_0[1]));
    wire [1:0] far_0_54_1;    relay_conn far_0_54_1_a(.in(far_0_54_0[0]), .out(far_0_54_1[0]));    relay_conn far_0_54_1_b(.in(far_0_54_0[1]), .out(far_0_54_1[1]));
    assign layer_0[54] = far_0_54_1[0] & ~far_0_54_1[1]; 
    wire [1:0] far_0_55_0;    relay_conn far_0_55_0_a(.in(in[66]), .out(far_0_55_0[0]));    relay_conn far_0_55_0_b(.in(in[186]), .out(far_0_55_0[1]));
    wire [1:0] far_0_55_1;    relay_conn far_0_55_1_a(.in(far_0_55_0[0]), .out(far_0_55_1[0]));    relay_conn far_0_55_1_b(.in(far_0_55_0[1]), .out(far_0_55_1[1]));
    wire [1:0] far_0_55_2;    relay_conn far_0_55_2_a(.in(far_0_55_1[0]), .out(far_0_55_2[0]));    relay_conn far_0_55_2_b(.in(far_0_55_1[1]), .out(far_0_55_2[1]));
    assign layer_0[55] = far_0_55_2[0] & far_0_55_2[1]; 
    wire [1:0] far_0_56_0;    relay_conn far_0_56_0_a(.in(in[17]), .out(far_0_56_0[0]));    relay_conn far_0_56_0_b(.in(in[55]), .out(far_0_56_0[1]));
    assign layer_0[56] = far_0_56_0[1]; 
    wire [1:0] far_0_57_0;    relay_conn far_0_57_0_a(.in(in[215]), .out(far_0_57_0[0]));    relay_conn far_0_57_0_b(.in(in[121]), .out(far_0_57_0[1]));
    wire [1:0] far_0_57_1;    relay_conn far_0_57_1_a(.in(far_0_57_0[0]), .out(far_0_57_1[0]));    relay_conn far_0_57_1_b(.in(far_0_57_0[1]), .out(far_0_57_1[1]));
    assign layer_0[57] = ~far_0_57_1[1] | (far_0_57_1[0] & far_0_57_1[1]); 
    wire [1:0] far_0_58_0;    relay_conn far_0_58_0_a(.in(in[133]), .out(far_0_58_0[0]));    relay_conn far_0_58_0_b(.in(in[247]), .out(far_0_58_0[1]));
    wire [1:0] far_0_58_1;    relay_conn far_0_58_1_a(.in(far_0_58_0[0]), .out(far_0_58_1[0]));    relay_conn far_0_58_1_b(.in(far_0_58_0[1]), .out(far_0_58_1[1]));
    wire [1:0] far_0_58_2;    relay_conn far_0_58_2_a(.in(far_0_58_1[0]), .out(far_0_58_2[0]));    relay_conn far_0_58_2_b(.in(far_0_58_1[1]), .out(far_0_58_2[1]));
    assign layer_0[58] = ~(far_0_58_2[0] ^ far_0_58_2[1]); 
    assign layer_0[59] = ~(in[18] | in[48]); 
    wire [1:0] far_0_60_0;    relay_conn far_0_60_0_a(.in(in[95]), .out(far_0_60_0[0]));    relay_conn far_0_60_0_b(.in(in[34]), .out(far_0_60_0[1]));
    assign layer_0[60] = ~far_0_60_0[1]; 
    wire [1:0] far_0_61_0;    relay_conn far_0_61_0_a(.in(in[88]), .out(far_0_61_0[0]));    relay_conn far_0_61_0_b(.in(in[199]), .out(far_0_61_0[1]));
    wire [1:0] far_0_61_1;    relay_conn far_0_61_1_a(.in(far_0_61_0[0]), .out(far_0_61_1[0]));    relay_conn far_0_61_1_b(.in(far_0_61_0[1]), .out(far_0_61_1[1]));
    wire [1:0] far_0_61_2;    relay_conn far_0_61_2_a(.in(far_0_61_1[0]), .out(far_0_61_2[0]));    relay_conn far_0_61_2_b(.in(far_0_61_1[1]), .out(far_0_61_2[1]));
    assign layer_0[61] = far_0_61_2[1] & ~far_0_61_2[0]; 
    wire [1:0] far_0_62_0;    relay_conn far_0_62_0_a(.in(in[74]), .out(far_0_62_0[0]));    relay_conn far_0_62_0_b(.in(in[121]), .out(far_0_62_0[1]));
    assign layer_0[62] = far_0_62_0[0] & ~far_0_62_0[1]; 
    wire [1:0] far_0_63_0;    relay_conn far_0_63_0_a(.in(in[202]), .out(far_0_63_0[0]));    relay_conn far_0_63_0_b(.in(in[250]), .out(far_0_63_0[1]));
    assign layer_0[63] = ~far_0_63_0[1]; 
    wire [1:0] far_0_64_0;    relay_conn far_0_64_0_a(.in(in[3]), .out(far_0_64_0[0]));    relay_conn far_0_64_0_b(.in(in[113]), .out(far_0_64_0[1]));
    wire [1:0] far_0_64_1;    relay_conn far_0_64_1_a(.in(far_0_64_0[0]), .out(far_0_64_1[0]));    relay_conn far_0_64_1_b(.in(far_0_64_0[1]), .out(far_0_64_1[1]));
    wire [1:0] far_0_64_2;    relay_conn far_0_64_2_a(.in(far_0_64_1[0]), .out(far_0_64_2[0]));    relay_conn far_0_64_2_b(.in(far_0_64_1[1]), .out(far_0_64_2[1]));
    assign layer_0[64] = far_0_64_2[0] & ~far_0_64_2[1]; 
    wire [1:0] far_0_65_0;    relay_conn far_0_65_0_a(.in(in[113]), .out(far_0_65_0[0]));    relay_conn far_0_65_0_b(.in(in[51]), .out(far_0_65_0[1]));
    assign layer_0[65] = far_0_65_0[0] | far_0_65_0[1]; 
    assign layer_0[66] = ~in[59] | (in[59] & in[89]); 
    wire [1:0] far_0_67_0;    relay_conn far_0_67_0_a(.in(in[0]), .out(far_0_67_0[0]));    relay_conn far_0_67_0_b(.in(in[125]), .out(far_0_67_0[1]));
    wire [1:0] far_0_67_1;    relay_conn far_0_67_1_a(.in(far_0_67_0[0]), .out(far_0_67_1[0]));    relay_conn far_0_67_1_b(.in(far_0_67_0[1]), .out(far_0_67_1[1]));
    wire [1:0] far_0_67_2;    relay_conn far_0_67_2_a(.in(far_0_67_1[0]), .out(far_0_67_2[0]));    relay_conn far_0_67_2_b(.in(far_0_67_1[1]), .out(far_0_67_2[1]));
    assign layer_0[67] = ~(far_0_67_2[0] ^ far_0_67_2[1]); 
    wire [1:0] far_0_68_0;    relay_conn far_0_68_0_a(.in(in[97]), .out(far_0_68_0[0]));    relay_conn far_0_68_0_b(.in(in[221]), .out(far_0_68_0[1]));
    wire [1:0] far_0_68_1;    relay_conn far_0_68_1_a(.in(far_0_68_0[0]), .out(far_0_68_1[0]));    relay_conn far_0_68_1_b(.in(far_0_68_0[1]), .out(far_0_68_1[1]));
    wire [1:0] far_0_68_2;    relay_conn far_0_68_2_a(.in(far_0_68_1[0]), .out(far_0_68_2[0]));    relay_conn far_0_68_2_b(.in(far_0_68_1[1]), .out(far_0_68_2[1]));
    assign layer_0[68] = far_0_68_2[0] & far_0_68_2[1]; 
    wire [1:0] far_0_69_0;    relay_conn far_0_69_0_a(.in(in[163]), .out(far_0_69_0[0]));    relay_conn far_0_69_0_b(.in(in[238]), .out(far_0_69_0[1]));
    wire [1:0] far_0_69_1;    relay_conn far_0_69_1_a(.in(far_0_69_0[0]), .out(far_0_69_1[0]));    relay_conn far_0_69_1_b(.in(far_0_69_0[1]), .out(far_0_69_1[1]));
    assign layer_0[69] = far_0_69_1[1]; 
    wire [1:0] far_0_70_0;    relay_conn far_0_70_0_a(.in(in[151]), .out(far_0_70_0[0]));    relay_conn far_0_70_0_b(.in(in[59]), .out(far_0_70_0[1]));
    wire [1:0] far_0_70_1;    relay_conn far_0_70_1_a(.in(far_0_70_0[0]), .out(far_0_70_1[0]));    relay_conn far_0_70_1_b(.in(far_0_70_0[1]), .out(far_0_70_1[1]));
    assign layer_0[70] = far_0_70_1[0] & ~far_0_70_1[1]; 
    wire [1:0] far_0_71_0;    relay_conn far_0_71_0_a(.in(in[239]), .out(far_0_71_0[0]));    relay_conn far_0_71_0_b(.in(in[164]), .out(far_0_71_0[1]));
    wire [1:0] far_0_71_1;    relay_conn far_0_71_1_a(.in(far_0_71_0[0]), .out(far_0_71_1[0]));    relay_conn far_0_71_1_b(.in(far_0_71_0[1]), .out(far_0_71_1[1]));
    assign layer_0[71] = ~far_0_71_1[1] | (far_0_71_1[0] & far_0_71_1[1]); 
    wire [1:0] far_0_72_0;    relay_conn far_0_72_0_a(.in(in[251]), .out(far_0_72_0[0]));    relay_conn far_0_72_0_b(.in(in[125]), .out(far_0_72_0[1]));
    wire [1:0] far_0_72_1;    relay_conn far_0_72_1_a(.in(far_0_72_0[0]), .out(far_0_72_1[0]));    relay_conn far_0_72_1_b(.in(far_0_72_0[1]), .out(far_0_72_1[1]));
    wire [1:0] far_0_72_2;    relay_conn far_0_72_2_a(.in(far_0_72_1[0]), .out(far_0_72_2[0]));    relay_conn far_0_72_2_b(.in(far_0_72_1[1]), .out(far_0_72_2[1]));
    assign layer_0[72] = far_0_72_2[0]; 
    wire [1:0] far_0_73_0;    relay_conn far_0_73_0_a(.in(in[166]), .out(far_0_73_0[0]));    relay_conn far_0_73_0_b(.in(in[122]), .out(far_0_73_0[1]));
    assign layer_0[73] = far_0_73_0[1] & ~far_0_73_0[0]; 
    wire [1:0] far_0_74_0;    relay_conn far_0_74_0_a(.in(in[239]), .out(far_0_74_0[0]));    relay_conn far_0_74_0_b(.in(in[199]), .out(far_0_74_0[1]));
    assign layer_0[74] = far_0_74_0[0] | far_0_74_0[1]; 
    wire [1:0] far_0_75_0;    relay_conn far_0_75_0_a(.in(in[5]), .out(far_0_75_0[0]));    relay_conn far_0_75_0_b(.in(in[102]), .out(far_0_75_0[1]));
    wire [1:0] far_0_75_1;    relay_conn far_0_75_1_a(.in(far_0_75_0[0]), .out(far_0_75_1[0]));    relay_conn far_0_75_1_b(.in(far_0_75_0[1]), .out(far_0_75_1[1]));
    wire [1:0] far_0_75_2;    relay_conn far_0_75_2_a(.in(far_0_75_1[0]), .out(far_0_75_2[0]));    relay_conn far_0_75_2_b(.in(far_0_75_1[1]), .out(far_0_75_2[1]));
    assign layer_0[75] = far_0_75_2[1]; 
    wire [1:0] far_0_76_0;    relay_conn far_0_76_0_a(.in(in[37]), .out(far_0_76_0[0]));    relay_conn far_0_76_0_b(.in(in[113]), .out(far_0_76_0[1]));
    wire [1:0] far_0_76_1;    relay_conn far_0_76_1_a(.in(far_0_76_0[0]), .out(far_0_76_1[0]));    relay_conn far_0_76_1_b(.in(far_0_76_0[1]), .out(far_0_76_1[1]));
    assign layer_0[76] = far_0_76_1[0]; 
    assign layer_0[77] = ~(in[174] ^ in[196]); 
    assign layer_0[78] = ~(in[188] ^ in[219]); 
    assign layer_0[79] = in[239] | in[236]; 
    wire [1:0] far_0_80_0;    relay_conn far_0_80_0_a(.in(in[175]), .out(far_0_80_0[0]));    relay_conn far_0_80_0_b(.in(in[109]), .out(far_0_80_0[1]));
    wire [1:0] far_0_80_1;    relay_conn far_0_80_1_a(.in(far_0_80_0[0]), .out(far_0_80_1[0]));    relay_conn far_0_80_1_b(.in(far_0_80_0[1]), .out(far_0_80_1[1]));
    assign layer_0[80] = ~(far_0_80_1[0] | far_0_80_1[1]); 
    wire [1:0] far_0_81_0;    relay_conn far_0_81_0_a(.in(in[121]), .out(far_0_81_0[0]));    relay_conn far_0_81_0_b(.in(in[174]), .out(far_0_81_0[1]));
    assign layer_0[81] = far_0_81_0[0]; 
    wire [1:0] far_0_82_0;    relay_conn far_0_82_0_a(.in(in[212]), .out(far_0_82_0[0]));    relay_conn far_0_82_0_b(.in(in[136]), .out(far_0_82_0[1]));
    wire [1:0] far_0_82_1;    relay_conn far_0_82_1_a(.in(far_0_82_0[0]), .out(far_0_82_1[0]));    relay_conn far_0_82_1_b(.in(far_0_82_0[1]), .out(far_0_82_1[1]));
    assign layer_0[82] = ~far_0_82_1[0]; 
    wire [1:0] far_0_83_0;    relay_conn far_0_83_0_a(.in(in[83]), .out(far_0_83_0[0]));    relay_conn far_0_83_0_b(.in(in[138]), .out(far_0_83_0[1]));
    assign layer_0[83] = ~far_0_83_0[0] | (far_0_83_0[0] & far_0_83_0[1]); 
    wire [1:0] far_0_84_0;    relay_conn far_0_84_0_a(.in(in[151]), .out(far_0_84_0[0]));    relay_conn far_0_84_0_b(.in(in[199]), .out(far_0_84_0[1]));
    assign layer_0[84] = ~(far_0_84_0[0] & far_0_84_0[1]); 
    assign layer_0[85] = in[215] & ~in[226]; 
    wire [1:0] far_0_86_0;    relay_conn far_0_86_0_a(.in(in[51]), .out(far_0_86_0[0]));    relay_conn far_0_86_0_b(.in(in[96]), .out(far_0_86_0[1]));
    assign layer_0[86] = ~(far_0_86_0[0] & far_0_86_0[1]); 
    wire [1:0] far_0_87_0;    relay_conn far_0_87_0_a(.in(in[72]), .out(far_0_87_0[0]));    relay_conn far_0_87_0_b(.in(in[199]), .out(far_0_87_0[1]));
    wire [1:0] far_0_87_1;    relay_conn far_0_87_1_a(.in(far_0_87_0[0]), .out(far_0_87_1[0]));    relay_conn far_0_87_1_b(.in(far_0_87_0[1]), .out(far_0_87_1[1]));
    wire [1:0] far_0_87_2;    relay_conn far_0_87_2_a(.in(far_0_87_1[0]), .out(far_0_87_2[0]));    relay_conn far_0_87_2_b(.in(far_0_87_1[1]), .out(far_0_87_2[1]));
    assign layer_0[87] = far_0_87_2[0] ^ far_0_87_2[1]; 
    assign layer_0[88] = ~(in[221] | in[212]); 
    assign layer_0[89] = in[10]; 
    wire [1:0] far_0_90_0;    relay_conn far_0_90_0_a(.in(in[199]), .out(far_0_90_0[0]));    relay_conn far_0_90_0_b(.in(in[254]), .out(far_0_90_0[1]));
    assign layer_0[90] = ~far_0_90_0[1] | (far_0_90_0[0] & far_0_90_0[1]); 
    assign layer_0[91] = in[213]; 
    wire [1:0] far_0_92_0;    relay_conn far_0_92_0_a(.in(in[125]), .out(far_0_92_0[0]));    relay_conn far_0_92_0_b(.in(in[207]), .out(far_0_92_0[1]));
    wire [1:0] far_0_92_1;    relay_conn far_0_92_1_a(.in(far_0_92_0[0]), .out(far_0_92_1[0]));    relay_conn far_0_92_1_b(.in(far_0_92_0[1]), .out(far_0_92_1[1]));
    assign layer_0[92] = ~far_0_92_1[1]; 
    wire [1:0] far_0_93_0;    relay_conn far_0_93_0_a(.in(in[89]), .out(far_0_93_0[0]));    relay_conn far_0_93_0_b(.in(in[56]), .out(far_0_93_0[1]));
    assign layer_0[93] = far_0_93_0[1]; 
    wire [1:0] far_0_94_0;    relay_conn far_0_94_0_a(.in(in[70]), .out(far_0_94_0[0]));    relay_conn far_0_94_0_b(.in(in[134]), .out(far_0_94_0[1]));
    wire [1:0] far_0_94_1;    relay_conn far_0_94_1_a(.in(far_0_94_0[0]), .out(far_0_94_1[0]));    relay_conn far_0_94_1_b(.in(far_0_94_0[1]), .out(far_0_94_1[1]));
    assign layer_0[94] = ~far_0_94_1[0]; 
    wire [1:0] far_0_95_0;    relay_conn far_0_95_0_a(.in(in[91]), .out(far_0_95_0[0]));    relay_conn far_0_95_0_b(.in(in[207]), .out(far_0_95_0[1]));
    wire [1:0] far_0_95_1;    relay_conn far_0_95_1_a(.in(far_0_95_0[0]), .out(far_0_95_1[0]));    relay_conn far_0_95_1_b(.in(far_0_95_0[1]), .out(far_0_95_1[1]));
    wire [1:0] far_0_95_2;    relay_conn far_0_95_2_a(.in(far_0_95_1[0]), .out(far_0_95_2[0]));    relay_conn far_0_95_2_b(.in(far_0_95_1[1]), .out(far_0_95_2[1]));
    assign layer_0[95] = far_0_95_2[0] & far_0_95_2[1]; 
    wire [1:0] far_0_96_0;    relay_conn far_0_96_0_a(.in(in[189]), .out(far_0_96_0[0]));    relay_conn far_0_96_0_b(.in(in[136]), .out(far_0_96_0[1]));
    assign layer_0[96] = far_0_96_0[0]; 
    assign layer_0[97] = in[117]; 
    wire [1:0] far_0_98_0;    relay_conn far_0_98_0_a(.in(in[173]), .out(far_0_98_0[0]));    relay_conn far_0_98_0_b(.in(in[111]), .out(far_0_98_0[1]));
    assign layer_0[98] = far_0_98_0[0] & ~far_0_98_0[1]; 
    assign layer_0[99] = in[101]; 
    wire [1:0] far_0_100_0;    relay_conn far_0_100_0_a(.in(in[198]), .out(far_0_100_0[0]));    relay_conn far_0_100_0_b(.in(in[150]), .out(far_0_100_0[1]));
    assign layer_0[100] = far_0_100_0[0] | far_0_100_0[1]; 
    assign layer_0[101] = ~(in[36] ^ in[38]); 
    wire [1:0] far_0_102_0;    relay_conn far_0_102_0_a(.in(in[133]), .out(far_0_102_0[0]));    relay_conn far_0_102_0_b(.in(in[29]), .out(far_0_102_0[1]));
    wire [1:0] far_0_102_1;    relay_conn far_0_102_1_a(.in(far_0_102_0[0]), .out(far_0_102_1[0]));    relay_conn far_0_102_1_b(.in(far_0_102_0[1]), .out(far_0_102_1[1]));
    wire [1:0] far_0_102_2;    relay_conn far_0_102_2_a(.in(far_0_102_1[0]), .out(far_0_102_2[0]));    relay_conn far_0_102_2_b(.in(far_0_102_1[1]), .out(far_0_102_2[1]));
    assign layer_0[102] = far_0_102_2[0] & ~far_0_102_2[1]; 
    wire [1:0] far_0_103_0;    relay_conn far_0_103_0_a(.in(in[48]), .out(far_0_103_0[0]));    relay_conn far_0_103_0_b(.in(in[157]), .out(far_0_103_0[1]));
    wire [1:0] far_0_103_1;    relay_conn far_0_103_1_a(.in(far_0_103_0[0]), .out(far_0_103_1[0]));    relay_conn far_0_103_1_b(.in(far_0_103_0[1]), .out(far_0_103_1[1]));
    wire [1:0] far_0_103_2;    relay_conn far_0_103_2_a(.in(far_0_103_1[0]), .out(far_0_103_2[0]));    relay_conn far_0_103_2_b(.in(far_0_103_1[1]), .out(far_0_103_2[1]));
    assign layer_0[103] = far_0_103_2[0] & far_0_103_2[1]; 
    wire [1:0] far_0_104_0;    relay_conn far_0_104_0_a(.in(in[241]), .out(far_0_104_0[0]));    relay_conn far_0_104_0_b(.in(in[164]), .out(far_0_104_0[1]));
    wire [1:0] far_0_104_1;    relay_conn far_0_104_1_a(.in(far_0_104_0[0]), .out(far_0_104_1[0]));    relay_conn far_0_104_1_b(.in(far_0_104_0[1]), .out(far_0_104_1[1]));
    assign layer_0[104] = far_0_104_1[1]; 
    wire [1:0] far_0_105_0;    relay_conn far_0_105_0_a(.in(in[108]), .out(far_0_105_0[0]));    relay_conn far_0_105_0_b(.in(in[17]), .out(far_0_105_0[1]));
    wire [1:0] far_0_105_1;    relay_conn far_0_105_1_a(.in(far_0_105_0[0]), .out(far_0_105_1[0]));    relay_conn far_0_105_1_b(.in(far_0_105_0[1]), .out(far_0_105_1[1]));
    assign layer_0[105] = ~(far_0_105_1[0] ^ far_0_105_1[1]); 
    wire [1:0] far_0_106_0;    relay_conn far_0_106_0_a(.in(in[211]), .out(far_0_106_0[0]));    relay_conn far_0_106_0_b(.in(in[247]), .out(far_0_106_0[1]));
    assign layer_0[106] = far_0_106_0[0] & ~far_0_106_0[1]; 
    wire [1:0] far_0_107_0;    relay_conn far_0_107_0_a(.in(in[84]), .out(far_0_107_0[0]));    relay_conn far_0_107_0_b(.in(in[166]), .out(far_0_107_0[1]));
    wire [1:0] far_0_107_1;    relay_conn far_0_107_1_a(.in(far_0_107_0[0]), .out(far_0_107_1[0]));    relay_conn far_0_107_1_b(.in(far_0_107_0[1]), .out(far_0_107_1[1]));
    assign layer_0[107] = far_0_107_1[0] | far_0_107_1[1]; 
    assign layer_0[108] = ~in[88] | (in[88] & in[78]); 
    wire [1:0] far_0_109_0;    relay_conn far_0_109_0_a(.in(in[253]), .out(far_0_109_0[0]));    relay_conn far_0_109_0_b(.in(in[219]), .out(far_0_109_0[1]));
    assign layer_0[109] = far_0_109_0[1] & ~far_0_109_0[0]; 
    assign layer_0[110] = ~in[183]; 
    wire [1:0] far_0_111_0;    relay_conn far_0_111_0_a(.in(in[97]), .out(far_0_111_0[0]));    relay_conn far_0_111_0_b(.in(in[34]), .out(far_0_111_0[1]));
    assign layer_0[111] = ~(far_0_111_0[0] & far_0_111_0[1]); 
    assign layer_0[112] = in[241] & ~in[249]; 
    assign layer_0[113] = in[199]; 
    wire [1:0] far_0_114_0;    relay_conn far_0_114_0_a(.in(in[150]), .out(far_0_114_0[0]));    relay_conn far_0_114_0_b(.in(in[254]), .out(far_0_114_0[1]));
    wire [1:0] far_0_114_1;    relay_conn far_0_114_1_a(.in(far_0_114_0[0]), .out(far_0_114_1[0]));    relay_conn far_0_114_1_b(.in(far_0_114_0[1]), .out(far_0_114_1[1]));
    wire [1:0] far_0_114_2;    relay_conn far_0_114_2_a(.in(far_0_114_1[0]), .out(far_0_114_2[0]));    relay_conn far_0_114_2_b(.in(far_0_114_1[1]), .out(far_0_114_2[1]));
    assign layer_0[114] = ~(far_0_114_2[0] & far_0_114_2[1]); 
    wire [1:0] far_0_115_0;    relay_conn far_0_115_0_a(.in(in[104]), .out(far_0_115_0[0]));    relay_conn far_0_115_0_b(.in(in[164]), .out(far_0_115_0[1]));
    assign layer_0[115] = ~(far_0_115_0[0] ^ far_0_115_0[1]); 
    assign layer_0[116] = ~(in[30] ^ in[28]); 
    assign layer_0[117] = in[138] & ~in[125]; 
    assign layer_0[118] = ~in[153] | (in[125] & in[153]); 
    wire [1:0] far_0_119_0;    relay_conn far_0_119_0_a(.in(in[132]), .out(far_0_119_0[0]));    relay_conn far_0_119_0_b(.in(in[199]), .out(far_0_119_0[1]));
    wire [1:0] far_0_119_1;    relay_conn far_0_119_1_a(.in(far_0_119_0[0]), .out(far_0_119_1[0]));    relay_conn far_0_119_1_b(.in(far_0_119_0[1]), .out(far_0_119_1[1]));
    assign layer_0[119] = ~far_0_119_1[0]; 
    wire [1:0] far_0_120_0;    relay_conn far_0_120_0_a(.in(in[216]), .out(far_0_120_0[0]));    relay_conn far_0_120_0_b(.in(in[167]), .out(far_0_120_0[1]));
    assign layer_0[120] = far_0_120_0[0] ^ far_0_120_0[1]; 
    assign layer_0[121] = ~(in[83] ^ in[81]); 
    wire [1:0] far_0_122_0;    relay_conn far_0_122_0_a(.in(in[199]), .out(far_0_122_0[0]));    relay_conn far_0_122_0_b(.in(in[149]), .out(far_0_122_0[1]));
    assign layer_0[122] = ~far_0_122_0[1] | (far_0_122_0[0] & far_0_122_0[1]); 
    wire [1:0] far_0_123_0;    relay_conn far_0_123_0_a(.in(in[99]), .out(far_0_123_0[0]));    relay_conn far_0_123_0_b(.in(in[186]), .out(far_0_123_0[1]));
    wire [1:0] far_0_123_1;    relay_conn far_0_123_1_a(.in(far_0_123_0[0]), .out(far_0_123_1[0]));    relay_conn far_0_123_1_b(.in(far_0_123_0[1]), .out(far_0_123_1[1]));
    assign layer_0[123] = far_0_123_1[0] & far_0_123_1[1]; 
    wire [1:0] far_0_124_0;    relay_conn far_0_124_0_a(.in(in[215]), .out(far_0_124_0[0]));    relay_conn far_0_124_0_b(.in(in[172]), .out(far_0_124_0[1]));
    assign layer_0[124] = far_0_124_0[0] | far_0_124_0[1]; 
    wire [1:0] far_0_125_0;    relay_conn far_0_125_0_a(.in(in[186]), .out(far_0_125_0[0]));    relay_conn far_0_125_0_b(.in(in[140]), .out(far_0_125_0[1]));
    assign layer_0[125] = far_0_125_0[1]; 
    wire [1:0] far_0_126_0;    relay_conn far_0_126_0_a(.in(in[63]), .out(far_0_126_0[0]));    relay_conn far_0_126_0_b(.in(in[113]), .out(far_0_126_0[1]));
    assign layer_0[126] = far_0_126_0[0] | far_0_126_0[1]; 
    assign layer_0[127] = in[56]; 
    assign layer_0[128] = ~in[31] | (in[48] & in[31]); 
    wire [1:0] far_0_129_0;    relay_conn far_0_129_0_a(.in(in[172]), .out(far_0_129_0[0]));    relay_conn far_0_129_0_b(.in(in[92]), .out(far_0_129_0[1]));
    wire [1:0] far_0_129_1;    relay_conn far_0_129_1_a(.in(far_0_129_0[0]), .out(far_0_129_1[0]));    relay_conn far_0_129_1_b(.in(far_0_129_0[1]), .out(far_0_129_1[1]));
    assign layer_0[129] = far_0_129_1[0] & far_0_129_1[1]; 
    wire [1:0] far_0_130_0;    relay_conn far_0_130_0_a(.in(in[205]), .out(far_0_130_0[0]));    relay_conn far_0_130_0_b(.in(in[135]), .out(far_0_130_0[1]));
    wire [1:0] far_0_130_1;    relay_conn far_0_130_1_a(.in(far_0_130_0[0]), .out(far_0_130_1[0]));    relay_conn far_0_130_1_b(.in(far_0_130_0[1]), .out(far_0_130_1[1]));
    assign layer_0[130] = far_0_130_1[1]; 
    wire [1:0] far_0_131_0;    relay_conn far_0_131_0_a(.in(in[169]), .out(far_0_131_0[0]));    relay_conn far_0_131_0_b(.in(in[57]), .out(far_0_131_0[1]));
    wire [1:0] far_0_131_1;    relay_conn far_0_131_1_a(.in(far_0_131_0[0]), .out(far_0_131_1[0]));    relay_conn far_0_131_1_b(.in(far_0_131_0[1]), .out(far_0_131_1[1]));
    wire [1:0] far_0_131_2;    relay_conn far_0_131_2_a(.in(far_0_131_1[0]), .out(far_0_131_2[0]));    relay_conn far_0_131_2_b(.in(far_0_131_1[1]), .out(far_0_131_2[1]));
    assign layer_0[131] = far_0_131_2[0] | far_0_131_2[1]; 
    wire [1:0] far_0_132_0;    relay_conn far_0_132_0_a(.in(in[42]), .out(far_0_132_0[0]));    relay_conn far_0_132_0_b(.in(in[157]), .out(far_0_132_0[1]));
    wire [1:0] far_0_132_1;    relay_conn far_0_132_1_a(.in(far_0_132_0[0]), .out(far_0_132_1[0]));    relay_conn far_0_132_1_b(.in(far_0_132_0[1]), .out(far_0_132_1[1]));
    wire [1:0] far_0_132_2;    relay_conn far_0_132_2_a(.in(far_0_132_1[0]), .out(far_0_132_2[0]));    relay_conn far_0_132_2_b(.in(far_0_132_1[1]), .out(far_0_132_2[1]));
    assign layer_0[132] = far_0_132_2[0] | far_0_132_2[1]; 
    wire [1:0] far_0_133_0;    relay_conn far_0_133_0_a(.in(in[222]), .out(far_0_133_0[0]));    relay_conn far_0_133_0_b(.in(in[185]), .out(far_0_133_0[1]));
    assign layer_0[133] = ~(far_0_133_0[0] & far_0_133_0[1]); 
    wire [1:0] far_0_134_0;    relay_conn far_0_134_0_a(.in(in[72]), .out(far_0_134_0[0]));    relay_conn far_0_134_0_b(.in(in[134]), .out(far_0_134_0[1]));
    assign layer_0[134] = ~(far_0_134_0[0] | far_0_134_0[1]); 
    wire [1:0] far_0_135_0;    relay_conn far_0_135_0_a(.in(in[84]), .out(far_0_135_0[0]));    relay_conn far_0_135_0_b(.in(in[199]), .out(far_0_135_0[1]));
    wire [1:0] far_0_135_1;    relay_conn far_0_135_1_a(.in(far_0_135_0[0]), .out(far_0_135_1[0]));    relay_conn far_0_135_1_b(.in(far_0_135_0[1]), .out(far_0_135_1[1]));
    wire [1:0] far_0_135_2;    relay_conn far_0_135_2_a(.in(far_0_135_1[0]), .out(far_0_135_2[0]));    relay_conn far_0_135_2_b(.in(far_0_135_1[1]), .out(far_0_135_2[1]));
    assign layer_0[135] = far_0_135_2[0] & ~far_0_135_2[1]; 
    wire [1:0] far_0_136_0;    relay_conn far_0_136_0_a(.in(in[172]), .out(far_0_136_0[0]));    relay_conn far_0_136_0_b(.in(in[66]), .out(far_0_136_0[1]));
    wire [1:0] far_0_136_1;    relay_conn far_0_136_1_a(.in(far_0_136_0[0]), .out(far_0_136_1[0]));    relay_conn far_0_136_1_b(.in(far_0_136_0[1]), .out(far_0_136_1[1]));
    wire [1:0] far_0_136_2;    relay_conn far_0_136_2_a(.in(far_0_136_1[0]), .out(far_0_136_2[0]));    relay_conn far_0_136_2_b(.in(far_0_136_1[1]), .out(far_0_136_2[1]));
    assign layer_0[136] = far_0_136_2[0] & far_0_136_2[1]; 
    wire [1:0] far_0_137_0;    relay_conn far_0_137_0_a(.in(in[117]), .out(far_0_137_0[0]));    relay_conn far_0_137_0_b(.in(in[176]), .out(far_0_137_0[1]));
    assign layer_0[137] = ~(far_0_137_0[0] ^ far_0_137_0[1]); 
    wire [1:0] far_0_138_0;    relay_conn far_0_138_0_a(.in(in[125]), .out(far_0_138_0[0]));    relay_conn far_0_138_0_b(.in(in[71]), .out(far_0_138_0[1]));
    assign layer_0[138] = ~(far_0_138_0[0] | far_0_138_0[1]); 
    wire [1:0] far_0_139_0;    relay_conn far_0_139_0_a(.in(in[102]), .out(far_0_139_0[0]));    relay_conn far_0_139_0_b(.in(in[221]), .out(far_0_139_0[1]));
    wire [1:0] far_0_139_1;    relay_conn far_0_139_1_a(.in(far_0_139_0[0]), .out(far_0_139_1[0]));    relay_conn far_0_139_1_b(.in(far_0_139_0[1]), .out(far_0_139_1[1]));
    wire [1:0] far_0_139_2;    relay_conn far_0_139_2_a(.in(far_0_139_1[0]), .out(far_0_139_2[0]));    relay_conn far_0_139_2_b(.in(far_0_139_1[1]), .out(far_0_139_2[1]));
    assign layer_0[139] = far_0_139_2[0] & far_0_139_2[1]; 
    wire [1:0] far_0_140_0;    relay_conn far_0_140_0_a(.in(in[130]), .out(far_0_140_0[0]));    relay_conn far_0_140_0_b(.in(in[234]), .out(far_0_140_0[1]));
    wire [1:0] far_0_140_1;    relay_conn far_0_140_1_a(.in(far_0_140_0[0]), .out(far_0_140_1[0]));    relay_conn far_0_140_1_b(.in(far_0_140_0[1]), .out(far_0_140_1[1]));
    wire [1:0] far_0_140_2;    relay_conn far_0_140_2_a(.in(far_0_140_1[0]), .out(far_0_140_2[0]));    relay_conn far_0_140_2_b(.in(far_0_140_1[1]), .out(far_0_140_2[1]));
    assign layer_0[140] = far_0_140_2[0]; 
    wire [1:0] far_0_141_0;    relay_conn far_0_141_0_a(.in(in[245]), .out(far_0_141_0[0]));    relay_conn far_0_141_0_b(.in(in[125]), .out(far_0_141_0[1]));
    wire [1:0] far_0_141_1;    relay_conn far_0_141_1_a(.in(far_0_141_0[0]), .out(far_0_141_1[0]));    relay_conn far_0_141_1_b(.in(far_0_141_0[1]), .out(far_0_141_1[1]));
    wire [1:0] far_0_141_2;    relay_conn far_0_141_2_a(.in(far_0_141_1[0]), .out(far_0_141_2[0]));    relay_conn far_0_141_2_b(.in(far_0_141_1[1]), .out(far_0_141_2[1]));
    assign layer_0[141] = far_0_141_2[0] & far_0_141_2[1]; 
    assign layer_0[142] = ~(in[16] & in[15]); 
    assign layer_0[143] = ~in[157] | (in[157] & in[158]); 
    assign layer_0[144] = in[21] & in[44]; 
    wire [1:0] far_0_145_0;    relay_conn far_0_145_0_a(.in(in[125]), .out(far_0_145_0[0]));    relay_conn far_0_145_0_b(.in(in[158]), .out(far_0_145_0[1]));
    assign layer_0[145] = far_0_145_0[0] ^ far_0_145_0[1]; 
    wire [1:0] far_0_146_0;    relay_conn far_0_146_0_a(.in(in[117]), .out(far_0_146_0[0]));    relay_conn far_0_146_0_b(.in(in[214]), .out(far_0_146_0[1]));
    wire [1:0] far_0_146_1;    relay_conn far_0_146_1_a(.in(far_0_146_0[0]), .out(far_0_146_1[0]));    relay_conn far_0_146_1_b(.in(far_0_146_0[1]), .out(far_0_146_1[1]));
    wire [1:0] far_0_146_2;    relay_conn far_0_146_2_a(.in(far_0_146_1[0]), .out(far_0_146_2[0]));    relay_conn far_0_146_2_b(.in(far_0_146_1[1]), .out(far_0_146_2[1]));
    assign layer_0[146] = ~far_0_146_2[0]; 
    wire [1:0] far_0_147_0;    relay_conn far_0_147_0_a(.in(in[142]), .out(far_0_147_0[0]));    relay_conn far_0_147_0_b(.in(in[87]), .out(far_0_147_0[1]));
    assign layer_0[147] = far_0_147_0[0] ^ far_0_147_0[1]; 
    wire [1:0] far_0_148_0;    relay_conn far_0_148_0_a(.in(in[17]), .out(far_0_148_0[0]));    relay_conn far_0_148_0_b(.in(in[87]), .out(far_0_148_0[1]));
    wire [1:0] far_0_148_1;    relay_conn far_0_148_1_a(.in(far_0_148_0[0]), .out(far_0_148_1[0]));    relay_conn far_0_148_1_b(.in(far_0_148_0[1]), .out(far_0_148_1[1]));
    assign layer_0[148] = far_0_148_1[1]; 
    assign layer_0[149] = in[214]; 
    assign layer_0[150] = in[221] ^ in[247]; 
    assign layer_0[151] = ~(in[119] ^ in[94]); 
    assign layer_0[152] = ~in[130] | (in[130] & in[119]); 
    assign layer_0[153] = ~(in[151] | in[142]); 
    wire [1:0] far_0_154_0;    relay_conn far_0_154_0_a(.in(in[187]), .out(far_0_154_0[0]));    relay_conn far_0_154_0_b(.in(in[251]), .out(far_0_154_0[1]));
    wire [1:0] far_0_154_1;    relay_conn far_0_154_1_a(.in(far_0_154_0[0]), .out(far_0_154_1[0]));    relay_conn far_0_154_1_b(.in(far_0_154_0[1]), .out(far_0_154_1[1]));
    assign layer_0[154] = far_0_154_1[0] | far_0_154_1[1]; 
    wire [1:0] far_0_155_0;    relay_conn far_0_155_0_a(.in(in[239]), .out(far_0_155_0[0]));    relay_conn far_0_155_0_b(.in(in[127]), .out(far_0_155_0[1]));
    wire [1:0] far_0_155_1;    relay_conn far_0_155_1_a(.in(far_0_155_0[0]), .out(far_0_155_1[0]));    relay_conn far_0_155_1_b(.in(far_0_155_0[1]), .out(far_0_155_1[1]));
    wire [1:0] far_0_155_2;    relay_conn far_0_155_2_a(.in(far_0_155_1[0]), .out(far_0_155_2[0]));    relay_conn far_0_155_2_b(.in(far_0_155_1[1]), .out(far_0_155_2[1]));
    assign layer_0[155] = ~(far_0_155_2[0] & far_0_155_2[1]); 
    assign layer_0[156] = ~(in[57] & in[51]); 
    wire [1:0] far_0_157_0;    relay_conn far_0_157_0_a(.in(in[176]), .out(far_0_157_0[0]));    relay_conn far_0_157_0_b(.in(in[243]), .out(far_0_157_0[1]));
    wire [1:0] far_0_157_1;    relay_conn far_0_157_1_a(.in(far_0_157_0[0]), .out(far_0_157_1[0]));    relay_conn far_0_157_1_b(.in(far_0_157_0[1]), .out(far_0_157_1[1]));
    assign layer_0[157] = ~far_0_157_1[0]; 
    wire [1:0] far_0_158_0;    relay_conn far_0_158_0_a(.in(in[30]), .out(far_0_158_0[0]));    relay_conn far_0_158_0_b(.in(in[125]), .out(far_0_158_0[1]));
    wire [1:0] far_0_158_1;    relay_conn far_0_158_1_a(.in(far_0_158_0[0]), .out(far_0_158_1[0]));    relay_conn far_0_158_1_b(.in(far_0_158_0[1]), .out(far_0_158_1[1]));
    assign layer_0[158] = far_0_158_1[0] & ~far_0_158_1[1]; 
    wire [1:0] far_0_159_0;    relay_conn far_0_159_0_a(.in(in[133]), .out(far_0_159_0[0]));    relay_conn far_0_159_0_b(.in(in[172]), .out(far_0_159_0[1]));
    assign layer_0[159] = ~far_0_159_0[0]; 
    wire [1:0] far_0_160_0;    relay_conn far_0_160_0_a(.in(in[53]), .out(far_0_160_0[0]));    relay_conn far_0_160_0_b(.in(in[181]), .out(far_0_160_0[1]));
    wire [1:0] far_0_160_1;    relay_conn far_0_160_1_a(.in(far_0_160_0[0]), .out(far_0_160_1[0]));    relay_conn far_0_160_1_b(.in(far_0_160_0[1]), .out(far_0_160_1[1]));
    wire [1:0] far_0_160_2;    relay_conn far_0_160_2_a(.in(far_0_160_1[0]), .out(far_0_160_2[0]));    relay_conn far_0_160_2_b(.in(far_0_160_1[1]), .out(far_0_160_2[1]));
    wire [1:0] far_0_160_3;    relay_conn far_0_160_3_a(.in(far_0_160_2[0]), .out(far_0_160_3[0]));    relay_conn far_0_160_3_b(.in(far_0_160_2[1]), .out(far_0_160_3[1]));
    assign layer_0[160] = ~far_0_160_3[1] | (far_0_160_3[0] & far_0_160_3[1]); 
    assign layer_0[161] = ~in[57]; 
    assign layer_0[162] = in[225] & ~in[255]; 
    wire [1:0] far_0_163_0;    relay_conn far_0_163_0_a(.in(in[57]), .out(far_0_163_0[0]));    relay_conn far_0_163_0_b(.in(in[151]), .out(far_0_163_0[1]));
    wire [1:0] far_0_163_1;    relay_conn far_0_163_1_a(.in(far_0_163_0[0]), .out(far_0_163_1[0]));    relay_conn far_0_163_1_b(.in(far_0_163_0[1]), .out(far_0_163_1[1]));
    assign layer_0[163] = far_0_163_1[0] | far_0_163_1[1]; 
    wire [1:0] far_0_164_0;    relay_conn far_0_164_0_a(.in(in[39]), .out(far_0_164_0[0]));    relay_conn far_0_164_0_b(.in(in[117]), .out(far_0_164_0[1]));
    wire [1:0] far_0_164_1;    relay_conn far_0_164_1_a(.in(far_0_164_0[0]), .out(far_0_164_1[0]));    relay_conn far_0_164_1_b(.in(far_0_164_0[1]), .out(far_0_164_1[1]));
    assign layer_0[164] = ~(far_0_164_1[0] ^ far_0_164_1[1]); 
    assign layer_0[165] = in[193]; 
    wire [1:0] far_0_166_0;    relay_conn far_0_166_0_a(.in(in[241]), .out(far_0_166_0[0]));    relay_conn far_0_166_0_b(.in(in[167]), .out(far_0_166_0[1]));
    wire [1:0] far_0_166_1;    relay_conn far_0_166_1_a(.in(far_0_166_0[0]), .out(far_0_166_1[0]));    relay_conn far_0_166_1_b(.in(far_0_166_0[1]), .out(far_0_166_1[1]));
    assign layer_0[166] = ~(far_0_166_1[0] ^ far_0_166_1[1]); 
    wire [1:0] far_0_167_0;    relay_conn far_0_167_0_a(.in(in[79]), .out(far_0_167_0[0]));    relay_conn far_0_167_0_b(.in(in[151]), .out(far_0_167_0[1]));
    wire [1:0] far_0_167_1;    relay_conn far_0_167_1_a(.in(far_0_167_0[0]), .out(far_0_167_1[0]));    relay_conn far_0_167_1_b(.in(far_0_167_0[1]), .out(far_0_167_1[1]));
    assign layer_0[167] = ~(far_0_167_1[0] | far_0_167_1[1]); 
    wire [1:0] far_0_168_0;    relay_conn far_0_168_0_a(.in(in[151]), .out(far_0_168_0[0]));    relay_conn far_0_168_0_b(.in(in[119]), .out(far_0_168_0[1]));
    assign layer_0[168] = ~(far_0_168_0[0] & far_0_168_0[1]); 
    wire [1:0] far_0_169_0;    relay_conn far_0_169_0_a(.in(in[197]), .out(far_0_169_0[0]));    relay_conn far_0_169_0_b(.in(in[151]), .out(far_0_169_0[1]));
    assign layer_0[169] = ~far_0_169_0[0]; 
    assign layer_0[170] = ~(in[57] | in[88]); 
    wire [1:0] far_0_171_0;    relay_conn far_0_171_0_a(.in(in[65]), .out(far_0_171_0[0]));    relay_conn far_0_171_0_b(.in(in[158]), .out(far_0_171_0[1]));
    wire [1:0] far_0_171_1;    relay_conn far_0_171_1_a(.in(far_0_171_0[0]), .out(far_0_171_1[0]));    relay_conn far_0_171_1_b(.in(far_0_171_0[1]), .out(far_0_171_1[1]));
    assign layer_0[171] = far_0_171_1[0]; 
    wire [1:0] far_0_172_0;    relay_conn far_0_172_0_a(.in(in[49]), .out(far_0_172_0[0]));    relay_conn far_0_172_0_b(.in(in[15]), .out(far_0_172_0[1]));
    assign layer_0[172] = ~far_0_172_0[1]; 
    wire [1:0] far_0_173_0;    relay_conn far_0_173_0_a(.in(in[181]), .out(far_0_173_0[0]));    relay_conn far_0_173_0_b(.in(in[250]), .out(far_0_173_0[1]));
    wire [1:0] far_0_173_1;    relay_conn far_0_173_1_a(.in(far_0_173_0[0]), .out(far_0_173_1[0]));    relay_conn far_0_173_1_b(.in(far_0_173_0[1]), .out(far_0_173_1[1]));
    assign layer_0[173] = ~far_0_173_1[0] | (far_0_173_1[0] & far_0_173_1[1]); 
    wire [1:0] far_0_174_0;    relay_conn far_0_174_0_a(.in(in[57]), .out(far_0_174_0[0]));    relay_conn far_0_174_0_b(.in(in[133]), .out(far_0_174_0[1]));
    wire [1:0] far_0_174_1;    relay_conn far_0_174_1_a(.in(far_0_174_0[0]), .out(far_0_174_1[0]));    relay_conn far_0_174_1_b(.in(far_0_174_0[1]), .out(far_0_174_1[1]));
    assign layer_0[174] = far_0_174_1[1]; 
    assign layer_0[175] = ~(in[186] ^ in[207]); 
    wire [1:0] far_0_176_0;    relay_conn far_0_176_0_a(.in(in[109]), .out(far_0_176_0[0]));    relay_conn far_0_176_0_b(.in(in[20]), .out(far_0_176_0[1]));
    wire [1:0] far_0_176_1;    relay_conn far_0_176_1_a(.in(far_0_176_0[0]), .out(far_0_176_1[0]));    relay_conn far_0_176_1_b(.in(far_0_176_0[1]), .out(far_0_176_1[1]));
    assign layer_0[176] = far_0_176_1[0] & far_0_176_1[1]; 
    assign layer_0[177] = ~(in[207] | in[188]); 
    wire [1:0] far_0_178_0;    relay_conn far_0_178_0_a(.in(in[172]), .out(far_0_178_0[0]));    relay_conn far_0_178_0_b(.in(in[250]), .out(far_0_178_0[1]));
    wire [1:0] far_0_178_1;    relay_conn far_0_178_1_a(.in(far_0_178_0[0]), .out(far_0_178_1[0]));    relay_conn far_0_178_1_b(.in(far_0_178_0[1]), .out(far_0_178_1[1]));
    assign layer_0[178] = far_0_178_1[0] & ~far_0_178_1[1]; 
    wire [1:0] far_0_179_0;    relay_conn far_0_179_0_a(.in(in[79]), .out(far_0_179_0[0]));    relay_conn far_0_179_0_b(.in(in[121]), .out(far_0_179_0[1]));
    assign layer_0[179] = far_0_179_0[0] & ~far_0_179_0[1]; 
    wire [1:0] far_0_180_0;    relay_conn far_0_180_0_a(.in(in[101]), .out(far_0_180_0[0]));    relay_conn far_0_180_0_b(.in(in[57]), .out(far_0_180_0[1]));
    assign layer_0[180] = far_0_180_0[0] ^ far_0_180_0[1]; 
    wire [1:0] far_0_181_0;    relay_conn far_0_181_0_a(.in(in[80]), .out(far_0_181_0[0]));    relay_conn far_0_181_0_b(.in(in[119]), .out(far_0_181_0[1]));
    assign layer_0[181] = ~(far_0_181_0[0] ^ far_0_181_0[1]); 
    wire [1:0] far_0_182_0;    relay_conn far_0_182_0_a(.in(in[121]), .out(far_0_182_0[0]));    relay_conn far_0_182_0_b(.in(in[70]), .out(far_0_182_0[1]));
    assign layer_0[182] = far_0_182_0[0] & far_0_182_0[1]; 
    assign layer_0[183] = in[136] ^ in[121]; 
    wire [1:0] far_0_184_0;    relay_conn far_0_184_0_a(.in(in[113]), .out(far_0_184_0[0]));    relay_conn far_0_184_0_b(.in(in[1]), .out(far_0_184_0[1]));
    wire [1:0] far_0_184_1;    relay_conn far_0_184_1_a(.in(far_0_184_0[0]), .out(far_0_184_1[0]));    relay_conn far_0_184_1_b(.in(far_0_184_0[1]), .out(far_0_184_1[1]));
    wire [1:0] far_0_184_2;    relay_conn far_0_184_2_a(.in(far_0_184_1[0]), .out(far_0_184_2[0]));    relay_conn far_0_184_2_b(.in(far_0_184_1[1]), .out(far_0_184_2[1]));
    assign layer_0[184] = far_0_184_2[1]; 
    wire [1:0] far_0_185_0;    relay_conn far_0_185_0_a(.in(in[136]), .out(far_0_185_0[0]));    relay_conn far_0_185_0_b(.in(in[216]), .out(far_0_185_0[1]));
    wire [1:0] far_0_185_1;    relay_conn far_0_185_1_a(.in(far_0_185_0[0]), .out(far_0_185_1[0]));    relay_conn far_0_185_1_b(.in(far_0_185_0[1]), .out(far_0_185_1[1]));
    assign layer_0[185] = far_0_185_1[0]; 
    wire [1:0] far_0_186_0;    relay_conn far_0_186_0_a(.in(in[207]), .out(far_0_186_0[0]));    relay_conn far_0_186_0_b(.in(in[156]), .out(far_0_186_0[1]));
    assign layer_0[186] = far_0_186_0[0] & ~far_0_186_0[1]; 
    wire [1:0] far_0_187_0;    relay_conn far_0_187_0_a(.in(in[207]), .out(far_0_187_0[0]));    relay_conn far_0_187_0_b(.in(in[125]), .out(far_0_187_0[1]));
    wire [1:0] far_0_187_1;    relay_conn far_0_187_1_a(.in(far_0_187_0[0]), .out(far_0_187_1[0]));    relay_conn far_0_187_1_b(.in(far_0_187_0[1]), .out(far_0_187_1[1]));
    assign layer_0[187] = ~far_0_187_1[1]; 
    assign layer_0[188] = ~in[186] | (in[186] & in[160]); 
    wire [1:0] far_0_189_0;    relay_conn far_0_189_0_a(.in(in[145]), .out(far_0_189_0[0]));    relay_conn far_0_189_0_b(.in(in[240]), .out(far_0_189_0[1]));
    wire [1:0] far_0_189_1;    relay_conn far_0_189_1_a(.in(far_0_189_0[0]), .out(far_0_189_1[0]));    relay_conn far_0_189_1_b(.in(far_0_189_0[1]), .out(far_0_189_1[1]));
    assign layer_0[189] = ~far_0_189_1[0] | (far_0_189_1[0] & far_0_189_1[1]); 
    assign layer_0[190] = ~in[123] | (in[151] & in[123]); 
    assign layer_0[191] = in[5] | in[19]; 
    wire [1:0] far_0_192_0;    relay_conn far_0_192_0_a(.in(in[23]), .out(far_0_192_0[0]));    relay_conn far_0_192_0_b(.in(in[76]), .out(far_0_192_0[1]));
    assign layer_0[192] = far_0_192_0[0] | far_0_192_0[1]; 
    wire [1:0] far_0_193_0;    relay_conn far_0_193_0_a(.in(in[8]), .out(far_0_193_0[0]));    relay_conn far_0_193_0_b(.in(in[73]), .out(far_0_193_0[1]));
    wire [1:0] far_0_193_1;    relay_conn far_0_193_1_a(.in(far_0_193_0[0]), .out(far_0_193_1[0]));    relay_conn far_0_193_1_b(.in(far_0_193_0[1]), .out(far_0_193_1[1]));
    assign layer_0[193] = far_0_193_1[0]; 
    wire [1:0] far_0_194_0;    relay_conn far_0_194_0_a(.in(in[254]), .out(far_0_194_0[0]));    relay_conn far_0_194_0_b(.in(in[202]), .out(far_0_194_0[1]));
    assign layer_0[194] = ~far_0_194_0[0]; 
    wire [1:0] far_0_195_0;    relay_conn far_0_195_0_a(.in(in[81]), .out(far_0_195_0[0]));    relay_conn far_0_195_0_b(.in(in[22]), .out(far_0_195_0[1]));
    assign layer_0[195] = ~(far_0_195_0[0] | far_0_195_0[1]); 
    wire [1:0] far_0_196_0;    relay_conn far_0_196_0_a(.in(in[181]), .out(far_0_196_0[0]));    relay_conn far_0_196_0_b(.in(in[215]), .out(far_0_196_0[1]));
    assign layer_0[196] = far_0_196_0[0] & far_0_196_0[1]; 
    wire [1:0] far_0_197_0;    relay_conn far_0_197_0_a(.in(in[179]), .out(far_0_197_0[0]));    relay_conn far_0_197_0_b(.in(in[80]), .out(far_0_197_0[1]));
    wire [1:0] far_0_197_1;    relay_conn far_0_197_1_a(.in(far_0_197_0[0]), .out(far_0_197_1[0]));    relay_conn far_0_197_1_b(.in(far_0_197_0[1]), .out(far_0_197_1[1]));
    wire [1:0] far_0_197_2;    relay_conn far_0_197_2_a(.in(far_0_197_1[0]), .out(far_0_197_2[0]));    relay_conn far_0_197_2_b(.in(far_0_197_1[1]), .out(far_0_197_2[1]));
    assign layer_0[197] = ~far_0_197_2[1]; 
    wire [1:0] far_0_198_0;    relay_conn far_0_198_0_a(.in(in[51]), .out(far_0_198_0[0]));    relay_conn far_0_198_0_b(.in(in[92]), .out(far_0_198_0[1]));
    assign layer_0[198] = far_0_198_0[0] & ~far_0_198_0[1]; 
    assign layer_0[199] = ~(in[34] ^ in[19]); 
    wire [1:0] far_0_200_0;    relay_conn far_0_200_0_a(.in(in[109]), .out(far_0_200_0[0]));    relay_conn far_0_200_0_b(.in(in[5]), .out(far_0_200_0[1]));
    wire [1:0] far_0_200_1;    relay_conn far_0_200_1_a(.in(far_0_200_0[0]), .out(far_0_200_1[0]));    relay_conn far_0_200_1_b(.in(far_0_200_0[1]), .out(far_0_200_1[1]));
    wire [1:0] far_0_200_2;    relay_conn far_0_200_2_a(.in(far_0_200_1[0]), .out(far_0_200_2[0]));    relay_conn far_0_200_2_b(.in(far_0_200_1[1]), .out(far_0_200_2[1]));
    assign layer_0[200] = far_0_200_2[0]; 
    wire [1:0] far_0_201_0;    relay_conn far_0_201_0_a(.in(in[79]), .out(far_0_201_0[0]));    relay_conn far_0_201_0_b(.in(in[137]), .out(far_0_201_0[1]));
    assign layer_0[201] = far_0_201_0[0] | far_0_201_0[1]; 
    wire [1:0] far_0_202_0;    relay_conn far_0_202_0_a(.in(in[13]), .out(far_0_202_0[0]));    relay_conn far_0_202_0_b(.in(in[109]), .out(far_0_202_0[1]));
    wire [1:0] far_0_202_1;    relay_conn far_0_202_1_a(.in(far_0_202_0[0]), .out(far_0_202_1[0]));    relay_conn far_0_202_1_b(.in(far_0_202_0[1]), .out(far_0_202_1[1]));
    wire [1:0] far_0_202_2;    relay_conn far_0_202_2_a(.in(far_0_202_1[0]), .out(far_0_202_2[0]));    relay_conn far_0_202_2_b(.in(far_0_202_1[1]), .out(far_0_202_2[1]));
    assign layer_0[202] = ~(far_0_202_2[0] | far_0_202_2[1]); 
    wire [1:0] far_0_203_0;    relay_conn far_0_203_0_a(.in(in[19]), .out(far_0_203_0[0]));    relay_conn far_0_203_0_b(.in(in[113]), .out(far_0_203_0[1]));
    wire [1:0] far_0_203_1;    relay_conn far_0_203_1_a(.in(far_0_203_0[0]), .out(far_0_203_1[0]));    relay_conn far_0_203_1_b(.in(far_0_203_0[1]), .out(far_0_203_1[1]));
    assign layer_0[203] = far_0_203_1[0] | far_0_203_1[1]; 
    wire [1:0] far_0_204_0;    relay_conn far_0_204_0_a(.in(in[136]), .out(far_0_204_0[0]));    relay_conn far_0_204_0_b(.in(in[172]), .out(far_0_204_0[1]));
    assign layer_0[204] = ~far_0_204_0[1] | (far_0_204_0[0] & far_0_204_0[1]); 
    wire [1:0] far_0_205_0;    relay_conn far_0_205_0_a(.in(in[207]), .out(far_0_205_0[0]));    relay_conn far_0_205_0_b(.in(in[151]), .out(far_0_205_0[1]));
    assign layer_0[205] = far_0_205_0[1]; 
    assign layer_0[206] = ~(in[186] ^ in[165]); 
    wire [1:0] far_0_207_0;    relay_conn far_0_207_0_a(.in(in[133]), .out(far_0_207_0[0]));    relay_conn far_0_207_0_b(.in(in[18]), .out(far_0_207_0[1]));
    wire [1:0] far_0_207_1;    relay_conn far_0_207_1_a(.in(far_0_207_0[0]), .out(far_0_207_1[0]));    relay_conn far_0_207_1_b(.in(far_0_207_0[1]), .out(far_0_207_1[1]));
    wire [1:0] far_0_207_2;    relay_conn far_0_207_2_a(.in(far_0_207_1[0]), .out(far_0_207_2[0]));    relay_conn far_0_207_2_b(.in(far_0_207_1[1]), .out(far_0_207_2[1]));
    assign layer_0[207] = far_0_207_2[0] ^ far_0_207_2[1]; 
    wire [1:0] far_0_208_0;    relay_conn far_0_208_0_a(.in(in[123]), .out(far_0_208_0[0]));    relay_conn far_0_208_0_b(.in(in[247]), .out(far_0_208_0[1]));
    wire [1:0] far_0_208_1;    relay_conn far_0_208_1_a(.in(far_0_208_0[0]), .out(far_0_208_1[0]));    relay_conn far_0_208_1_b(.in(far_0_208_0[1]), .out(far_0_208_1[1]));
    wire [1:0] far_0_208_2;    relay_conn far_0_208_2_a(.in(far_0_208_1[0]), .out(far_0_208_2[0]));    relay_conn far_0_208_2_b(.in(far_0_208_1[1]), .out(far_0_208_2[1]));
    assign layer_0[208] = ~far_0_208_2[1]; 
    assign layer_0[209] = in[188] | in[209]; 
    assign layer_0[210] = in[139]; 
    wire [1:0] far_0_211_0;    relay_conn far_0_211_0_a(.in(in[99]), .out(far_0_211_0[0]));    relay_conn far_0_211_0_b(.in(in[199]), .out(far_0_211_0[1]));
    wire [1:0] far_0_211_1;    relay_conn far_0_211_1_a(.in(far_0_211_0[0]), .out(far_0_211_1[0]));    relay_conn far_0_211_1_b(.in(far_0_211_0[1]), .out(far_0_211_1[1]));
    wire [1:0] far_0_211_2;    relay_conn far_0_211_2_a(.in(far_0_211_1[0]), .out(far_0_211_2[0]));    relay_conn far_0_211_2_b(.in(far_0_211_1[1]), .out(far_0_211_2[1]));
    assign layer_0[211] = far_0_211_2[0] & ~far_0_211_2[1]; 
    wire [1:0] far_0_212_0;    relay_conn far_0_212_0_a(.in(in[109]), .out(far_0_212_0[0]));    relay_conn far_0_212_0_b(.in(in[174]), .out(far_0_212_0[1]));
    wire [1:0] far_0_212_1;    relay_conn far_0_212_1_a(.in(far_0_212_0[0]), .out(far_0_212_1[0]));    relay_conn far_0_212_1_b(.in(far_0_212_0[1]), .out(far_0_212_1[1]));
    assign layer_0[212] = far_0_212_1[1]; 
    wire [1:0] far_0_213_0;    relay_conn far_0_213_0_a(.in(in[33]), .out(far_0_213_0[0]));    relay_conn far_0_213_0_b(.in(in[134]), .out(far_0_213_0[1]));
    wire [1:0] far_0_213_1;    relay_conn far_0_213_1_a(.in(far_0_213_0[0]), .out(far_0_213_1[0]));    relay_conn far_0_213_1_b(.in(far_0_213_0[1]), .out(far_0_213_1[1]));
    wire [1:0] far_0_213_2;    relay_conn far_0_213_2_a(.in(far_0_213_1[0]), .out(far_0_213_2[0]));    relay_conn far_0_213_2_b(.in(far_0_213_1[1]), .out(far_0_213_2[1]));
    assign layer_0[213] = far_0_213_2[0] & far_0_213_2[1]; 
    assign layer_0[214] = in[70] & ~in[53]; 
    wire [1:0] far_0_215_0;    relay_conn far_0_215_0_a(.in(in[175]), .out(far_0_215_0[0]));    relay_conn far_0_215_0_b(.in(in[79]), .out(far_0_215_0[1]));
    wire [1:0] far_0_215_1;    relay_conn far_0_215_1_a(.in(far_0_215_0[0]), .out(far_0_215_1[0]));    relay_conn far_0_215_1_b(.in(far_0_215_0[1]), .out(far_0_215_1[1]));
    wire [1:0] far_0_215_2;    relay_conn far_0_215_2_a(.in(far_0_215_1[0]), .out(far_0_215_2[0]));    relay_conn far_0_215_2_b(.in(far_0_215_1[1]), .out(far_0_215_2[1]));
    assign layer_0[215] = ~far_0_215_2[1] | (far_0_215_2[0] & far_0_215_2[1]); 
    assign layer_0[216] = ~in[99]; 
    wire [1:0] far_0_217_0;    relay_conn far_0_217_0_a(.in(in[105]), .out(far_0_217_0[0]));    relay_conn far_0_217_0_b(.in(in[182]), .out(far_0_217_0[1]));
    wire [1:0] far_0_217_1;    relay_conn far_0_217_1_a(.in(far_0_217_0[0]), .out(far_0_217_1[0]));    relay_conn far_0_217_1_b(.in(far_0_217_0[1]), .out(far_0_217_1[1]));
    assign layer_0[217] = far_0_217_1[0] & far_0_217_1[1]; 
    wire [1:0] far_0_218_0;    relay_conn far_0_218_0_a(.in(in[111]), .out(far_0_218_0[0]));    relay_conn far_0_218_0_b(.in(in[208]), .out(far_0_218_0[1]));
    wire [1:0] far_0_218_1;    relay_conn far_0_218_1_a(.in(far_0_218_0[0]), .out(far_0_218_1[0]));    relay_conn far_0_218_1_b(.in(far_0_218_0[1]), .out(far_0_218_1[1]));
    wire [1:0] far_0_218_2;    relay_conn far_0_218_2_a(.in(far_0_218_1[0]), .out(far_0_218_2[0]));    relay_conn far_0_218_2_b(.in(far_0_218_1[1]), .out(far_0_218_2[1]));
    assign layer_0[218] = far_0_218_2[0] | far_0_218_2[1]; 
    assign layer_0[219] = ~in[212] | (in[199] & in[212]); 
    wire [1:0] far_0_220_0;    relay_conn far_0_220_0_a(.in(in[167]), .out(far_0_220_0[0]));    relay_conn far_0_220_0_b(.in(in[120]), .out(far_0_220_0[1]));
    assign layer_0[220] = ~far_0_220_0[1] | (far_0_220_0[0] & far_0_220_0[1]); 
    wire [1:0] far_0_221_0;    relay_conn far_0_221_0_a(.in(in[252]), .out(far_0_221_0[0]));    relay_conn far_0_221_0_b(.in(in[210]), .out(far_0_221_0[1]));
    assign layer_0[221] = far_0_221_0[0] ^ far_0_221_0[1]; 
    assign layer_0[222] = ~(in[88] | in[112]); 
    assign layer_0[223] = ~(in[197] & in[188]); 
    wire [1:0] far_0_224_0;    relay_conn far_0_224_0_a(.in(in[18]), .out(far_0_224_0[0]));    relay_conn far_0_224_0_b(.in(in[71]), .out(far_0_224_0[1]));
    assign layer_0[224] = far_0_224_0[0] & ~far_0_224_0[1]; 
    wire [1:0] far_0_225_0;    relay_conn far_0_225_0_a(.in(in[81]), .out(far_0_225_0[0]));    relay_conn far_0_225_0_b(.in(in[172]), .out(far_0_225_0[1]));
    wire [1:0] far_0_225_1;    relay_conn far_0_225_1_a(.in(far_0_225_0[0]), .out(far_0_225_1[0]));    relay_conn far_0_225_1_b(.in(far_0_225_0[1]), .out(far_0_225_1[1]));
    assign layer_0[225] = ~far_0_225_1[1] | (far_0_225_1[0] & far_0_225_1[1]); 
    wire [1:0] far_0_226_0;    relay_conn far_0_226_0_a(.in(in[85]), .out(far_0_226_0[0]));    relay_conn far_0_226_0_b(.in(in[137]), .out(far_0_226_0[1]));
    assign layer_0[226] = far_0_226_0[0] & ~far_0_226_0[1]; 
    assign layer_0[227] = in[239]; 
    wire [1:0] far_0_228_0;    relay_conn far_0_228_0_a(.in(in[202]), .out(far_0_228_0[0]));    relay_conn far_0_228_0_b(.in(in[142]), .out(far_0_228_0[1]));
    assign layer_0[228] = ~(far_0_228_0[0] & far_0_228_0[1]); 
    assign layer_0[229] = in[139] & ~in[134]; 
    assign layer_0[230] = ~in[199]; 
    wire [1:0] far_0_231_0;    relay_conn far_0_231_0_a(.in(in[139]), .out(far_0_231_0[0]));    relay_conn far_0_231_0_b(.in(in[16]), .out(far_0_231_0[1]));
    wire [1:0] far_0_231_1;    relay_conn far_0_231_1_a(.in(far_0_231_0[0]), .out(far_0_231_1[0]));    relay_conn far_0_231_1_b(.in(far_0_231_0[1]), .out(far_0_231_1[1]));
    wire [1:0] far_0_231_2;    relay_conn far_0_231_2_a(.in(far_0_231_1[0]), .out(far_0_231_2[0]));    relay_conn far_0_231_2_b(.in(far_0_231_1[1]), .out(far_0_231_2[1]));
    assign layer_0[231] = ~far_0_231_2[1]; 
    assign layer_0[232] = in[197] & ~in[215]; 
    assign layer_0[233] = in[29] & in[31]; 
    wire [1:0] far_0_234_0;    relay_conn far_0_234_0_a(.in(in[105]), .out(far_0_234_0[0]));    relay_conn far_0_234_0_b(.in(in[157]), .out(far_0_234_0[1]));
    assign layer_0[234] = ~(far_0_234_0[0] & far_0_234_0[1]); 
    wire [1:0] far_0_235_0;    relay_conn far_0_235_0_a(.in(in[79]), .out(far_0_235_0[0]));    relay_conn far_0_235_0_b(.in(in[132]), .out(far_0_235_0[1]));
    assign layer_0[235] = far_0_235_0[0] & far_0_235_0[1]; 
    wire [1:0] far_0_236_0;    relay_conn far_0_236_0_a(.in(in[17]), .out(far_0_236_0[0]));    relay_conn far_0_236_0_b(.in(in[99]), .out(far_0_236_0[1]));
    wire [1:0] far_0_236_1;    relay_conn far_0_236_1_a(.in(far_0_236_0[0]), .out(far_0_236_1[0]));    relay_conn far_0_236_1_b(.in(far_0_236_0[1]), .out(far_0_236_1[1]));
    assign layer_0[236] = far_0_236_1[0] & ~far_0_236_1[1]; 
    wire [1:0] far_0_237_0;    relay_conn far_0_237_0_a(.in(in[159]), .out(far_0_237_0[0]));    relay_conn far_0_237_0_b(.in(in[247]), .out(far_0_237_0[1]));
    wire [1:0] far_0_237_1;    relay_conn far_0_237_1_a(.in(far_0_237_0[0]), .out(far_0_237_1[0]));    relay_conn far_0_237_1_b(.in(far_0_237_0[1]), .out(far_0_237_1[1]));
    assign layer_0[237] = far_0_237_1[0] & ~far_0_237_1[1]; 
    wire [1:0] far_0_238_0;    relay_conn far_0_238_0_a(.in(in[134]), .out(far_0_238_0[0]));    relay_conn far_0_238_0_b(.in(in[101]), .out(far_0_238_0[1]));
    assign layer_0[238] = ~far_0_238_0[1] | (far_0_238_0[0] & far_0_238_0[1]); 
    wire [1:0] far_0_239_0;    relay_conn far_0_239_0_a(.in(in[154]), .out(far_0_239_0[0]));    relay_conn far_0_239_0_b(.in(in[28]), .out(far_0_239_0[1]));
    wire [1:0] far_0_239_1;    relay_conn far_0_239_1_a(.in(far_0_239_0[0]), .out(far_0_239_1[0]));    relay_conn far_0_239_1_b(.in(far_0_239_0[1]), .out(far_0_239_1[1]));
    wire [1:0] far_0_239_2;    relay_conn far_0_239_2_a(.in(far_0_239_1[0]), .out(far_0_239_2[0]));    relay_conn far_0_239_2_b(.in(far_0_239_1[1]), .out(far_0_239_2[1]));
    assign layer_0[239] = ~(far_0_239_2[0] ^ far_0_239_2[1]); 
    wire [1:0] far_0_240_0;    relay_conn far_0_240_0_a(.in(in[207]), .out(far_0_240_0[0]));    relay_conn far_0_240_0_b(.in(in[113]), .out(far_0_240_0[1]));
    wire [1:0] far_0_240_1;    relay_conn far_0_240_1_a(.in(far_0_240_0[0]), .out(far_0_240_1[0]));    relay_conn far_0_240_1_b(.in(far_0_240_0[1]), .out(far_0_240_1[1]));
    assign layer_0[240] = far_0_240_1[0] | far_0_240_1[1]; 
    wire [1:0] far_0_241_0;    relay_conn far_0_241_0_a(.in(in[57]), .out(far_0_241_0[0]));    relay_conn far_0_241_0_b(.in(in[17]), .out(far_0_241_0[1]));
    assign layer_0[241] = ~(far_0_241_0[0] & far_0_241_0[1]); 
    assign layer_0[242] = in[164]; 
    wire [1:0] far_0_243_0;    relay_conn far_0_243_0_a(.in(in[254]), .out(far_0_243_0[0]));    relay_conn far_0_243_0_b(.in(in[197]), .out(far_0_243_0[1]));
    assign layer_0[243] = ~(far_0_243_0[0] ^ far_0_243_0[1]); 
    wire [1:0] far_0_244_0;    relay_conn far_0_244_0_a(.in(in[15]), .out(far_0_244_0[0]));    relay_conn far_0_244_0_b(.in(in[57]), .out(far_0_244_0[1]));
    assign layer_0[244] = ~far_0_244_0[1]; 
    wire [1:0] far_0_245_0;    relay_conn far_0_245_0_a(.in(in[82]), .out(far_0_245_0[0]));    relay_conn far_0_245_0_b(.in(in[172]), .out(far_0_245_0[1]));
    wire [1:0] far_0_245_1;    relay_conn far_0_245_1_a(.in(far_0_245_0[0]), .out(far_0_245_1[0]));    relay_conn far_0_245_1_b(.in(far_0_245_0[1]), .out(far_0_245_1[1]));
    assign layer_0[245] = far_0_245_1[0] & ~far_0_245_1[1]; 
    wire [1:0] far_0_246_0;    relay_conn far_0_246_0_a(.in(in[204]), .out(far_0_246_0[0]));    relay_conn far_0_246_0_b(.in(in[111]), .out(far_0_246_0[1]));
    wire [1:0] far_0_246_1;    relay_conn far_0_246_1_a(.in(far_0_246_0[0]), .out(far_0_246_1[0]));    relay_conn far_0_246_1_b(.in(far_0_246_0[1]), .out(far_0_246_1[1]));
    assign layer_0[246] = ~(far_0_246_1[0] & far_0_246_1[1]); 
    assign layer_0[247] = ~(in[87] | in[63]); 
    wire [1:0] far_0_248_0;    relay_conn far_0_248_0_a(.in(in[111]), .out(far_0_248_0[0]));    relay_conn far_0_248_0_b(.in(in[181]), .out(far_0_248_0[1]));
    wire [1:0] far_0_248_1;    relay_conn far_0_248_1_a(.in(far_0_248_0[0]), .out(far_0_248_1[0]));    relay_conn far_0_248_1_b(.in(far_0_248_0[1]), .out(far_0_248_1[1]));
    assign layer_0[248] = far_0_248_1[0]; 
    wire [1:0] far_0_249_0;    relay_conn far_0_249_0_a(.in(in[97]), .out(far_0_249_0[0]));    relay_conn far_0_249_0_b(.in(in[167]), .out(far_0_249_0[1]));
    wire [1:0] far_0_249_1;    relay_conn far_0_249_1_a(.in(far_0_249_0[0]), .out(far_0_249_1[0]));    relay_conn far_0_249_1_b(.in(far_0_249_0[1]), .out(far_0_249_1[1]));
    assign layer_0[249] = ~(far_0_249_1[0] | far_0_249_1[1]); 
    wire [1:0] far_0_250_0;    relay_conn far_0_250_0_a(.in(in[57]), .out(far_0_250_0[0]));    relay_conn far_0_250_0_b(.in(in[162]), .out(far_0_250_0[1]));
    wire [1:0] far_0_250_1;    relay_conn far_0_250_1_a(.in(far_0_250_0[0]), .out(far_0_250_1[0]));    relay_conn far_0_250_1_b(.in(far_0_250_0[1]), .out(far_0_250_1[1]));
    wire [1:0] far_0_250_2;    relay_conn far_0_250_2_a(.in(far_0_250_1[0]), .out(far_0_250_2[0]));    relay_conn far_0_250_2_b(.in(far_0_250_1[1]), .out(far_0_250_2[1]));
    assign layer_0[250] = ~(far_0_250_2[0] ^ far_0_250_2[1]); 
    assign layer_0[251] = ~in[207]; 
    wire [1:0] far_0_252_0;    relay_conn far_0_252_0_a(.in(in[57]), .out(far_0_252_0[0]));    relay_conn far_0_252_0_b(.in(in[110]), .out(far_0_252_0[1]));
    assign layer_0[252] = ~far_0_252_0[1] | (far_0_252_0[0] & far_0_252_0[1]); 
    wire [1:0] far_0_253_0;    relay_conn far_0_253_0_a(.in(in[186]), .out(far_0_253_0[0]));    relay_conn far_0_253_0_b(.in(in[140]), .out(far_0_253_0[1]));
    assign layer_0[253] = far_0_253_0[0]; 
    assign layer_0[254] = ~in[220]; 
    assign layer_0[255] = ~(in[212] & in[181]); 
    wire [1:0] far_0_256_0;    relay_conn far_0_256_0_a(.in(in[138]), .out(far_0_256_0[0]));    relay_conn far_0_256_0_b(.in(in[79]), .out(far_0_256_0[1]));
    assign layer_0[256] = far_0_256_0[0] & ~far_0_256_0[1]; 
    wire [1:0] far_0_257_0;    relay_conn far_0_257_0_a(.in(in[165]), .out(far_0_257_0[0]));    relay_conn far_0_257_0_b(.in(in[237]), .out(far_0_257_0[1]));
    wire [1:0] far_0_257_1;    relay_conn far_0_257_1_a(.in(far_0_257_0[0]), .out(far_0_257_1[0]));    relay_conn far_0_257_1_b(.in(far_0_257_0[1]), .out(far_0_257_1[1]));
    assign layer_0[257] = far_0_257_1[0] & ~far_0_257_1[1]; 
    wire [1:0] far_0_258_0;    relay_conn far_0_258_0_a(.in(in[132]), .out(far_0_258_0[0]));    relay_conn far_0_258_0_b(.in(in[164]), .out(far_0_258_0[1]));
    assign layer_0[258] = ~(far_0_258_0[0] & far_0_258_0[1]); 
    wire [1:0] far_0_259_0;    relay_conn far_0_259_0_a(.in(in[121]), .out(far_0_259_0[0]));    relay_conn far_0_259_0_b(.in(in[239]), .out(far_0_259_0[1]));
    wire [1:0] far_0_259_1;    relay_conn far_0_259_1_a(.in(far_0_259_0[0]), .out(far_0_259_1[0]));    relay_conn far_0_259_1_b(.in(far_0_259_0[1]), .out(far_0_259_1[1]));
    wire [1:0] far_0_259_2;    relay_conn far_0_259_2_a(.in(far_0_259_1[0]), .out(far_0_259_2[0]));    relay_conn far_0_259_2_b(.in(far_0_259_1[1]), .out(far_0_259_2[1]));
    assign layer_0[259] = far_0_259_2[1]; 
    assign layer_0[260] = in[216]; 
    wire [1:0] far_0_261_0;    relay_conn far_0_261_0_a(.in(in[120]), .out(far_0_261_0[0]));    relay_conn far_0_261_0_b(.in(in[28]), .out(far_0_261_0[1]));
    wire [1:0] far_0_261_1;    relay_conn far_0_261_1_a(.in(far_0_261_0[0]), .out(far_0_261_1[0]));    relay_conn far_0_261_1_b(.in(far_0_261_0[1]), .out(far_0_261_1[1]));
    assign layer_0[261] = ~(far_0_261_1[0] | far_0_261_1[1]); 
    wire [1:0] far_0_262_0;    relay_conn far_0_262_0_a(.in(in[113]), .out(far_0_262_0[0]));    relay_conn far_0_262_0_b(.in(in[162]), .out(far_0_262_0[1]));
    assign layer_0[262] = far_0_262_0[0] & ~far_0_262_0[1]; 
    assign layer_0[263] = in[30] & in[51]; 
    assign layer_0[264] = ~in[241]; 
    wire [1:0] far_0_265_0;    relay_conn far_0_265_0_a(.in(in[59]), .out(far_0_265_0[0]));    relay_conn far_0_265_0_b(.in(in[151]), .out(far_0_265_0[1]));
    wire [1:0] far_0_265_1;    relay_conn far_0_265_1_a(.in(far_0_265_0[0]), .out(far_0_265_1[0]));    relay_conn far_0_265_1_b(.in(far_0_265_0[1]), .out(far_0_265_1[1]));
    assign layer_0[265] = ~far_0_265_1[1] | (far_0_265_1[0] & far_0_265_1[1]); 
    assign layer_0[266] = ~(in[86] & in[101]); 
    wire [1:0] far_0_267_0;    relay_conn far_0_267_0_a(.in(in[158]), .out(far_0_267_0[0]));    relay_conn far_0_267_0_b(.in(in[66]), .out(far_0_267_0[1]));
    wire [1:0] far_0_267_1;    relay_conn far_0_267_1_a(.in(far_0_267_0[0]), .out(far_0_267_1[0]));    relay_conn far_0_267_1_b(.in(far_0_267_0[1]), .out(far_0_267_1[1]));
    assign layer_0[267] = ~far_0_267_1[1]; 
    wire [1:0] far_0_268_0;    relay_conn far_0_268_0_a(.in(in[177]), .out(far_0_268_0[0]));    relay_conn far_0_268_0_b(.in(in[73]), .out(far_0_268_0[1]));
    wire [1:0] far_0_268_1;    relay_conn far_0_268_1_a(.in(far_0_268_0[0]), .out(far_0_268_1[0]));    relay_conn far_0_268_1_b(.in(far_0_268_0[1]), .out(far_0_268_1[1]));
    wire [1:0] far_0_268_2;    relay_conn far_0_268_2_a(.in(far_0_268_1[0]), .out(far_0_268_2[0]));    relay_conn far_0_268_2_b(.in(far_0_268_1[1]), .out(far_0_268_2[1]));
    assign layer_0[268] = ~(far_0_268_2[0] & far_0_268_2[1]); 
    assign layer_0[269] = ~in[137] | (in[109] & in[137]); 
    wire [1:0] far_0_270_0;    relay_conn far_0_270_0_a(.in(in[15]), .out(far_0_270_0[0]));    relay_conn far_0_270_0_b(.in(in[105]), .out(far_0_270_0[1]));
    wire [1:0] far_0_270_1;    relay_conn far_0_270_1_a(.in(far_0_270_0[0]), .out(far_0_270_1[0]));    relay_conn far_0_270_1_b(.in(far_0_270_0[1]), .out(far_0_270_1[1]));
    assign layer_0[270] = ~(far_0_270_1[0] & far_0_270_1[1]); 
    wire [1:0] far_0_271_0;    relay_conn far_0_271_0_a(.in(in[66]), .out(far_0_271_0[0]));    relay_conn far_0_271_0_b(.in(in[172]), .out(far_0_271_0[1]));
    wire [1:0] far_0_271_1;    relay_conn far_0_271_1_a(.in(far_0_271_0[0]), .out(far_0_271_1[0]));    relay_conn far_0_271_1_b(.in(far_0_271_0[1]), .out(far_0_271_1[1]));
    wire [1:0] far_0_271_2;    relay_conn far_0_271_2_a(.in(far_0_271_1[0]), .out(far_0_271_2[0]));    relay_conn far_0_271_2_b(.in(far_0_271_1[1]), .out(far_0_271_2[1]));
    assign layer_0[271] = far_0_271_2[1]; 
    wire [1:0] far_0_272_0;    relay_conn far_0_272_0_a(.in(in[111]), .out(far_0_272_0[0]));    relay_conn far_0_272_0_b(.in(in[143]), .out(far_0_272_0[1]));
    assign layer_0[272] = ~(far_0_272_0[0] | far_0_272_0[1]); 
    wire [1:0] far_0_273_0;    relay_conn far_0_273_0_a(.in(in[59]), .out(far_0_273_0[0]));    relay_conn far_0_273_0_b(.in(in[18]), .out(far_0_273_0[1]));
    assign layer_0[273] = ~(far_0_273_0[0] & far_0_273_0[1]); 
    wire [1:0] far_0_274_0;    relay_conn far_0_274_0_a(.in(in[88]), .out(far_0_274_0[0]));    relay_conn far_0_274_0_b(.in(in[188]), .out(far_0_274_0[1]));
    wire [1:0] far_0_274_1;    relay_conn far_0_274_1_a(.in(far_0_274_0[0]), .out(far_0_274_1[0]));    relay_conn far_0_274_1_b(.in(far_0_274_0[1]), .out(far_0_274_1[1]));
    wire [1:0] far_0_274_2;    relay_conn far_0_274_2_a(.in(far_0_274_1[0]), .out(far_0_274_2[0]));    relay_conn far_0_274_2_b(.in(far_0_274_1[1]), .out(far_0_274_2[1]));
    assign layer_0[274] = far_0_274_2[0] ^ far_0_274_2[1]; 
    wire [1:0] far_0_275_0;    relay_conn far_0_275_0_a(.in(in[164]), .out(far_0_275_0[0]));    relay_conn far_0_275_0_b(.in(in[119]), .out(far_0_275_0[1]));
    assign layer_0[275] = ~far_0_275_0[0] | (far_0_275_0[0] & far_0_275_0[1]); 
    assign layer_0[276] = ~in[86]; 
    wire [1:0] far_0_277_0;    relay_conn far_0_277_0_a(.in(in[131]), .out(far_0_277_0[0]));    relay_conn far_0_277_0_b(.in(in[179]), .out(far_0_277_0[1]));
    assign layer_0[277] = far_0_277_0[0] & far_0_277_0[1]; 
    wire [1:0] far_0_278_0;    relay_conn far_0_278_0_a(.in(in[113]), .out(far_0_278_0[0]));    relay_conn far_0_278_0_b(.in(in[158]), .out(far_0_278_0[1]));
    assign layer_0[278] = ~far_0_278_0[0]; 
    wire [1:0] far_0_279_0;    relay_conn far_0_279_0_a(.in(in[204]), .out(far_0_279_0[0]));    relay_conn far_0_279_0_b(.in(in[97]), .out(far_0_279_0[1]));
    wire [1:0] far_0_279_1;    relay_conn far_0_279_1_a(.in(far_0_279_0[0]), .out(far_0_279_1[0]));    relay_conn far_0_279_1_b(.in(far_0_279_0[1]), .out(far_0_279_1[1]));
    wire [1:0] far_0_279_2;    relay_conn far_0_279_2_a(.in(far_0_279_1[0]), .out(far_0_279_2[0]));    relay_conn far_0_279_2_b(.in(far_0_279_1[1]), .out(far_0_279_2[1]));
    assign layer_0[279] = far_0_279_2[0] ^ far_0_279_2[1]; 
    assign layer_0[280] = ~in[132]; 
    wire [1:0] far_0_281_0;    relay_conn far_0_281_0_a(.in(in[57]), .out(far_0_281_0[0]));    relay_conn far_0_281_0_b(.in(in[174]), .out(far_0_281_0[1]));
    wire [1:0] far_0_281_1;    relay_conn far_0_281_1_a(.in(far_0_281_0[0]), .out(far_0_281_1[0]));    relay_conn far_0_281_1_b(.in(far_0_281_0[1]), .out(far_0_281_1[1]));
    wire [1:0] far_0_281_2;    relay_conn far_0_281_2_a(.in(far_0_281_1[0]), .out(far_0_281_2[0]));    relay_conn far_0_281_2_b(.in(far_0_281_1[1]), .out(far_0_281_2[1]));
    assign layer_0[281] = far_0_281_2[0] | far_0_281_2[1]; 
    assign layer_0[282] = in[113] & ~in[142]; 
    wire [1:0] far_0_283_0;    relay_conn far_0_283_0_a(.in(in[88]), .out(far_0_283_0[0]));    relay_conn far_0_283_0_b(.in(in[19]), .out(far_0_283_0[1]));
    wire [1:0] far_0_283_1;    relay_conn far_0_283_1_a(.in(far_0_283_0[0]), .out(far_0_283_1[0]));    relay_conn far_0_283_1_b(.in(far_0_283_0[1]), .out(far_0_283_1[1]));
    assign layer_0[283] = ~far_0_283_1[1]; 
    assign layer_0[284] = in[28] ^ in[56]; 
    assign layer_0[285] = in[35]; 
    wire [1:0] far_0_286_0;    relay_conn far_0_286_0_a(.in(in[211]), .out(far_0_286_0[0]));    relay_conn far_0_286_0_b(.in(in[134]), .out(far_0_286_0[1]));
    wire [1:0] far_0_286_1;    relay_conn far_0_286_1_a(.in(far_0_286_0[0]), .out(far_0_286_1[0]));    relay_conn far_0_286_1_b(.in(far_0_286_0[1]), .out(far_0_286_1[1]));
    assign layer_0[286] = ~(far_0_286_1[0] | far_0_286_1[1]); 
    wire [1:0] far_0_287_0;    relay_conn far_0_287_0_a(.in(in[239]), .out(far_0_287_0[0]));    relay_conn far_0_287_0_b(.in(in[113]), .out(far_0_287_0[1]));
    wire [1:0] far_0_287_1;    relay_conn far_0_287_1_a(.in(far_0_287_0[0]), .out(far_0_287_1[0]));    relay_conn far_0_287_1_b(.in(far_0_287_0[1]), .out(far_0_287_1[1]));
    wire [1:0] far_0_287_2;    relay_conn far_0_287_2_a(.in(far_0_287_1[0]), .out(far_0_287_2[0]));    relay_conn far_0_287_2_b(.in(far_0_287_1[1]), .out(far_0_287_2[1]));
    assign layer_0[287] = ~far_0_287_2[0] | (far_0_287_2[0] & far_0_287_2[1]); 
    assign layer_0[288] = in[234] & ~in[239]; 
    wire [1:0] far_0_289_0;    relay_conn far_0_289_0_a(.in(in[72]), .out(far_0_289_0[0]));    relay_conn far_0_289_0_b(.in(in[142]), .out(far_0_289_0[1]));
    wire [1:0] far_0_289_1;    relay_conn far_0_289_1_a(.in(far_0_289_0[0]), .out(far_0_289_1[0]));    relay_conn far_0_289_1_b(.in(far_0_289_0[1]), .out(far_0_289_1[1]));
    assign layer_0[289] = far_0_289_1[0] & far_0_289_1[1]; 
    wire [1:0] far_0_290_0;    relay_conn far_0_290_0_a(.in(in[59]), .out(far_0_290_0[0]));    relay_conn far_0_290_0_b(.in(in[0]), .out(far_0_290_0[1]));
    assign layer_0[290] = far_0_290_0[0] & far_0_290_0[1]; 
    assign layer_0[291] = in[151] | in[180]; 
    wire [1:0] far_0_292_0;    relay_conn far_0_292_0_a(.in(in[212]), .out(far_0_292_0[0]));    relay_conn far_0_292_0_b(.in(in[92]), .out(far_0_292_0[1]));
    wire [1:0] far_0_292_1;    relay_conn far_0_292_1_a(.in(far_0_292_0[0]), .out(far_0_292_1[0]));    relay_conn far_0_292_1_b(.in(far_0_292_0[1]), .out(far_0_292_1[1]));
    wire [1:0] far_0_292_2;    relay_conn far_0_292_2_a(.in(far_0_292_1[0]), .out(far_0_292_2[0]));    relay_conn far_0_292_2_b(.in(far_0_292_1[1]), .out(far_0_292_2[1]));
    assign layer_0[292] = ~far_0_292_2[0] | (far_0_292_2[0] & far_0_292_2[1]); 
    wire [1:0] far_0_293_0;    relay_conn far_0_293_0_a(.in(in[221]), .out(far_0_293_0[0]));    relay_conn far_0_293_0_b(.in(in[132]), .out(far_0_293_0[1]));
    wire [1:0] far_0_293_1;    relay_conn far_0_293_1_a(.in(far_0_293_0[0]), .out(far_0_293_1[0]));    relay_conn far_0_293_1_b(.in(far_0_293_0[1]), .out(far_0_293_1[1]));
    assign layer_0[293] = ~far_0_293_1[0]; 
    assign layer_0[294] = in[86] ^ in[70]; 
    assign layer_0[295] = in[215]; 
    wire [1:0] far_0_296_0;    relay_conn far_0_296_0_a(.in(in[113]), .out(far_0_296_0[0]));    relay_conn far_0_296_0_b(.in(in[188]), .out(far_0_296_0[1]));
    wire [1:0] far_0_296_1;    relay_conn far_0_296_1_a(.in(far_0_296_0[0]), .out(far_0_296_1[0]));    relay_conn far_0_296_1_b(.in(far_0_296_0[1]), .out(far_0_296_1[1]));
    assign layer_0[296] = far_0_296_1[0] ^ far_0_296_1[1]; 
    assign layer_0[297] = in[81]; 
    assign layer_0[298] = in[80] & in[104]; 
    wire [1:0] far_0_299_0;    relay_conn far_0_299_0_a(.in(in[48]), .out(far_0_299_0[0]));    relay_conn far_0_299_0_b(.in(in[90]), .out(far_0_299_0[1]));
    assign layer_0[299] = far_0_299_0[0] & far_0_299_0[1]; 
    wire [1:0] far_0_300_0;    relay_conn far_0_300_0_a(.in(in[104]), .out(far_0_300_0[0]));    relay_conn far_0_300_0_b(.in(in[7]), .out(far_0_300_0[1]));
    wire [1:0] far_0_300_1;    relay_conn far_0_300_1_a(.in(far_0_300_0[0]), .out(far_0_300_1[0]));    relay_conn far_0_300_1_b(.in(far_0_300_0[1]), .out(far_0_300_1[1]));
    wire [1:0] far_0_300_2;    relay_conn far_0_300_2_a(.in(far_0_300_1[0]), .out(far_0_300_2[0]));    relay_conn far_0_300_2_b(.in(far_0_300_1[1]), .out(far_0_300_2[1]));
    assign layer_0[300] = ~far_0_300_2[0] | (far_0_300_2[0] & far_0_300_2[1]); 
    wire [1:0] far_0_301_0;    relay_conn far_0_301_0_a(.in(in[189]), .out(far_0_301_0[0]));    relay_conn far_0_301_0_b(.in(in[241]), .out(far_0_301_0[1]));
    assign layer_0[301] = far_0_301_0[1]; 
    assign layer_0[302] = in[52] & ~in[81]; 
    assign layer_0[303] = in[172] & ~in[149]; 
    assign layer_0[304] = in[151] & ~in[133]; 
    wire [1:0] far_0_305_0;    relay_conn far_0_305_0_a(.in(in[36]), .out(far_0_305_0[0]));    relay_conn far_0_305_0_b(.in(in[113]), .out(far_0_305_0[1]));
    wire [1:0] far_0_305_1;    relay_conn far_0_305_1_a(.in(far_0_305_0[0]), .out(far_0_305_1[0]));    relay_conn far_0_305_1_b(.in(far_0_305_0[1]), .out(far_0_305_1[1]));
    assign layer_0[305] = far_0_305_1[0] | far_0_305_1[1]; 
    assign layer_0[306] = ~in[19]; 
    wire [1:0] far_0_307_0;    relay_conn far_0_307_0_a(.in(in[121]), .out(far_0_307_0[0]));    relay_conn far_0_307_0_b(.in(in[87]), .out(far_0_307_0[1]));
    assign layer_0[307] = far_0_307_0[0]; 
    wire [1:0] far_0_308_0;    relay_conn far_0_308_0_a(.in(in[212]), .out(far_0_308_0[0]));    relay_conn far_0_308_0_b(.in(in[175]), .out(far_0_308_0[1]));
    assign layer_0[308] = ~far_0_308_0[0] | (far_0_308_0[0] & far_0_308_0[1]); 
    wire [1:0] far_0_309_0;    relay_conn far_0_309_0_a(.in(in[55]), .out(far_0_309_0[0]));    relay_conn far_0_309_0_b(.in(in[164]), .out(far_0_309_0[1]));
    wire [1:0] far_0_309_1;    relay_conn far_0_309_1_a(.in(far_0_309_0[0]), .out(far_0_309_1[0]));    relay_conn far_0_309_1_b(.in(far_0_309_0[1]), .out(far_0_309_1[1]));
    wire [1:0] far_0_309_2;    relay_conn far_0_309_2_a(.in(far_0_309_1[0]), .out(far_0_309_2[0]));    relay_conn far_0_309_2_b(.in(far_0_309_1[1]), .out(far_0_309_2[1]));
    assign layer_0[309] = far_0_309_2[1]; 
    assign layer_0[310] = ~in[207]; 
    wire [1:0] far_0_311_0;    relay_conn far_0_311_0_a(.in(in[239]), .out(far_0_311_0[0]));    relay_conn far_0_311_0_b(.in(in[165]), .out(far_0_311_0[1]));
    wire [1:0] far_0_311_1;    relay_conn far_0_311_1_a(.in(far_0_311_0[0]), .out(far_0_311_1[0]));    relay_conn far_0_311_1_b(.in(far_0_311_0[1]), .out(far_0_311_1[1]));
    assign layer_0[311] = far_0_311_1[0] | far_0_311_1[1]; 
    assign layer_0[312] = ~in[77]; 
    wire [1:0] far_0_313_0;    relay_conn far_0_313_0_a(.in(in[57]), .out(far_0_313_0[0]));    relay_conn far_0_313_0_b(.in(in[121]), .out(far_0_313_0[1]));
    wire [1:0] far_0_313_1;    relay_conn far_0_313_1_a(.in(far_0_313_0[0]), .out(far_0_313_1[0]));    relay_conn far_0_313_1_b(.in(far_0_313_0[1]), .out(far_0_313_1[1]));
    assign layer_0[313] = far_0_313_1[0] | far_0_313_1[1]; 
    assign layer_0[314] = ~in[173]; 
    wire [1:0] far_0_315_0;    relay_conn far_0_315_0_a(.in(in[32]), .out(far_0_315_0[0]));    relay_conn far_0_315_0_b(.in(in[76]), .out(far_0_315_0[1]));
    assign layer_0[315] = ~far_0_315_0[0] | (far_0_315_0[0] & far_0_315_0[1]); 
    wire [1:0] far_0_316_0;    relay_conn far_0_316_0_a(.in(in[89]), .out(far_0_316_0[0]));    relay_conn far_0_316_0_b(.in(in[48]), .out(far_0_316_0[1]));
    assign layer_0[316] = far_0_316_0[1] & ~far_0_316_0[0]; 
    assign layer_0[317] = in[158] ^ in[187]; 
    wire [1:0] far_0_318_0;    relay_conn far_0_318_0_a(.in(in[94]), .out(far_0_318_0[0]));    relay_conn far_0_318_0_b(.in(in[136]), .out(far_0_318_0[1]));
    assign layer_0[318] = ~(far_0_318_0[0] & far_0_318_0[1]); 
    assign layer_0[319] = ~(in[49] & in[36]); 
    assign layer_0[320] = ~(in[98] ^ in[99]); 
    wire [1:0] far_0_321_0;    relay_conn far_0_321_0_a(.in(in[163]), .out(far_0_321_0[0]));    relay_conn far_0_321_0_b(.in(in[43]), .out(far_0_321_0[1]));
    wire [1:0] far_0_321_1;    relay_conn far_0_321_1_a(.in(far_0_321_0[0]), .out(far_0_321_1[0]));    relay_conn far_0_321_1_b(.in(far_0_321_0[1]), .out(far_0_321_1[1]));
    wire [1:0] far_0_321_2;    relay_conn far_0_321_2_a(.in(far_0_321_1[0]), .out(far_0_321_2[0]));    relay_conn far_0_321_2_b(.in(far_0_321_1[1]), .out(far_0_321_2[1]));
    assign layer_0[321] = far_0_321_2[0] | far_0_321_2[1]; 
    assign layer_0[322] = in[199] & ~in[181]; 
    wire [1:0] far_0_323_0;    relay_conn far_0_323_0_a(.in(in[10]), .out(far_0_323_0[0]));    relay_conn far_0_323_0_b(.in(in[127]), .out(far_0_323_0[1]));
    wire [1:0] far_0_323_1;    relay_conn far_0_323_1_a(.in(far_0_323_0[0]), .out(far_0_323_1[0]));    relay_conn far_0_323_1_b(.in(far_0_323_0[1]), .out(far_0_323_1[1]));
    wire [1:0] far_0_323_2;    relay_conn far_0_323_2_a(.in(far_0_323_1[0]), .out(far_0_323_2[0]));    relay_conn far_0_323_2_b(.in(far_0_323_1[1]), .out(far_0_323_2[1]));
    assign layer_0[323] = ~(far_0_323_2[0] | far_0_323_2[1]); 
    wire [1:0] far_0_324_0;    relay_conn far_0_324_0_a(.in(in[213]), .out(far_0_324_0[0]));    relay_conn far_0_324_0_b(.in(in[132]), .out(far_0_324_0[1]));
    wire [1:0] far_0_324_1;    relay_conn far_0_324_1_a(.in(far_0_324_0[0]), .out(far_0_324_1[0]));    relay_conn far_0_324_1_b(.in(far_0_324_0[1]), .out(far_0_324_1[1]));
    assign layer_0[324] = ~(far_0_324_1[0] & far_0_324_1[1]); 
    wire [1:0] far_0_325_0;    relay_conn far_0_325_0_a(.in(in[117]), .out(far_0_325_0[0]));    relay_conn far_0_325_0_b(.in(in[164]), .out(far_0_325_0[1]));
    assign layer_0[325] = ~(far_0_325_0[0] | far_0_325_0[1]); 
    wire [1:0] far_0_326_0;    relay_conn far_0_326_0_a(.in(in[241]), .out(far_0_326_0[0]));    relay_conn far_0_326_0_b(.in(in[122]), .out(far_0_326_0[1]));
    wire [1:0] far_0_326_1;    relay_conn far_0_326_1_a(.in(far_0_326_0[0]), .out(far_0_326_1[0]));    relay_conn far_0_326_1_b(.in(far_0_326_0[1]), .out(far_0_326_1[1]));
    wire [1:0] far_0_326_2;    relay_conn far_0_326_2_a(.in(far_0_326_1[0]), .out(far_0_326_2[0]));    relay_conn far_0_326_2_b(.in(far_0_326_1[1]), .out(far_0_326_2[1]));
    assign layer_0[326] = ~far_0_326_2[0] | (far_0_326_2[0] & far_0_326_2[1]); 
    wire [1:0] far_0_327_0;    relay_conn far_0_327_0_a(.in(in[109]), .out(far_0_327_0[0]));    relay_conn far_0_327_0_b(.in(in[187]), .out(far_0_327_0[1]));
    wire [1:0] far_0_327_1;    relay_conn far_0_327_1_a(.in(far_0_327_0[0]), .out(far_0_327_1[0]));    relay_conn far_0_327_1_b(.in(far_0_327_0[1]), .out(far_0_327_1[1]));
    assign layer_0[327] = ~(far_0_327_1[0] | far_0_327_1[1]); 
    wire [1:0] far_0_328_0;    relay_conn far_0_328_0_a(.in(in[121]), .out(far_0_328_0[0]));    relay_conn far_0_328_0_b(.in(in[157]), .out(far_0_328_0[1]));
    assign layer_0[328] = far_0_328_0[0] & far_0_328_0[1]; 
    assign layer_0[329] = ~(in[187] | in[164]); 
    assign layer_0[330] = ~in[122]; 
    wire [1:0] far_0_331_0;    relay_conn far_0_331_0_a(.in(in[20]), .out(far_0_331_0[0]));    relay_conn far_0_331_0_b(.in(in[66]), .out(far_0_331_0[1]));
    assign layer_0[331] = ~(far_0_331_0[0] ^ far_0_331_0[1]); 
    assign layer_0[332] = ~(in[188] & in[212]); 
    assign layer_0[333] = ~(in[157] | in[150]); 
    wire [1:0] far_0_334_0;    relay_conn far_0_334_0_a(.in(in[190]), .out(far_0_334_0[0]));    relay_conn far_0_334_0_b(.in(in[117]), .out(far_0_334_0[1]));
    wire [1:0] far_0_334_1;    relay_conn far_0_334_1_a(.in(far_0_334_0[0]), .out(far_0_334_1[0]));    relay_conn far_0_334_1_b(.in(far_0_334_0[1]), .out(far_0_334_1[1]));
    assign layer_0[334] = ~far_0_334_1[0] | (far_0_334_1[0] & far_0_334_1[1]); 
    wire [1:0] far_0_335_0;    relay_conn far_0_335_0_a(.in(in[121]), .out(far_0_335_0[0]));    relay_conn far_0_335_0_b(.in(in[59]), .out(far_0_335_0[1]));
    assign layer_0[335] = ~(far_0_335_0[0] | far_0_335_0[1]); 
    assign layer_0[336] = ~(in[172] | in[170]); 
    wire [1:0] far_0_337_0;    relay_conn far_0_337_0_a(.in(in[186]), .out(far_0_337_0[0]));    relay_conn far_0_337_0_b(.in(in[226]), .out(far_0_337_0[1]));
    assign layer_0[337] = far_0_337_0[1]; 
    assign layer_0[338] = ~in[212] | (in[212] & in[239]); 
    wire [1:0] far_0_339_0;    relay_conn far_0_339_0_a(.in(in[117]), .out(far_0_339_0[0]));    relay_conn far_0_339_0_b(.in(in[233]), .out(far_0_339_0[1]));
    wire [1:0] far_0_339_1;    relay_conn far_0_339_1_a(.in(far_0_339_0[0]), .out(far_0_339_1[0]));    relay_conn far_0_339_1_b(.in(far_0_339_0[1]), .out(far_0_339_1[1]));
    wire [1:0] far_0_339_2;    relay_conn far_0_339_2_a(.in(far_0_339_1[0]), .out(far_0_339_2[0]));    relay_conn far_0_339_2_b(.in(far_0_339_1[1]), .out(far_0_339_2[1]));
    assign layer_0[339] = ~far_0_339_2[0]; 
    wire [1:0] far_0_340_0;    relay_conn far_0_340_0_a(.in(in[40]), .out(far_0_340_0[0]));    relay_conn far_0_340_0_b(.in(in[88]), .out(far_0_340_0[1]));
    assign layer_0[340] = ~(far_0_340_0[0] | far_0_340_0[1]); 
    wire [1:0] far_0_341_0;    relay_conn far_0_341_0_a(.in(in[132]), .out(far_0_341_0[0]));    relay_conn far_0_341_0_b(.in(in[225]), .out(far_0_341_0[1]));
    wire [1:0] far_0_341_1;    relay_conn far_0_341_1_a(.in(far_0_341_0[0]), .out(far_0_341_1[0]));    relay_conn far_0_341_1_b(.in(far_0_341_0[1]), .out(far_0_341_1[1]));
    assign layer_0[341] = far_0_341_1[0] & far_0_341_1[1]; 
    assign layer_0[342] = in[179] | in[156]; 
    wire [1:0] far_0_343_0;    relay_conn far_0_343_0_a(.in(in[207]), .out(far_0_343_0[0]));    relay_conn far_0_343_0_b(.in(in[151]), .out(far_0_343_0[1]));
    assign layer_0[343] = far_0_343_0[1]; 
    wire [1:0] far_0_344_0;    relay_conn far_0_344_0_a(.in(in[151]), .out(far_0_344_0[0]));    relay_conn far_0_344_0_b(.in(in[212]), .out(far_0_344_0[1]));
    assign layer_0[344] = ~(far_0_344_0[0] | far_0_344_0[1]); 
    assign layer_0[345] = ~(in[87] | in[79]); 
    assign layer_0[346] = ~(in[188] & in[211]); 
    assign layer_0[347] = ~(in[22] | in[28]); 
    wire [1:0] far_0_348_0;    relay_conn far_0_348_0_a(.in(in[37]), .out(far_0_348_0[0]));    relay_conn far_0_348_0_b(.in(in[72]), .out(far_0_348_0[1]));
    assign layer_0[348] = far_0_348_0[1] & ~far_0_348_0[0]; 
    wire [1:0] far_0_349_0;    relay_conn far_0_349_0_a(.in(in[82]), .out(far_0_349_0[0]));    relay_conn far_0_349_0_b(.in(in[127]), .out(far_0_349_0[1]));
    assign layer_0[349] = ~far_0_349_0[0] | (far_0_349_0[0] & far_0_349_0[1]); 
    wire [1:0] far_0_350_0;    relay_conn far_0_350_0_a(.in(in[113]), .out(far_0_350_0[0]));    relay_conn far_0_350_0_b(.in(in[172]), .out(far_0_350_0[1]));
    assign layer_0[350] = ~far_0_350_0[0]; 
    wire [1:0] far_0_351_0;    relay_conn far_0_351_0_a(.in(in[210]), .out(far_0_351_0[0]));    relay_conn far_0_351_0_b(.in(in[84]), .out(far_0_351_0[1]));
    wire [1:0] far_0_351_1;    relay_conn far_0_351_1_a(.in(far_0_351_0[0]), .out(far_0_351_1[0]));    relay_conn far_0_351_1_b(.in(far_0_351_0[1]), .out(far_0_351_1[1]));
    wire [1:0] far_0_351_2;    relay_conn far_0_351_2_a(.in(far_0_351_1[0]), .out(far_0_351_2[0]));    relay_conn far_0_351_2_b(.in(far_0_351_1[1]), .out(far_0_351_2[1]));
    assign layer_0[351] = ~(far_0_351_2[0] & far_0_351_2[1]); 
    wire [1:0] far_0_352_0;    relay_conn far_0_352_0_a(.in(in[181]), .out(far_0_352_0[0]));    relay_conn far_0_352_0_b(.in(in[61]), .out(far_0_352_0[1]));
    wire [1:0] far_0_352_1;    relay_conn far_0_352_1_a(.in(far_0_352_0[0]), .out(far_0_352_1[0]));    relay_conn far_0_352_1_b(.in(far_0_352_0[1]), .out(far_0_352_1[1]));
    wire [1:0] far_0_352_2;    relay_conn far_0_352_2_a(.in(far_0_352_1[0]), .out(far_0_352_2[0]));    relay_conn far_0_352_2_b(.in(far_0_352_1[1]), .out(far_0_352_2[1]));
    assign layer_0[352] = far_0_352_2[1] & ~far_0_352_2[0]; 
    wire [1:0] far_0_353_0;    relay_conn far_0_353_0_a(.in(in[229]), .out(far_0_353_0[0]));    relay_conn far_0_353_0_b(.in(in[181]), .out(far_0_353_0[1]));
    assign layer_0[353] = ~far_0_353_0[1]; 
    assign layer_0[354] = ~in[17]; 
    wire [1:0] far_0_355_0;    relay_conn far_0_355_0_a(.in(in[165]), .out(far_0_355_0[0]));    relay_conn far_0_355_0_b(.in(in[84]), .out(far_0_355_0[1]));
    wire [1:0] far_0_355_1;    relay_conn far_0_355_1_a(.in(far_0_355_0[0]), .out(far_0_355_1[0]));    relay_conn far_0_355_1_b(.in(far_0_355_0[1]), .out(far_0_355_1[1]));
    assign layer_0[355] = ~far_0_355_1[1] | (far_0_355_1[0] & far_0_355_1[1]); 
    wire [1:0] far_0_356_0;    relay_conn far_0_356_0_a(.in(in[211]), .out(far_0_356_0[0]));    relay_conn far_0_356_0_b(.in(in[149]), .out(far_0_356_0[1]));
    assign layer_0[356] = ~far_0_356_0[1] | (far_0_356_0[0] & far_0_356_0[1]); 
    wire [1:0] far_0_357_0;    relay_conn far_0_357_0_a(.in(in[151]), .out(far_0_357_0[0]));    relay_conn far_0_357_0_b(.in(in[110]), .out(far_0_357_0[1]));
    assign layer_0[357] = ~far_0_357_0[0] | (far_0_357_0[0] & far_0_357_0[1]); 
    wire [1:0] far_0_358_0;    relay_conn far_0_358_0_a(.in(in[175]), .out(far_0_358_0[0]));    relay_conn far_0_358_0_b(.in(in[82]), .out(far_0_358_0[1]));
    wire [1:0] far_0_358_1;    relay_conn far_0_358_1_a(.in(far_0_358_0[0]), .out(far_0_358_1[0]));    relay_conn far_0_358_1_b(.in(far_0_358_0[1]), .out(far_0_358_1[1]));
    assign layer_0[358] = ~far_0_358_1[0] | (far_0_358_1[0] & far_0_358_1[1]); 
    wire [1:0] far_0_359_0;    relay_conn far_0_359_0_a(.in(in[150]), .out(far_0_359_0[0]));    relay_conn far_0_359_0_b(.in(in[213]), .out(far_0_359_0[1]));
    assign layer_0[359] = ~far_0_359_0[0] | (far_0_359_0[0] & far_0_359_0[1]); 
    wire [1:0] far_0_360_0;    relay_conn far_0_360_0_a(.in(in[88]), .out(far_0_360_0[0]));    relay_conn far_0_360_0_b(.in(in[215]), .out(far_0_360_0[1]));
    wire [1:0] far_0_360_1;    relay_conn far_0_360_1_a(.in(far_0_360_0[0]), .out(far_0_360_1[0]));    relay_conn far_0_360_1_b(.in(far_0_360_0[1]), .out(far_0_360_1[1]));
    wire [1:0] far_0_360_2;    relay_conn far_0_360_2_a(.in(far_0_360_1[0]), .out(far_0_360_2[0]));    relay_conn far_0_360_2_b(.in(far_0_360_1[1]), .out(far_0_360_2[1]));
    assign layer_0[360] = far_0_360_2[0] | far_0_360_2[1]; 
    wire [1:0] far_0_361_0;    relay_conn far_0_361_0_a(.in(in[53]), .out(far_0_361_0[0]));    relay_conn far_0_361_0_b(.in(in[136]), .out(far_0_361_0[1]));
    wire [1:0] far_0_361_1;    relay_conn far_0_361_1_a(.in(far_0_361_0[0]), .out(far_0_361_1[0]));    relay_conn far_0_361_1_b(.in(far_0_361_0[1]), .out(far_0_361_1[1]));
    assign layer_0[361] = far_0_361_1[1]; 
    assign layer_0[362] = ~in[138]; 
    wire [1:0] far_0_363_0;    relay_conn far_0_363_0_a(.in(in[137]), .out(far_0_363_0[0]));    relay_conn far_0_363_0_b(.in(in[25]), .out(far_0_363_0[1]));
    wire [1:0] far_0_363_1;    relay_conn far_0_363_1_a(.in(far_0_363_0[0]), .out(far_0_363_1[0]));    relay_conn far_0_363_1_b(.in(far_0_363_0[1]), .out(far_0_363_1[1]));
    wire [1:0] far_0_363_2;    relay_conn far_0_363_2_a(.in(far_0_363_1[0]), .out(far_0_363_2[0]));    relay_conn far_0_363_2_b(.in(far_0_363_1[1]), .out(far_0_363_2[1]));
    assign layer_0[363] = far_0_363_2[0] ^ far_0_363_2[1]; 
    wire [1:0] far_0_364_0;    relay_conn far_0_364_0_a(.in(in[199]), .out(far_0_364_0[0]));    relay_conn far_0_364_0_b(.in(in[249]), .out(far_0_364_0[1]));
    assign layer_0[364] = far_0_364_0[1]; 
    wire [1:0] far_0_365_0;    relay_conn far_0_365_0_a(.in(in[215]), .out(far_0_365_0[0]));    relay_conn far_0_365_0_b(.in(in[110]), .out(far_0_365_0[1]));
    wire [1:0] far_0_365_1;    relay_conn far_0_365_1_a(.in(far_0_365_0[0]), .out(far_0_365_1[0]));    relay_conn far_0_365_1_b(.in(far_0_365_0[1]), .out(far_0_365_1[1]));
    wire [1:0] far_0_365_2;    relay_conn far_0_365_2_a(.in(far_0_365_1[0]), .out(far_0_365_2[0]));    relay_conn far_0_365_2_b(.in(far_0_365_1[1]), .out(far_0_365_2[1]));
    assign layer_0[365] = far_0_365_2[0]; 
    assign layer_0[366] = in[65]; 
    wire [1:0] far_0_367_0;    relay_conn far_0_367_0_a(.in(in[121]), .out(far_0_367_0[0]));    relay_conn far_0_367_0_b(.in(in[75]), .out(far_0_367_0[1]));
    assign layer_0[367] = far_0_367_0[0]; 
    wire [1:0] far_0_368_0;    relay_conn far_0_368_0_a(.in(in[125]), .out(far_0_368_0[0]));    relay_conn far_0_368_0_b(.in(in[164]), .out(far_0_368_0[1]));
    assign layer_0[368] = ~(far_0_368_0[0] ^ far_0_368_0[1]); 
    assign layer_0[369] = in[221] & ~in[223]; 
    assign layer_0[370] = in[189] & in[197]; 
    wire [1:0] far_0_371_0;    relay_conn far_0_371_0_a(.in(in[150]), .out(far_0_371_0[0]));    relay_conn far_0_371_0_b(.in(in[109]), .out(far_0_371_0[1]));
    assign layer_0[371] = ~(far_0_371_0[0] & far_0_371_0[1]); 
    assign layer_0[372] = in[212] ^ in[241]; 
    wire [1:0] far_0_373_0;    relay_conn far_0_373_0_a(.in(in[196]), .out(far_0_373_0[0]));    relay_conn far_0_373_0_b(.in(in[239]), .out(far_0_373_0[1]));
    assign layer_0[373] = ~(far_0_373_0[0] & far_0_373_0[1]); 
    wire [1:0] far_0_374_0;    relay_conn far_0_374_0_a(.in(in[121]), .out(far_0_374_0[0]));    relay_conn far_0_374_0_b(.in(in[49]), .out(far_0_374_0[1]));
    wire [1:0] far_0_374_1;    relay_conn far_0_374_1_a(.in(far_0_374_0[0]), .out(far_0_374_1[0]));    relay_conn far_0_374_1_b(.in(far_0_374_0[1]), .out(far_0_374_1[1]));
    assign layer_0[374] = far_0_374_1[1]; 
    assign layer_0[375] = ~in[237] | (in[237] & in[251]); 
    assign layer_0[376] = in[164] & in[151]; 
    wire [1:0] far_0_377_0;    relay_conn far_0_377_0_a(.in(in[202]), .out(far_0_377_0[0]));    relay_conn far_0_377_0_b(.in(in[109]), .out(far_0_377_0[1]));
    wire [1:0] far_0_377_1;    relay_conn far_0_377_1_a(.in(far_0_377_0[0]), .out(far_0_377_1[0]));    relay_conn far_0_377_1_b(.in(far_0_377_0[1]), .out(far_0_377_1[1]));
    assign layer_0[377] = far_0_377_1[1]; 
    wire [1:0] far_0_378_0;    relay_conn far_0_378_0_a(.in(in[25]), .out(far_0_378_0[0]));    relay_conn far_0_378_0_b(.in(in[87]), .out(far_0_378_0[1]));
    assign layer_0[378] = ~(far_0_378_0[0] | far_0_378_0[1]); 
    wire [1:0] far_0_379_0;    relay_conn far_0_379_0_a(.in(in[112]), .out(far_0_379_0[0]));    relay_conn far_0_379_0_b(.in(in[65]), .out(far_0_379_0[1]));
    assign layer_0[379] = ~(far_0_379_0[0] & far_0_379_0[1]); 
    wire [1:0] far_0_380_0;    relay_conn far_0_380_0_a(.in(in[136]), .out(far_0_380_0[0]));    relay_conn far_0_380_0_b(.in(in[20]), .out(far_0_380_0[1]));
    wire [1:0] far_0_380_1;    relay_conn far_0_380_1_a(.in(far_0_380_0[0]), .out(far_0_380_1[0]));    relay_conn far_0_380_1_b(.in(far_0_380_0[1]), .out(far_0_380_1[1]));
    wire [1:0] far_0_380_2;    relay_conn far_0_380_2_a(.in(far_0_380_1[0]), .out(far_0_380_2[0]));    relay_conn far_0_380_2_b(.in(far_0_380_1[1]), .out(far_0_380_2[1]));
    assign layer_0[380] = far_0_380_2[0] | far_0_380_2[1]; 
    wire [1:0] far_0_381_0;    relay_conn far_0_381_0_a(.in(in[57]), .out(far_0_381_0[0]));    relay_conn far_0_381_0_b(.in(in[17]), .out(far_0_381_0[1]));
    assign layer_0[381] = ~far_0_381_0[1] | (far_0_381_0[0] & far_0_381_0[1]); 
    wire [1:0] far_0_382_0;    relay_conn far_0_382_0_a(.in(in[102]), .out(far_0_382_0[0]));    relay_conn far_0_382_0_b(.in(in[203]), .out(far_0_382_0[1]));
    wire [1:0] far_0_382_1;    relay_conn far_0_382_1_a(.in(far_0_382_0[0]), .out(far_0_382_1[0]));    relay_conn far_0_382_1_b(.in(far_0_382_0[1]), .out(far_0_382_1[1]));
    wire [1:0] far_0_382_2;    relay_conn far_0_382_2_a(.in(far_0_382_1[0]), .out(far_0_382_2[0]));    relay_conn far_0_382_2_b(.in(far_0_382_1[1]), .out(far_0_382_2[1]));
    assign layer_0[382] = far_0_382_2[0]; 
    assign layer_0[383] = in[51] | in[22]; 
    wire [1:0] far_0_384_0;    relay_conn far_0_384_0_a(.in(in[181]), .out(far_0_384_0[0]));    relay_conn far_0_384_0_b(.in(in[117]), .out(far_0_384_0[1]));
    wire [1:0] far_0_384_1;    relay_conn far_0_384_1_a(.in(far_0_384_0[0]), .out(far_0_384_1[0]));    relay_conn far_0_384_1_b(.in(far_0_384_0[1]), .out(far_0_384_1[1]));
    assign layer_0[384] = far_0_384_1[0] | far_0_384_1[1]; 
    wire [1:0] far_0_385_0;    relay_conn far_0_385_0_a(.in(in[0]), .out(far_0_385_0[0]));    relay_conn far_0_385_0_b(.in(in[98]), .out(far_0_385_0[1]));
    wire [1:0] far_0_385_1;    relay_conn far_0_385_1_a(.in(far_0_385_0[0]), .out(far_0_385_1[0]));    relay_conn far_0_385_1_b(.in(far_0_385_0[1]), .out(far_0_385_1[1]));
    wire [1:0] far_0_385_2;    relay_conn far_0_385_2_a(.in(far_0_385_1[0]), .out(far_0_385_2[0]));    relay_conn far_0_385_2_b(.in(far_0_385_1[1]), .out(far_0_385_2[1]));
    assign layer_0[385] = ~(far_0_385_2[0] ^ far_0_385_2[1]); 
    wire [1:0] far_0_386_0;    relay_conn far_0_386_0_a(.in(in[104]), .out(far_0_386_0[0]));    relay_conn far_0_386_0_b(.in(in[57]), .out(far_0_386_0[1]));
    assign layer_0[386] = ~far_0_386_0[0]; 
    wire [1:0] far_0_387_0;    relay_conn far_0_387_0_a(.in(in[150]), .out(far_0_387_0[0]));    relay_conn far_0_387_0_b(.in(in[199]), .out(far_0_387_0[1]));
    assign layer_0[387] = far_0_387_0[1] & ~far_0_387_0[0]; 
    wire [1:0] far_0_388_0;    relay_conn far_0_388_0_a(.in(in[255]), .out(far_0_388_0[0]));    relay_conn far_0_388_0_b(.in(in[185]), .out(far_0_388_0[1]));
    wire [1:0] far_0_388_1;    relay_conn far_0_388_1_a(.in(far_0_388_0[0]), .out(far_0_388_1[0]));    relay_conn far_0_388_1_b(.in(far_0_388_0[1]), .out(far_0_388_1[1]));
    assign layer_0[388] = far_0_388_1[1]; 
    wire [1:0] far_0_389_0;    relay_conn far_0_389_0_a(.in(in[72]), .out(far_0_389_0[0]));    relay_conn far_0_389_0_b(.in(in[157]), .out(far_0_389_0[1]));
    wire [1:0] far_0_389_1;    relay_conn far_0_389_1_a(.in(far_0_389_0[0]), .out(far_0_389_1[0]));    relay_conn far_0_389_1_b(.in(far_0_389_0[1]), .out(far_0_389_1[1]));
    assign layer_0[389] = ~far_0_389_1[0] | (far_0_389_1[0] & far_0_389_1[1]); 
    wire [1:0] far_0_390_0;    relay_conn far_0_390_0_a(.in(in[37]), .out(far_0_390_0[0]));    relay_conn far_0_390_0_b(.in(in[164]), .out(far_0_390_0[1]));
    wire [1:0] far_0_390_1;    relay_conn far_0_390_1_a(.in(far_0_390_0[0]), .out(far_0_390_1[0]));    relay_conn far_0_390_1_b(.in(far_0_390_0[1]), .out(far_0_390_1[1]));
    wire [1:0] far_0_390_2;    relay_conn far_0_390_2_a(.in(far_0_390_1[0]), .out(far_0_390_2[0]));    relay_conn far_0_390_2_b(.in(far_0_390_1[1]), .out(far_0_390_2[1]));
    assign layer_0[390] = ~far_0_390_2[0] | (far_0_390_2[0] & far_0_390_2[1]); 
    wire [1:0] far_0_391_0;    relay_conn far_0_391_0_a(.in(in[68]), .out(far_0_391_0[0]));    relay_conn far_0_391_0_b(.in(in[121]), .out(far_0_391_0[1]));
    assign layer_0[391] = ~far_0_391_0[1] | (far_0_391_0[0] & far_0_391_0[1]); 
    wire [1:0] far_0_392_0;    relay_conn far_0_392_0_a(.in(in[130]), .out(far_0_392_0[0]));    relay_conn far_0_392_0_b(.in(in[196]), .out(far_0_392_0[1]));
    wire [1:0] far_0_392_1;    relay_conn far_0_392_1_a(.in(far_0_392_0[0]), .out(far_0_392_1[0]));    relay_conn far_0_392_1_b(.in(far_0_392_0[1]), .out(far_0_392_1[1]));
    assign layer_0[392] = ~(far_0_392_1[0] & far_0_392_1[1]); 
    wire [1:0] far_0_393_0;    relay_conn far_0_393_0_a(.in(in[99]), .out(far_0_393_0[0]));    relay_conn far_0_393_0_b(.in(in[153]), .out(far_0_393_0[1]));
    assign layer_0[393] = far_0_393_0[0] | far_0_393_0[1]; 
    wire [1:0] far_0_394_0;    relay_conn far_0_394_0_a(.in(in[57]), .out(far_0_394_0[0]));    relay_conn far_0_394_0_b(.in(in[125]), .out(far_0_394_0[1]));
    wire [1:0] far_0_394_1;    relay_conn far_0_394_1_a(.in(far_0_394_0[0]), .out(far_0_394_1[0]));    relay_conn far_0_394_1_b(.in(far_0_394_0[1]), .out(far_0_394_1[1]));
    assign layer_0[394] = ~(far_0_394_1[0] ^ far_0_394_1[1]); 
    assign layer_0[395] = ~(in[128] | in[119]); 
    wire [1:0] far_0_396_0;    relay_conn far_0_396_0_a(.in(in[174]), .out(far_0_396_0[0]));    relay_conn far_0_396_0_b(.in(in[133]), .out(far_0_396_0[1]));
    assign layer_0[396] = far_0_396_0[0] | far_0_396_0[1]; 
    wire [1:0] far_0_397_0;    relay_conn far_0_397_0_a(.in(in[241]), .out(far_0_397_0[0]));    relay_conn far_0_397_0_b(.in(in[132]), .out(far_0_397_0[1]));
    wire [1:0] far_0_397_1;    relay_conn far_0_397_1_a(.in(far_0_397_0[0]), .out(far_0_397_1[0]));    relay_conn far_0_397_1_b(.in(far_0_397_0[1]), .out(far_0_397_1[1]));
    wire [1:0] far_0_397_2;    relay_conn far_0_397_2_a(.in(far_0_397_1[0]), .out(far_0_397_2[0]));    relay_conn far_0_397_2_b(.in(far_0_397_1[1]), .out(far_0_397_2[1]));
    assign layer_0[397] = far_0_397_2[0] & far_0_397_2[1]; 
    wire [1:0] far_0_398_0;    relay_conn far_0_398_0_a(.in(in[164]), .out(far_0_398_0[0]));    relay_conn far_0_398_0_b(.in(in[93]), .out(far_0_398_0[1]));
    wire [1:0] far_0_398_1;    relay_conn far_0_398_1_a(.in(far_0_398_0[0]), .out(far_0_398_1[0]));    relay_conn far_0_398_1_b(.in(far_0_398_0[1]), .out(far_0_398_1[1]));
    assign layer_0[398] = ~(far_0_398_1[0] & far_0_398_1[1]); 
    wire [1:0] far_0_399_0;    relay_conn far_0_399_0_a(.in(in[167]), .out(far_0_399_0[0]));    relay_conn far_0_399_0_b(.in(in[72]), .out(far_0_399_0[1]));
    wire [1:0] far_0_399_1;    relay_conn far_0_399_1_a(.in(far_0_399_0[0]), .out(far_0_399_1[0]));    relay_conn far_0_399_1_b(.in(far_0_399_0[1]), .out(far_0_399_1[1]));
    assign layer_0[399] = far_0_399_1[0] | far_0_399_1[1]; 
    assign layer_0[400] = ~in[133]; 
    wire [1:0] far_0_401_0;    relay_conn far_0_401_0_a(.in(in[249]), .out(far_0_401_0[0]));    relay_conn far_0_401_0_b(.in(in[207]), .out(far_0_401_0[1]));
    assign layer_0[401] = ~(far_0_401_0[0] ^ far_0_401_0[1]); 
    wire [1:0] far_0_402_0;    relay_conn far_0_402_0_a(.in(in[199]), .out(far_0_402_0[0]));    relay_conn far_0_402_0_b(.in(in[72]), .out(far_0_402_0[1]));
    wire [1:0] far_0_402_1;    relay_conn far_0_402_1_a(.in(far_0_402_0[0]), .out(far_0_402_1[0]));    relay_conn far_0_402_1_b(.in(far_0_402_0[1]), .out(far_0_402_1[1]));
    wire [1:0] far_0_402_2;    relay_conn far_0_402_2_a(.in(far_0_402_1[0]), .out(far_0_402_2[0]));    relay_conn far_0_402_2_b(.in(far_0_402_1[1]), .out(far_0_402_2[1]));
    assign layer_0[402] = far_0_402_2[1] & ~far_0_402_2[0]; 
    wire [1:0] far_0_403_0;    relay_conn far_0_403_0_a(.in(in[57]), .out(far_0_403_0[0]));    relay_conn far_0_403_0_b(.in(in[3]), .out(far_0_403_0[1]));
    assign layer_0[403] = far_0_403_0[1] & ~far_0_403_0[0]; 
    assign layer_0[404] = in[151] & in[122]; 
    wire [1:0] far_0_405_0;    relay_conn far_0_405_0_a(.in(in[67]), .out(far_0_405_0[0]));    relay_conn far_0_405_0_b(.in(in[170]), .out(far_0_405_0[1]));
    wire [1:0] far_0_405_1;    relay_conn far_0_405_1_a(.in(far_0_405_0[0]), .out(far_0_405_1[0]));    relay_conn far_0_405_1_b(.in(far_0_405_0[1]), .out(far_0_405_1[1]));
    wire [1:0] far_0_405_2;    relay_conn far_0_405_2_a(.in(far_0_405_1[0]), .out(far_0_405_2[0]));    relay_conn far_0_405_2_b(.in(far_0_405_1[1]), .out(far_0_405_2[1]));
    assign layer_0[405] = ~(far_0_405_2[0] ^ far_0_405_2[1]); 
    wire [1:0] far_0_406_0;    relay_conn far_0_406_0_a(.in(in[30]), .out(far_0_406_0[0]));    relay_conn far_0_406_0_b(.in(in[134]), .out(far_0_406_0[1]));
    wire [1:0] far_0_406_1;    relay_conn far_0_406_1_a(.in(far_0_406_0[0]), .out(far_0_406_1[0]));    relay_conn far_0_406_1_b(.in(far_0_406_0[1]), .out(far_0_406_1[1]));
    wire [1:0] far_0_406_2;    relay_conn far_0_406_2_a(.in(far_0_406_1[0]), .out(far_0_406_2[0]));    relay_conn far_0_406_2_b(.in(far_0_406_1[1]), .out(far_0_406_2[1]));
    assign layer_0[406] = ~(far_0_406_2[0] & far_0_406_2[1]); 
    wire [1:0] far_0_407_0;    relay_conn far_0_407_0_a(.in(in[169]), .out(far_0_407_0[0]));    relay_conn far_0_407_0_b(.in(in[99]), .out(far_0_407_0[1]));
    wire [1:0] far_0_407_1;    relay_conn far_0_407_1_a(.in(far_0_407_0[0]), .out(far_0_407_1[0]));    relay_conn far_0_407_1_b(.in(far_0_407_0[1]), .out(far_0_407_1[1]));
    assign layer_0[407] = far_0_407_1[0] & far_0_407_1[1]; 
    assign layer_0[408] = in[214] & ~in[191]; 
    wire [1:0] far_0_409_0;    relay_conn far_0_409_0_a(.in(in[131]), .out(far_0_409_0[0]));    relay_conn far_0_409_0_b(.in(in[167]), .out(far_0_409_0[1]));
    assign layer_0[409] = ~far_0_409_0[1]; 
    assign layer_0[410] = in[100]; 
    assign layer_0[411] = in[37] | in[52]; 
    wire [1:0] far_0_412_0;    relay_conn far_0_412_0_a(.in(in[125]), .out(far_0_412_0[0]));    relay_conn far_0_412_0_b(.in(in[199]), .out(far_0_412_0[1]));
    wire [1:0] far_0_412_1;    relay_conn far_0_412_1_a(.in(far_0_412_0[0]), .out(far_0_412_1[0]));    relay_conn far_0_412_1_b(.in(far_0_412_0[1]), .out(far_0_412_1[1]));
    assign layer_0[412] = far_0_412_1[0] & ~far_0_412_1[1]; 
    assign layer_0[413] = ~in[207] | (in[211] & in[207]); 
    wire [1:0] far_0_414_0;    relay_conn far_0_414_0_a(.in(in[6]), .out(far_0_414_0[0]));    relay_conn far_0_414_0_b(.in(in[133]), .out(far_0_414_0[1]));
    wire [1:0] far_0_414_1;    relay_conn far_0_414_1_a(.in(far_0_414_0[0]), .out(far_0_414_1[0]));    relay_conn far_0_414_1_b(.in(far_0_414_0[1]), .out(far_0_414_1[1]));
    wire [1:0] far_0_414_2;    relay_conn far_0_414_2_a(.in(far_0_414_1[0]), .out(far_0_414_2[0]));    relay_conn far_0_414_2_b(.in(far_0_414_1[1]), .out(far_0_414_2[1]));
    assign layer_0[414] = ~far_0_414_2[1]; 
    wire [1:0] far_0_415_0;    relay_conn far_0_415_0_a(.in(in[188]), .out(far_0_415_0[0]));    relay_conn far_0_415_0_b(.in(in[239]), .out(far_0_415_0[1]));
    assign layer_0[415] = ~(far_0_415_0[0] & far_0_415_0[1]); 
    wire [1:0] far_0_416_0;    relay_conn far_0_416_0_a(.in(in[207]), .out(far_0_416_0[0]));    relay_conn far_0_416_0_b(.in(in[130]), .out(far_0_416_0[1]));
    wire [1:0] far_0_416_1;    relay_conn far_0_416_1_a(.in(far_0_416_0[0]), .out(far_0_416_1[0]));    relay_conn far_0_416_1_b(.in(far_0_416_0[1]), .out(far_0_416_1[1]));
    assign layer_0[416] = far_0_416_1[0]; 
    assign layer_0[417] = ~(in[239] | in[240]); 
    wire [1:0] far_0_418_0;    relay_conn far_0_418_0_a(.in(in[142]), .out(far_0_418_0[0]));    relay_conn far_0_418_0_b(.in(in[239]), .out(far_0_418_0[1]));
    wire [1:0] far_0_418_1;    relay_conn far_0_418_1_a(.in(far_0_418_0[0]), .out(far_0_418_1[0]));    relay_conn far_0_418_1_b(.in(far_0_418_0[1]), .out(far_0_418_1[1]));
    wire [1:0] far_0_418_2;    relay_conn far_0_418_2_a(.in(far_0_418_1[0]), .out(far_0_418_2[0]));    relay_conn far_0_418_2_b(.in(far_0_418_1[1]), .out(far_0_418_2[1]));
    assign layer_0[418] = ~far_0_418_2[0]; 
    wire [1:0] far_0_419_0;    relay_conn far_0_419_0_a(.in(in[32]), .out(far_0_419_0[0]));    relay_conn far_0_419_0_b(.in(in[113]), .out(far_0_419_0[1]));
    wire [1:0] far_0_419_1;    relay_conn far_0_419_1_a(.in(far_0_419_0[0]), .out(far_0_419_1[0]));    relay_conn far_0_419_1_b(.in(far_0_419_0[1]), .out(far_0_419_1[1]));
    assign layer_0[419] = far_0_419_1[1] & ~far_0_419_1[0]; 
    wire [1:0] far_0_420_0;    relay_conn far_0_420_0_a(.in(in[132]), .out(far_0_420_0[0]));    relay_conn far_0_420_0_b(.in(in[176]), .out(far_0_420_0[1]));
    assign layer_0[420] = ~(far_0_420_0[0] ^ far_0_420_0[1]); 
    wire [1:0] far_0_421_0;    relay_conn far_0_421_0_a(.in(in[244]), .out(far_0_421_0[0]));    relay_conn far_0_421_0_b(.in(in[151]), .out(far_0_421_0[1]));
    wire [1:0] far_0_421_1;    relay_conn far_0_421_1_a(.in(far_0_421_0[0]), .out(far_0_421_1[0]));    relay_conn far_0_421_1_b(.in(far_0_421_0[1]), .out(far_0_421_1[1]));
    assign layer_0[421] = far_0_421_1[0] | far_0_421_1[1]; 
    assign layer_0[422] = ~(in[149] ^ in[121]); 
    assign layer_0[423] = ~in[236]; 
    assign layer_0[424] = in[151] | in[172]; 
    wire [1:0] far_0_425_0;    relay_conn far_0_425_0_a(.in(in[10]), .out(far_0_425_0[0]));    relay_conn far_0_425_0_b(.in(in[79]), .out(far_0_425_0[1]));
    wire [1:0] far_0_425_1;    relay_conn far_0_425_1_a(.in(far_0_425_0[0]), .out(far_0_425_1[0]));    relay_conn far_0_425_1_b(.in(far_0_425_0[1]), .out(far_0_425_1[1]));
    assign layer_0[425] = far_0_425_1[0] & ~far_0_425_1[1]; 
    wire [1:0] far_0_426_0;    relay_conn far_0_426_0_a(.in(in[245]), .out(far_0_426_0[0]));    relay_conn far_0_426_0_b(.in(in[138]), .out(far_0_426_0[1]));
    wire [1:0] far_0_426_1;    relay_conn far_0_426_1_a(.in(far_0_426_0[0]), .out(far_0_426_1[0]));    relay_conn far_0_426_1_b(.in(far_0_426_0[1]), .out(far_0_426_1[1]));
    wire [1:0] far_0_426_2;    relay_conn far_0_426_2_a(.in(far_0_426_1[0]), .out(far_0_426_2[0]));    relay_conn far_0_426_2_b(.in(far_0_426_1[1]), .out(far_0_426_2[1]));
    assign layer_0[426] = far_0_426_2[0] & far_0_426_2[1]; 
    assign layer_0[427] = in[13]; 
    assign layer_0[428] = in[211] & in[241]; 
    wire [1:0] far_0_429_0;    relay_conn far_0_429_0_a(.in(in[109]), .out(far_0_429_0[0]));    relay_conn far_0_429_0_b(.in(in[34]), .out(far_0_429_0[1]));
    wire [1:0] far_0_429_1;    relay_conn far_0_429_1_a(.in(far_0_429_0[0]), .out(far_0_429_1[0]));    relay_conn far_0_429_1_b(.in(far_0_429_0[1]), .out(far_0_429_1[1]));
    assign layer_0[429] = far_0_429_1[0] & ~far_0_429_1[1]; 
    wire [1:0] far_0_430_0;    relay_conn far_0_430_0_a(.in(in[73]), .out(far_0_430_0[0]));    relay_conn far_0_430_0_b(.in(in[107]), .out(far_0_430_0[1]));
    assign layer_0[430] = ~(far_0_430_0[0] | far_0_430_0[1]); 
    wire [1:0] far_0_431_0;    relay_conn far_0_431_0_a(.in(in[79]), .out(far_0_431_0[0]));    relay_conn far_0_431_0_b(.in(in[165]), .out(far_0_431_0[1]));
    wire [1:0] far_0_431_1;    relay_conn far_0_431_1_a(.in(far_0_431_0[0]), .out(far_0_431_1[0]));    relay_conn far_0_431_1_b(.in(far_0_431_0[1]), .out(far_0_431_1[1]));
    assign layer_0[431] = ~far_0_431_1[1] | (far_0_431_1[0] & far_0_431_1[1]); 
    wire [1:0] far_0_432_0;    relay_conn far_0_432_0_a(.in(in[101]), .out(far_0_432_0[0]));    relay_conn far_0_432_0_b(.in(in[188]), .out(far_0_432_0[1]));
    wire [1:0] far_0_432_1;    relay_conn far_0_432_1_a(.in(far_0_432_0[0]), .out(far_0_432_1[0]));    relay_conn far_0_432_1_b(.in(far_0_432_0[1]), .out(far_0_432_1[1]));
    assign layer_0[432] = far_0_432_1[0] & far_0_432_1[1]; 
    wire [1:0] far_0_433_0;    relay_conn far_0_433_0_a(.in(in[187]), .out(far_0_433_0[0]));    relay_conn far_0_433_0_b(.in(in[233]), .out(far_0_433_0[1]));
    assign layer_0[433] = ~(far_0_433_0[0] & far_0_433_0[1]); 
    assign layer_0[434] = ~in[43]; 
    assign layer_0[435] = ~(in[111] | in[125]); 
    wire [1:0] far_0_436_0;    relay_conn far_0_436_0_a(.in(in[3]), .out(far_0_436_0[0]));    relay_conn far_0_436_0_b(.in(in[105]), .out(far_0_436_0[1]));
    wire [1:0] far_0_436_1;    relay_conn far_0_436_1_a(.in(far_0_436_0[0]), .out(far_0_436_1[0]));    relay_conn far_0_436_1_b(.in(far_0_436_0[1]), .out(far_0_436_1[1]));
    wire [1:0] far_0_436_2;    relay_conn far_0_436_2_a(.in(far_0_436_1[0]), .out(far_0_436_2[0]));    relay_conn far_0_436_2_b(.in(far_0_436_1[1]), .out(far_0_436_2[1]));
    assign layer_0[436] = far_0_436_2[0] ^ far_0_436_2[1]; 
    wire [1:0] far_0_437_0;    relay_conn far_0_437_0_a(.in(in[57]), .out(far_0_437_0[0]));    relay_conn far_0_437_0_b(.in(in[178]), .out(far_0_437_0[1]));
    wire [1:0] far_0_437_1;    relay_conn far_0_437_1_a(.in(far_0_437_0[0]), .out(far_0_437_1[0]));    relay_conn far_0_437_1_b(.in(far_0_437_0[1]), .out(far_0_437_1[1]));
    wire [1:0] far_0_437_2;    relay_conn far_0_437_2_a(.in(far_0_437_1[0]), .out(far_0_437_2[0]));    relay_conn far_0_437_2_b(.in(far_0_437_1[1]), .out(far_0_437_2[1]));
    assign layer_0[437] = far_0_437_2[1]; 
    wire [1:0] far_0_438_0;    relay_conn far_0_438_0_a(.in(in[82]), .out(far_0_438_0[0]));    relay_conn far_0_438_0_b(.in(in[158]), .out(far_0_438_0[1]));
    wire [1:0] far_0_438_1;    relay_conn far_0_438_1_a(.in(far_0_438_0[0]), .out(far_0_438_1[0]));    relay_conn far_0_438_1_b(.in(far_0_438_0[1]), .out(far_0_438_1[1]));
    assign layer_0[438] = far_0_438_1[0] ^ far_0_438_1[1]; 
    wire [1:0] far_0_439_0;    relay_conn far_0_439_0_a(.in(in[164]), .out(far_0_439_0[0]));    relay_conn far_0_439_0_b(.in(in[202]), .out(far_0_439_0[1]));
    assign layer_0[439] = ~far_0_439_0[1] | (far_0_439_0[0] & far_0_439_0[1]); 
    assign layer_0[440] = ~in[233] | (in[233] & in[211]); 
    assign layer_0[441] = ~in[137]; 
    assign layer_0[442] = ~in[56] | (in[72] & in[56]); 
    wire [1:0] far_0_443_0;    relay_conn far_0_443_0_a(.in(in[34]), .out(far_0_443_0[0]));    relay_conn far_0_443_0_b(.in(in[69]), .out(far_0_443_0[1]));
    assign layer_0[443] = ~far_0_443_0[0] | (far_0_443_0[0] & far_0_443_0[1]); 
    wire [1:0] far_0_444_0;    relay_conn far_0_444_0_a(.in(in[97]), .out(far_0_444_0[0]));    relay_conn far_0_444_0_b(.in(in[158]), .out(far_0_444_0[1]));
    assign layer_0[444] = far_0_444_0[1]; 
    wire [1:0] far_0_445_0;    relay_conn far_0_445_0_a(.in(in[103]), .out(far_0_445_0[0]));    relay_conn far_0_445_0_b(.in(in[215]), .out(far_0_445_0[1]));
    wire [1:0] far_0_445_1;    relay_conn far_0_445_1_a(.in(far_0_445_0[0]), .out(far_0_445_1[0]));    relay_conn far_0_445_1_b(.in(far_0_445_0[1]), .out(far_0_445_1[1]));
    wire [1:0] far_0_445_2;    relay_conn far_0_445_2_a(.in(far_0_445_1[0]), .out(far_0_445_2[0]));    relay_conn far_0_445_2_b(.in(far_0_445_1[1]), .out(far_0_445_2[1]));
    assign layer_0[445] = ~far_0_445_2[0] | (far_0_445_2[0] & far_0_445_2[1]); 
    assign layer_0[446] = in[73]; 
    wire [1:0] far_0_447_0;    relay_conn far_0_447_0_a(.in(in[23]), .out(far_0_447_0[0]));    relay_conn far_0_447_0_b(.in(in[75]), .out(far_0_447_0[1]));
    assign layer_0[447] = ~(far_0_447_0[0] | far_0_447_0[1]); 
    wire [1:0] far_0_448_0;    relay_conn far_0_448_0_a(.in(in[222]), .out(far_0_448_0[0]));    relay_conn far_0_448_0_b(.in(in[111]), .out(far_0_448_0[1]));
    wire [1:0] far_0_448_1;    relay_conn far_0_448_1_a(.in(far_0_448_0[0]), .out(far_0_448_1[0]));    relay_conn far_0_448_1_b(.in(far_0_448_0[1]), .out(far_0_448_1[1]));
    wire [1:0] far_0_448_2;    relay_conn far_0_448_2_a(.in(far_0_448_1[0]), .out(far_0_448_2[0]));    relay_conn far_0_448_2_b(.in(far_0_448_1[1]), .out(far_0_448_2[1]));
    assign layer_0[448] = ~(far_0_448_2[0] | far_0_448_2[1]); 
    wire [1:0] far_0_449_0;    relay_conn far_0_449_0_a(.in(in[136]), .out(far_0_449_0[0]));    relay_conn far_0_449_0_b(.in(in[72]), .out(far_0_449_0[1]));
    wire [1:0] far_0_449_1;    relay_conn far_0_449_1_a(.in(far_0_449_0[0]), .out(far_0_449_1[0]));    relay_conn far_0_449_1_b(.in(far_0_449_0[1]), .out(far_0_449_1[1]));
    assign layer_0[449] = ~far_0_449_1[1] | (far_0_449_1[0] & far_0_449_1[1]); 
    wire [1:0] far_0_450_0;    relay_conn far_0_450_0_a(.in(in[38]), .out(far_0_450_0[0]));    relay_conn far_0_450_0_b(.in(in[151]), .out(far_0_450_0[1]));
    wire [1:0] far_0_450_1;    relay_conn far_0_450_1_a(.in(far_0_450_0[0]), .out(far_0_450_1[0]));    relay_conn far_0_450_1_b(.in(far_0_450_0[1]), .out(far_0_450_1[1]));
    wire [1:0] far_0_450_2;    relay_conn far_0_450_2_a(.in(far_0_450_1[0]), .out(far_0_450_2[0]));    relay_conn far_0_450_2_b(.in(far_0_450_1[1]), .out(far_0_450_2[1]));
    assign layer_0[450] = far_0_450_2[1]; 
    wire [1:0] far_0_451_0;    relay_conn far_0_451_0_a(.in(in[87]), .out(far_0_451_0[0]));    relay_conn far_0_451_0_b(.in(in[133]), .out(far_0_451_0[1]));
    assign layer_0[451] = ~(far_0_451_0[0] ^ far_0_451_0[1]); 
    assign layer_0[452] = in[186] | in[167]; 
    wire [1:0] far_0_453_0;    relay_conn far_0_453_0_a(.in(in[198]), .out(far_0_453_0[0]));    relay_conn far_0_453_0_b(.in(in[113]), .out(far_0_453_0[1]));
    wire [1:0] far_0_453_1;    relay_conn far_0_453_1_a(.in(far_0_453_0[0]), .out(far_0_453_1[0]));    relay_conn far_0_453_1_b(.in(far_0_453_0[1]), .out(far_0_453_1[1]));
    assign layer_0[453] = ~(far_0_453_1[0] ^ far_0_453_1[1]); 
    wire [1:0] far_0_454_0;    relay_conn far_0_454_0_a(.in(in[97]), .out(far_0_454_0[0]));    relay_conn far_0_454_0_b(.in(in[23]), .out(far_0_454_0[1]));
    wire [1:0] far_0_454_1;    relay_conn far_0_454_1_a(.in(far_0_454_0[0]), .out(far_0_454_1[0]));    relay_conn far_0_454_1_b(.in(far_0_454_0[1]), .out(far_0_454_1[1]));
    assign layer_0[454] = far_0_454_1[0] & ~far_0_454_1[1]; 
    wire [1:0] far_0_455_0;    relay_conn far_0_455_0_a(.in(in[96]), .out(far_0_455_0[0]));    relay_conn far_0_455_0_b(.in(in[35]), .out(far_0_455_0[1]));
    assign layer_0[455] = far_0_455_0[0] & far_0_455_0[1]; 
    assign layer_0[456] = in[119] & ~in[109]; 
    assign layer_0[457] = ~in[113] | (in[113] & in[88]); 
    wire [1:0] far_0_458_0;    relay_conn far_0_458_0_a(.in(in[199]), .out(far_0_458_0[0]));    relay_conn far_0_458_0_b(.in(in[87]), .out(far_0_458_0[1]));
    wire [1:0] far_0_458_1;    relay_conn far_0_458_1_a(.in(far_0_458_0[0]), .out(far_0_458_1[0]));    relay_conn far_0_458_1_b(.in(far_0_458_0[1]), .out(far_0_458_1[1]));
    wire [1:0] far_0_458_2;    relay_conn far_0_458_2_a(.in(far_0_458_1[0]), .out(far_0_458_2[0]));    relay_conn far_0_458_2_b(.in(far_0_458_1[1]), .out(far_0_458_2[1]));
    assign layer_0[458] = far_0_458_2[0] & far_0_458_2[1]; 
    wire [1:0] far_0_459_0;    relay_conn far_0_459_0_a(.in(in[208]), .out(far_0_459_0[0]));    relay_conn far_0_459_0_b(.in(in[134]), .out(far_0_459_0[1]));
    wire [1:0] far_0_459_1;    relay_conn far_0_459_1_a(.in(far_0_459_0[0]), .out(far_0_459_1[0]));    relay_conn far_0_459_1_b(.in(far_0_459_0[1]), .out(far_0_459_1[1]));
    assign layer_0[459] = ~far_0_459_1[0]; 
    wire [1:0] far_0_460_0;    relay_conn far_0_460_0_a(.in(in[91]), .out(far_0_460_0[0]));    relay_conn far_0_460_0_b(.in(in[25]), .out(far_0_460_0[1]));
    wire [1:0] far_0_460_1;    relay_conn far_0_460_1_a(.in(far_0_460_0[0]), .out(far_0_460_1[0]));    relay_conn far_0_460_1_b(.in(far_0_460_0[1]), .out(far_0_460_1[1]));
    assign layer_0[460] = far_0_460_1[0] ^ far_0_460_1[1]; 
    assign layer_0[461] = ~in[18]; 
    assign layer_0[462] = in[185] | in[172]; 
    wire [1:0] far_0_463_0;    relay_conn far_0_463_0_a(.in(in[215]), .out(far_0_463_0[0]));    relay_conn far_0_463_0_b(.in(in[133]), .out(far_0_463_0[1]));
    wire [1:0] far_0_463_1;    relay_conn far_0_463_1_a(.in(far_0_463_0[0]), .out(far_0_463_1[0]));    relay_conn far_0_463_1_b(.in(far_0_463_0[1]), .out(far_0_463_1[1]));
    assign layer_0[463] = far_0_463_1[0] | far_0_463_1[1]; 
    assign layer_0[464] = ~in[34]; 
    wire [1:0] far_0_465_0;    relay_conn far_0_465_0_a(.in(in[158]), .out(far_0_465_0[0]));    relay_conn far_0_465_0_b(.in(in[247]), .out(far_0_465_0[1]));
    wire [1:0] far_0_465_1;    relay_conn far_0_465_1_a(.in(far_0_465_0[0]), .out(far_0_465_1[0]));    relay_conn far_0_465_1_b(.in(far_0_465_0[1]), .out(far_0_465_1[1]));
    assign layer_0[465] = ~(far_0_465_1[0] ^ far_0_465_1[1]); 
    wire [1:0] far_0_466_0;    relay_conn far_0_466_0_a(.in(in[88]), .out(far_0_466_0[0]));    relay_conn far_0_466_0_b(.in(in[32]), .out(far_0_466_0[1]));
    assign layer_0[466] = ~(far_0_466_0[0] & far_0_466_0[1]); 
    wire [1:0] far_0_467_0;    relay_conn far_0_467_0_a(.in(in[172]), .out(far_0_467_0[0]));    relay_conn far_0_467_0_b(.in(in[215]), .out(far_0_467_0[1]));
    assign layer_0[467] = far_0_467_0[0] | far_0_467_0[1]; 
    wire [1:0] far_0_468_0;    relay_conn far_0_468_0_a(.in(in[145]), .out(far_0_468_0[0]));    relay_conn far_0_468_0_b(.in(in[241]), .out(far_0_468_0[1]));
    wire [1:0] far_0_468_1;    relay_conn far_0_468_1_a(.in(far_0_468_0[0]), .out(far_0_468_1[0]));    relay_conn far_0_468_1_b(.in(far_0_468_0[1]), .out(far_0_468_1[1]));
    wire [1:0] far_0_468_2;    relay_conn far_0_468_2_a(.in(far_0_468_1[0]), .out(far_0_468_2[0]));    relay_conn far_0_468_2_b(.in(far_0_468_1[1]), .out(far_0_468_2[1]));
    assign layer_0[468] = far_0_468_2[0] & far_0_468_2[1]; 
    wire [1:0] far_0_469_0;    relay_conn far_0_469_0_a(.in(in[48]), .out(far_0_469_0[0]));    relay_conn far_0_469_0_b(.in(in[143]), .out(far_0_469_0[1]));
    wire [1:0] far_0_469_1;    relay_conn far_0_469_1_a(.in(far_0_469_0[0]), .out(far_0_469_1[0]));    relay_conn far_0_469_1_b(.in(far_0_469_0[1]), .out(far_0_469_1[1]));
    assign layer_0[469] = far_0_469_1[0] | far_0_469_1[1]; 
    assign layer_0[470] = ~in[30] | (in[30] & in[57]); 
    wire [1:0] far_0_471_0;    relay_conn far_0_471_0_a(.in(in[199]), .out(far_0_471_0[0]));    relay_conn far_0_471_0_b(.in(in[132]), .out(far_0_471_0[1]));
    wire [1:0] far_0_471_1;    relay_conn far_0_471_1_a(.in(far_0_471_0[0]), .out(far_0_471_1[0]));    relay_conn far_0_471_1_b(.in(far_0_471_0[1]), .out(far_0_471_1[1]));
    assign layer_0[471] = ~far_0_471_1[1] | (far_0_471_1[0] & far_0_471_1[1]); 
    wire [1:0] far_0_472_0;    relay_conn far_0_472_0_a(.in(in[189]), .out(far_0_472_0[0]));    relay_conn far_0_472_0_b(.in(in[132]), .out(far_0_472_0[1]));
    assign layer_0[472] = far_0_472_0[0] & far_0_472_0[1]; 
    assign layer_0[473] = in[223] & in[212]; 
    assign layer_0[474] = ~in[197] | (in[225] & in[197]); 
    wire [1:0] far_0_475_0;    relay_conn far_0_475_0_a(.in(in[122]), .out(far_0_475_0[0]));    relay_conn far_0_475_0_b(.in(in[213]), .out(far_0_475_0[1]));
    wire [1:0] far_0_475_1;    relay_conn far_0_475_1_a(.in(far_0_475_0[0]), .out(far_0_475_1[0]));    relay_conn far_0_475_1_b(.in(far_0_475_0[1]), .out(far_0_475_1[1]));
    assign layer_0[475] = far_0_475_1[0] & far_0_475_1[1]; 
    wire [1:0] far_0_476_0;    relay_conn far_0_476_0_a(.in(in[30]), .out(far_0_476_0[0]));    relay_conn far_0_476_0_b(.in(in[132]), .out(far_0_476_0[1]));
    wire [1:0] far_0_476_1;    relay_conn far_0_476_1_a(.in(far_0_476_0[0]), .out(far_0_476_1[0]));    relay_conn far_0_476_1_b(.in(far_0_476_0[1]), .out(far_0_476_1[1]));
    wire [1:0] far_0_476_2;    relay_conn far_0_476_2_a(.in(far_0_476_1[0]), .out(far_0_476_2[0]));    relay_conn far_0_476_2_b(.in(far_0_476_1[1]), .out(far_0_476_2[1]));
    assign layer_0[476] = ~far_0_476_2[1] | (far_0_476_2[0] & far_0_476_2[1]); 
    assign layer_0[477] = ~in[113] | (in[113] & in[138]); 
    wire [1:0] far_0_478_0;    relay_conn far_0_478_0_a(.in(in[226]), .out(far_0_478_0[0]));    relay_conn far_0_478_0_b(.in(in[109]), .out(far_0_478_0[1]));
    wire [1:0] far_0_478_1;    relay_conn far_0_478_1_a(.in(far_0_478_0[0]), .out(far_0_478_1[0]));    relay_conn far_0_478_1_b(.in(far_0_478_0[1]), .out(far_0_478_1[1]));
    wire [1:0] far_0_478_2;    relay_conn far_0_478_2_a(.in(far_0_478_1[0]), .out(far_0_478_2[0]));    relay_conn far_0_478_2_b(.in(far_0_478_1[1]), .out(far_0_478_2[1]));
    assign layer_0[478] = ~far_0_478_2[0]; 
    wire [1:0] far_0_479_0;    relay_conn far_0_479_0_a(.in(in[188]), .out(far_0_479_0[0]));    relay_conn far_0_479_0_b(.in(in[230]), .out(far_0_479_0[1]));
    assign layer_0[479] = far_0_479_0[1]; 
    wire [1:0] far_0_480_0;    relay_conn far_0_480_0_a(.in(in[150]), .out(far_0_480_0[0]));    relay_conn far_0_480_0_b(.in(in[71]), .out(far_0_480_0[1]));
    wire [1:0] far_0_480_1;    relay_conn far_0_480_1_a(.in(far_0_480_0[0]), .out(far_0_480_1[0]));    relay_conn far_0_480_1_b(.in(far_0_480_0[1]), .out(far_0_480_1[1]));
    assign layer_0[480] = far_0_480_1[0] & ~far_0_480_1[1]; 
    assign layer_0[481] = ~in[233]; 
    wire [1:0] far_0_482_0;    relay_conn far_0_482_0_a(.in(in[199]), .out(far_0_482_0[0]));    relay_conn far_0_482_0_b(.in(in[148]), .out(far_0_482_0[1]));
    assign layer_0[482] = far_0_482_0[0] ^ far_0_482_0[1]; 
    wire [1:0] far_0_483_0;    relay_conn far_0_483_0_a(.in(in[229]), .out(far_0_483_0[0]));    relay_conn far_0_483_0_b(.in(in[117]), .out(far_0_483_0[1]));
    wire [1:0] far_0_483_1;    relay_conn far_0_483_1_a(.in(far_0_483_0[0]), .out(far_0_483_1[0]));    relay_conn far_0_483_1_b(.in(far_0_483_0[1]), .out(far_0_483_1[1]));
    wire [1:0] far_0_483_2;    relay_conn far_0_483_2_a(.in(far_0_483_1[0]), .out(far_0_483_2[0]));    relay_conn far_0_483_2_b(.in(far_0_483_1[1]), .out(far_0_483_2[1]));
    assign layer_0[483] = ~(far_0_483_2[0] ^ far_0_483_2[1]); 
    assign layer_0[484] = in[71] ^ in[41]; 
    wire [1:0] far_0_485_0;    relay_conn far_0_485_0_a(.in(in[113]), .out(far_0_485_0[0]));    relay_conn far_0_485_0_b(.in(in[173]), .out(far_0_485_0[1]));
    assign layer_0[485] = far_0_485_0[1] & ~far_0_485_0[0]; 
    wire [1:0] far_0_486_0;    relay_conn far_0_486_0_a(.in(in[135]), .out(far_0_486_0[0]));    relay_conn far_0_486_0_b(.in(in[203]), .out(far_0_486_0[1]));
    wire [1:0] far_0_486_1;    relay_conn far_0_486_1_a(.in(far_0_486_0[0]), .out(far_0_486_1[0]));    relay_conn far_0_486_1_b(.in(far_0_486_0[1]), .out(far_0_486_1[1]));
    assign layer_0[486] = far_0_486_1[0] | far_0_486_1[1]; 
    assign layer_0[487] = in[66]; 
    assign layer_0[488] = ~in[191]; 
    assign layer_0[489] = in[199]; 
    assign layer_0[490] = ~in[18]; 
    wire [1:0] far_0_491_0;    relay_conn far_0_491_0_a(.in(in[134]), .out(far_0_491_0[0]));    relay_conn far_0_491_0_b(.in(in[189]), .out(far_0_491_0[1]));
    assign layer_0[491] = far_0_491_0[0] & far_0_491_0[1]; 
    assign layer_0[492] = in[185] | in[188]; 
    wire [1:0] far_0_493_0;    relay_conn far_0_493_0_a(.in(in[74]), .out(far_0_493_0[0]));    relay_conn far_0_493_0_b(.in(in[41]), .out(far_0_493_0[1]));
    assign layer_0[493] = ~(far_0_493_0[0] | far_0_493_0[1]); 
    wire [1:0] far_0_494_0;    relay_conn far_0_494_0_a(.in(in[82]), .out(far_0_494_0[0]));    relay_conn far_0_494_0_b(.in(in[15]), .out(far_0_494_0[1]));
    wire [1:0] far_0_494_1;    relay_conn far_0_494_1_a(.in(far_0_494_0[0]), .out(far_0_494_1[0]));    relay_conn far_0_494_1_b(.in(far_0_494_0[1]), .out(far_0_494_1[1]));
    assign layer_0[494] = far_0_494_1[0] | far_0_494_1[1]; 
    assign layer_0[495] = in[117] | in[87]; 
    wire [1:0] far_0_496_0;    relay_conn far_0_496_0_a(.in(in[27]), .out(far_0_496_0[0]));    relay_conn far_0_496_0_b(.in(in[87]), .out(far_0_496_0[1]));
    assign layer_0[496] = far_0_496_0[1] & ~far_0_496_0[0]; 
    assign layer_0[497] = in[203] & in[188]; 
    wire [1:0] far_0_498_0;    relay_conn far_0_498_0_a(.in(in[61]), .out(far_0_498_0[0]));    relay_conn far_0_498_0_b(.in(in[95]), .out(far_0_498_0[1]));
    assign layer_0[498] = far_0_498_0[0] ^ far_0_498_0[1]; 
    assign layer_0[499] = in[127]; 
    wire [1:0] far_0_500_0;    relay_conn far_0_500_0_a(.in(in[57]), .out(far_0_500_0[0]));    relay_conn far_0_500_0_b(.in(in[117]), .out(far_0_500_0[1]));
    assign layer_0[500] = ~far_0_500_0[0] | (far_0_500_0[0] & far_0_500_0[1]); 
    wire [1:0] far_0_501_0;    relay_conn far_0_501_0_a(.in(in[79]), .out(far_0_501_0[0]));    relay_conn far_0_501_0_b(.in(in[151]), .out(far_0_501_0[1]));
    wire [1:0] far_0_501_1;    relay_conn far_0_501_1_a(.in(far_0_501_0[0]), .out(far_0_501_1[0]));    relay_conn far_0_501_1_b(.in(far_0_501_0[1]), .out(far_0_501_1[1]));
    assign layer_0[501] = far_0_501_1[1] & ~far_0_501_1[0]; 
    wire [1:0] far_0_502_0;    relay_conn far_0_502_0_a(.in(in[6]), .out(far_0_502_0[0]));    relay_conn far_0_502_0_b(.in(in[79]), .out(far_0_502_0[1]));
    wire [1:0] far_0_502_1;    relay_conn far_0_502_1_a(.in(far_0_502_0[0]), .out(far_0_502_1[0]));    relay_conn far_0_502_1_b(.in(far_0_502_0[1]), .out(far_0_502_1[1]));
    assign layer_0[502] = ~far_0_502_1[0] | (far_0_502_1[0] & far_0_502_1[1]); 
    assign layer_0[503] = ~in[0] | (in[0] & in[29]); 
    wire [1:0] far_0_504_0;    relay_conn far_0_504_0_a(.in(in[199]), .out(far_0_504_0[0]));    relay_conn far_0_504_0_b(.in(in[135]), .out(far_0_504_0[1]));
    wire [1:0] far_0_504_1;    relay_conn far_0_504_1_a(.in(far_0_504_0[0]), .out(far_0_504_1[0]));    relay_conn far_0_504_1_b(.in(far_0_504_0[1]), .out(far_0_504_1[1]));
    assign layer_0[504] = far_0_504_1[1]; 
    assign layer_0[505] = in[223]; 
    wire [1:0] far_0_506_0;    relay_conn far_0_506_0_a(.in(in[110]), .out(far_0_506_0[0]));    relay_conn far_0_506_0_b(.in(in[202]), .out(far_0_506_0[1]));
    wire [1:0] far_0_506_1;    relay_conn far_0_506_1_a(.in(far_0_506_0[0]), .out(far_0_506_1[0]));    relay_conn far_0_506_1_b(.in(far_0_506_0[1]), .out(far_0_506_1[1]));
    assign layer_0[506] = ~(far_0_506_1[0] | far_0_506_1[1]); 
    assign layer_0[507] = ~(in[65] | in[73]); 
    assign layer_0[508] = ~in[171] | (in[171] & in[188]); 
    assign layer_0[509] = in[185] & ~in[172]; 
    wire [1:0] far_0_510_0;    relay_conn far_0_510_0_a(.in(in[87]), .out(far_0_510_0[0]));    relay_conn far_0_510_0_b(.in(in[194]), .out(far_0_510_0[1]));
    wire [1:0] far_0_510_1;    relay_conn far_0_510_1_a(.in(far_0_510_0[0]), .out(far_0_510_1[0]));    relay_conn far_0_510_1_b(.in(far_0_510_0[1]), .out(far_0_510_1[1]));
    wire [1:0] far_0_510_2;    relay_conn far_0_510_2_a(.in(far_0_510_1[0]), .out(far_0_510_2[0]));    relay_conn far_0_510_2_b(.in(far_0_510_1[1]), .out(far_0_510_2[1]));
    assign layer_0[510] = far_0_510_2[1]; 
    wire [1:0] far_0_511_0;    relay_conn far_0_511_0_a(.in(in[199]), .out(far_0_511_0[0]));    relay_conn far_0_511_0_b(.in(in[112]), .out(far_0_511_0[1]));
    wire [1:0] far_0_511_1;    relay_conn far_0_511_1_a(.in(far_0_511_0[0]), .out(far_0_511_1[0]));    relay_conn far_0_511_1_b(.in(far_0_511_0[1]), .out(far_0_511_1[1]));
    assign layer_0[511] = ~far_0_511_1[1] | (far_0_511_1[0] & far_0_511_1[1]); 
    wire [1:0] far_0_512_0;    relay_conn far_0_512_0_a(.in(in[41]), .out(far_0_512_0[0]));    relay_conn far_0_512_0_b(.in(in[113]), .out(far_0_512_0[1]));
    wire [1:0] far_0_512_1;    relay_conn far_0_512_1_a(.in(far_0_512_0[0]), .out(far_0_512_1[0]));    relay_conn far_0_512_1_b(.in(far_0_512_0[1]), .out(far_0_512_1[1]));
    assign layer_0[512] = ~far_0_512_1[0]; 
    wire [1:0] far_0_513_0;    relay_conn far_0_513_0_a(.in(in[148]), .out(far_0_513_0[0]));    relay_conn far_0_513_0_b(.in(in[116]), .out(far_0_513_0[1]));
    assign layer_0[513] = ~far_0_513_0[0] | (far_0_513_0[0] & far_0_513_0[1]); 
    assign layer_0[514] = in[202]; 
    wire [1:0] far_0_515_0;    relay_conn far_0_515_0_a(.in(in[37]), .out(far_0_515_0[0]));    relay_conn far_0_515_0_b(.in(in[134]), .out(far_0_515_0[1]));
    wire [1:0] far_0_515_1;    relay_conn far_0_515_1_a(.in(far_0_515_0[0]), .out(far_0_515_1[0]));    relay_conn far_0_515_1_b(.in(far_0_515_0[1]), .out(far_0_515_1[1]));
    wire [1:0] far_0_515_2;    relay_conn far_0_515_2_a(.in(far_0_515_1[0]), .out(far_0_515_2[0]));    relay_conn far_0_515_2_b(.in(far_0_515_1[1]), .out(far_0_515_2[1]));
    assign layer_0[515] = ~(far_0_515_2[0] & far_0_515_2[1]); 
    wire [1:0] far_0_516_0;    relay_conn far_0_516_0_a(.in(in[77]), .out(far_0_516_0[0]));    relay_conn far_0_516_0_b(.in(in[138]), .out(far_0_516_0[1]));
    assign layer_0[516] = far_0_516_0[0]; 
    assign layer_0[517] = in[173]; 
    assign layer_0[518] = in[61] ^ in[73]; 
    wire [1:0] far_0_519_0;    relay_conn far_0_519_0_a(.in(in[34]), .out(far_0_519_0[0]));    relay_conn far_0_519_0_b(.in(in[0]), .out(far_0_519_0[1]));
    assign layer_0[519] = ~(far_0_519_0[0] | far_0_519_0[1]); 
    assign layer_0[520] = in[181] & ~in[178]; 
    assign layer_0[521] = in[3] & in[13]; 
    assign layer_0[522] = ~in[181]; 
    assign layer_0[523] = ~(in[25] & in[3]); 
    wire [1:0] far_0_524_0;    relay_conn far_0_524_0_a(.in(in[165]), .out(far_0_524_0[0]));    relay_conn far_0_524_0_b(.in(in[77]), .out(far_0_524_0[1]));
    wire [1:0] far_0_524_1;    relay_conn far_0_524_1_a(.in(far_0_524_0[0]), .out(far_0_524_1[0]));    relay_conn far_0_524_1_b(.in(far_0_524_0[1]), .out(far_0_524_1[1]));
    assign layer_0[524] = far_0_524_1[0] & ~far_0_524_1[1]; 
    wire [1:0] far_0_525_0;    relay_conn far_0_525_0_a(.in(in[7]), .out(far_0_525_0[0]));    relay_conn far_0_525_0_b(.in(in[72]), .out(far_0_525_0[1]));
    wire [1:0] far_0_525_1;    relay_conn far_0_525_1_a(.in(far_0_525_0[0]), .out(far_0_525_1[0]));    relay_conn far_0_525_1_b(.in(far_0_525_0[1]), .out(far_0_525_1[1]));
    assign layer_0[525] = ~(far_0_525_1[0] | far_0_525_1[1]); 
    wire [1:0] far_0_526_0;    relay_conn far_0_526_0_a(.in(in[125]), .out(far_0_526_0[0]));    relay_conn far_0_526_0_b(.in(in[66]), .out(far_0_526_0[1]));
    assign layer_0[526] = far_0_526_0[0] ^ far_0_526_0[1]; 
    assign layer_0[527] = ~in[79]; 
    wire [1:0] far_0_528_0;    relay_conn far_0_528_0_a(.in(in[250]), .out(far_0_528_0[0]));    relay_conn far_0_528_0_b(.in(in[152]), .out(far_0_528_0[1]));
    wire [1:0] far_0_528_1;    relay_conn far_0_528_1_a(.in(far_0_528_0[0]), .out(far_0_528_1[0]));    relay_conn far_0_528_1_b(.in(far_0_528_0[1]), .out(far_0_528_1[1]));
    wire [1:0] far_0_528_2;    relay_conn far_0_528_2_a(.in(far_0_528_1[0]), .out(far_0_528_2[0]));    relay_conn far_0_528_2_b(.in(far_0_528_1[1]), .out(far_0_528_2[1]));
    assign layer_0[528] = far_0_528_2[0] | far_0_528_2[1]; 
    wire [1:0] far_0_529_0;    relay_conn far_0_529_0_a(.in(in[211]), .out(far_0_529_0[0]));    relay_conn far_0_529_0_b(.in(in[172]), .out(far_0_529_0[1]));
    assign layer_0[529] = far_0_529_0[0] ^ far_0_529_0[1]; 
    wire [1:0] far_0_530_0;    relay_conn far_0_530_0_a(.in(in[135]), .out(far_0_530_0[0]));    relay_conn far_0_530_0_b(.in(in[191]), .out(far_0_530_0[1]));
    assign layer_0[530] = ~(far_0_530_0[0] ^ far_0_530_0[1]); 
    wire [1:0] far_0_531_0;    relay_conn far_0_531_0_a(.in(in[25]), .out(far_0_531_0[0]));    relay_conn far_0_531_0_b(.in(in[117]), .out(far_0_531_0[1]));
    wire [1:0] far_0_531_1;    relay_conn far_0_531_1_a(.in(far_0_531_0[0]), .out(far_0_531_1[0]));    relay_conn far_0_531_1_b(.in(far_0_531_0[1]), .out(far_0_531_1[1]));
    assign layer_0[531] = far_0_531_1[0] | far_0_531_1[1]; 
    wire [1:0] far_0_532_0;    relay_conn far_0_532_0_a(.in(in[13]), .out(far_0_532_0[0]));    relay_conn far_0_532_0_b(.in(in[99]), .out(far_0_532_0[1]));
    wire [1:0] far_0_532_1;    relay_conn far_0_532_1_a(.in(far_0_532_0[0]), .out(far_0_532_1[0]));    relay_conn far_0_532_1_b(.in(far_0_532_0[1]), .out(far_0_532_1[1]));
    assign layer_0[532] = far_0_532_1[1] & ~far_0_532_1[0]; 
    wire [1:0] far_0_533_0;    relay_conn far_0_533_0_a(.in(in[102]), .out(far_0_533_0[0]));    relay_conn far_0_533_0_b(.in(in[165]), .out(far_0_533_0[1]));
    assign layer_0[533] = far_0_533_0[1]; 
    wire [1:0] far_0_534_0;    relay_conn far_0_534_0_a(.in(in[74]), .out(far_0_534_0[0]));    relay_conn far_0_534_0_b(.in(in[157]), .out(far_0_534_0[1]));
    wire [1:0] far_0_534_1;    relay_conn far_0_534_1_a(.in(far_0_534_0[0]), .out(far_0_534_1[0]));    relay_conn far_0_534_1_b(.in(far_0_534_0[1]), .out(far_0_534_1[1]));
    assign layer_0[534] = ~far_0_534_1[0] | (far_0_534_1[0] & far_0_534_1[1]); 
    wire [1:0] far_0_535_0;    relay_conn far_0_535_0_a(.in(in[57]), .out(far_0_535_0[0]));    relay_conn far_0_535_0_b(.in(in[158]), .out(far_0_535_0[1]));
    wire [1:0] far_0_535_1;    relay_conn far_0_535_1_a(.in(far_0_535_0[0]), .out(far_0_535_1[0]));    relay_conn far_0_535_1_b(.in(far_0_535_0[1]), .out(far_0_535_1[1]));
    wire [1:0] far_0_535_2;    relay_conn far_0_535_2_a(.in(far_0_535_1[0]), .out(far_0_535_2[0]));    relay_conn far_0_535_2_b(.in(far_0_535_1[1]), .out(far_0_535_2[1]));
    assign layer_0[535] = far_0_535_2[1] & ~far_0_535_2[0]; 
    wire [1:0] far_0_536_0;    relay_conn far_0_536_0_a(.in(in[111]), .out(far_0_536_0[0]));    relay_conn far_0_536_0_b(.in(in[236]), .out(far_0_536_0[1]));
    wire [1:0] far_0_536_1;    relay_conn far_0_536_1_a(.in(far_0_536_0[0]), .out(far_0_536_1[0]));    relay_conn far_0_536_1_b(.in(far_0_536_0[1]), .out(far_0_536_1[1]));
    wire [1:0] far_0_536_2;    relay_conn far_0_536_2_a(.in(far_0_536_1[0]), .out(far_0_536_2[0]));    relay_conn far_0_536_2_b(.in(far_0_536_1[1]), .out(far_0_536_2[1]));
    assign layer_0[536] = far_0_536_2[0] | far_0_536_2[1]; 
    wire [1:0] far_0_537_0;    relay_conn far_0_537_0_a(.in(in[196]), .out(far_0_537_0[0]));    relay_conn far_0_537_0_b(.in(in[99]), .out(far_0_537_0[1]));
    wire [1:0] far_0_537_1;    relay_conn far_0_537_1_a(.in(far_0_537_0[0]), .out(far_0_537_1[0]));    relay_conn far_0_537_1_b(.in(far_0_537_0[1]), .out(far_0_537_1[1]));
    wire [1:0] far_0_537_2;    relay_conn far_0_537_2_a(.in(far_0_537_1[0]), .out(far_0_537_2[0]));    relay_conn far_0_537_2_b(.in(far_0_537_1[1]), .out(far_0_537_2[1]));
    assign layer_0[537] = far_0_537_2[1] & ~far_0_537_2[0]; 
    assign layer_0[538] = in[99] & ~in[113]; 
    wire [1:0] far_0_539_0;    relay_conn far_0_539_0_a(.in(in[195]), .out(far_0_539_0[0]));    relay_conn far_0_539_0_b(.in(in[233]), .out(far_0_539_0[1]));
    assign layer_0[539] = ~far_0_539_0[1]; 
    assign layer_0[540] = in[241] ^ in[223]; 
    wire [1:0] far_0_541_0;    relay_conn far_0_541_0_a(.in(in[221]), .out(far_0_541_0[0]));    relay_conn far_0_541_0_b(.in(in[136]), .out(far_0_541_0[1]));
    wire [1:0] far_0_541_1;    relay_conn far_0_541_1_a(.in(far_0_541_0[0]), .out(far_0_541_1[0]));    relay_conn far_0_541_1_b(.in(far_0_541_0[1]), .out(far_0_541_1[1]));
    assign layer_0[541] = far_0_541_1[1]; 
    wire [1:0] far_0_542_0;    relay_conn far_0_542_0_a(.in(in[202]), .out(far_0_542_0[0]));    relay_conn far_0_542_0_b(.in(in[120]), .out(far_0_542_0[1]));
    wire [1:0] far_0_542_1;    relay_conn far_0_542_1_a(.in(far_0_542_0[0]), .out(far_0_542_1[0]));    relay_conn far_0_542_1_b(.in(far_0_542_0[1]), .out(far_0_542_1[1]));
    assign layer_0[542] = ~far_0_542_1[0]; 
    assign layer_0[543] = in[187] & ~in[182]; 
    wire [1:0] far_0_544_0;    relay_conn far_0_544_0_a(.in(in[239]), .out(far_0_544_0[0]));    relay_conn far_0_544_0_b(.in(in[207]), .out(far_0_544_0[1]));
    assign layer_0[544] = ~(far_0_544_0[0] ^ far_0_544_0[1]); 
    wire [1:0] far_0_545_0;    relay_conn far_0_545_0_a(.in(in[157]), .out(far_0_545_0[0]));    relay_conn far_0_545_0_b(.in(in[43]), .out(far_0_545_0[1]));
    wire [1:0] far_0_545_1;    relay_conn far_0_545_1_a(.in(far_0_545_0[0]), .out(far_0_545_1[0]));    relay_conn far_0_545_1_b(.in(far_0_545_0[1]), .out(far_0_545_1[1]));
    wire [1:0] far_0_545_2;    relay_conn far_0_545_2_a(.in(far_0_545_1[0]), .out(far_0_545_2[0]));    relay_conn far_0_545_2_b(.in(far_0_545_1[1]), .out(far_0_545_2[1]));
    assign layer_0[545] = ~far_0_545_2[0]; 
    assign layer_0[546] = ~(in[57] ^ in[28]); 
    assign layer_0[547] = ~(in[42] | in[43]); 
    wire [1:0] far_0_548_0;    relay_conn far_0_548_0_a(.in(in[181]), .out(far_0_548_0[0]));    relay_conn far_0_548_0_b(.in(in[215]), .out(far_0_548_0[1]));
    assign layer_0[548] = ~far_0_548_0[0]; 
    assign layer_0[549] = ~in[132]; 
    wire [1:0] far_0_550_0;    relay_conn far_0_550_0_a(.in(in[71]), .out(far_0_550_0[0]));    relay_conn far_0_550_0_b(.in(in[165]), .out(far_0_550_0[1]));
    wire [1:0] far_0_550_1;    relay_conn far_0_550_1_a(.in(far_0_550_0[0]), .out(far_0_550_1[0]));    relay_conn far_0_550_1_b(.in(far_0_550_0[1]), .out(far_0_550_1[1]));
    assign layer_0[550] = far_0_550_1[0] | far_0_550_1[1]; 
    wire [1:0] far_0_551_0;    relay_conn far_0_551_0_a(.in(in[196]), .out(far_0_551_0[0]));    relay_conn far_0_551_0_b(.in(in[236]), .out(far_0_551_0[1]));
    assign layer_0[551] = ~far_0_551_0[1]; 
    wire [1:0] far_0_552_0;    relay_conn far_0_552_0_a(.in(in[115]), .out(far_0_552_0[0]));    relay_conn far_0_552_0_b(.in(in[165]), .out(far_0_552_0[1]));
    assign layer_0[552] = far_0_552_0[1]; 
    wire [1:0] far_0_553_0;    relay_conn far_0_553_0_a(.in(in[247]), .out(far_0_553_0[0]));    relay_conn far_0_553_0_b(.in(in[151]), .out(far_0_553_0[1]));
    wire [1:0] far_0_553_1;    relay_conn far_0_553_1_a(.in(far_0_553_0[0]), .out(far_0_553_1[0]));    relay_conn far_0_553_1_b(.in(far_0_553_0[1]), .out(far_0_553_1[1]));
    wire [1:0] far_0_553_2;    relay_conn far_0_553_2_a(.in(far_0_553_1[0]), .out(far_0_553_2[0]));    relay_conn far_0_553_2_b(.in(far_0_553_1[1]), .out(far_0_553_2[1]));
    assign layer_0[553] = ~far_0_553_2[0] | (far_0_553_2[0] & far_0_553_2[1]); 
    wire [1:0] far_0_554_0;    relay_conn far_0_554_0_a(.in(in[87]), .out(far_0_554_0[0]));    relay_conn far_0_554_0_b(.in(in[214]), .out(far_0_554_0[1]));
    wire [1:0] far_0_554_1;    relay_conn far_0_554_1_a(.in(far_0_554_0[0]), .out(far_0_554_1[0]));    relay_conn far_0_554_1_b(.in(far_0_554_0[1]), .out(far_0_554_1[1]));
    wire [1:0] far_0_554_2;    relay_conn far_0_554_2_a(.in(far_0_554_1[0]), .out(far_0_554_2[0]));    relay_conn far_0_554_2_b(.in(far_0_554_1[1]), .out(far_0_554_2[1]));
    assign layer_0[554] = far_0_554_2[0] | far_0_554_2[1]; 
    wire [1:0] far_0_555_0;    relay_conn far_0_555_0_a(.in(in[199]), .out(far_0_555_0[0]));    relay_conn far_0_555_0_b(.in(in[132]), .out(far_0_555_0[1]));
    wire [1:0] far_0_555_1;    relay_conn far_0_555_1_a(.in(far_0_555_0[0]), .out(far_0_555_1[0]));    relay_conn far_0_555_1_b(.in(far_0_555_0[1]), .out(far_0_555_1[1]));
    assign layer_0[555] = far_0_555_1[0] | far_0_555_1[1]; 
    wire [1:0] far_0_556_0;    relay_conn far_0_556_0_a(.in(in[61]), .out(far_0_556_0[0]));    relay_conn far_0_556_0_b(.in(in[157]), .out(far_0_556_0[1]));
    wire [1:0] far_0_556_1;    relay_conn far_0_556_1_a(.in(far_0_556_0[0]), .out(far_0_556_1[0]));    relay_conn far_0_556_1_b(.in(far_0_556_0[1]), .out(far_0_556_1[1]));
    wire [1:0] far_0_556_2;    relay_conn far_0_556_2_a(.in(far_0_556_1[0]), .out(far_0_556_2[0]));    relay_conn far_0_556_2_b(.in(far_0_556_1[1]), .out(far_0_556_2[1]));
    assign layer_0[556] = ~far_0_556_2[1] | (far_0_556_2[0] & far_0_556_2[1]); 
    assign layer_0[557] = ~in[88] | (in[116] & in[88]); 
    assign layer_0[558] = ~in[5] | (in[5] & in[6]); 
    assign layer_0[559] = ~in[51] | (in[48] & in[51]); 
    wire [1:0] far_0_560_0;    relay_conn far_0_560_0_a(.in(in[125]), .out(far_0_560_0[0]));    relay_conn far_0_560_0_b(.in(in[199]), .out(far_0_560_0[1]));
    wire [1:0] far_0_560_1;    relay_conn far_0_560_1_a(.in(far_0_560_0[0]), .out(far_0_560_1[0]));    relay_conn far_0_560_1_b(.in(far_0_560_0[1]), .out(far_0_560_1[1]));
    assign layer_0[560] = ~(far_0_560_1[0] | far_0_560_1[1]); 
    wire [1:0] far_0_561_0;    relay_conn far_0_561_0_a(.in(in[99]), .out(far_0_561_0[0]));    relay_conn far_0_561_0_b(.in(in[158]), .out(far_0_561_0[1]));
    assign layer_0[561] = far_0_561_0[0] | far_0_561_0[1]; 
    assign layer_0[562] = ~(in[88] | in[79]); 
    wire [1:0] far_0_563_0;    relay_conn far_0_563_0_a(.in(in[54]), .out(far_0_563_0[0]));    relay_conn far_0_563_0_b(.in(in[127]), .out(far_0_563_0[1]));
    wire [1:0] far_0_563_1;    relay_conn far_0_563_1_a(.in(far_0_563_0[0]), .out(far_0_563_1[0]));    relay_conn far_0_563_1_b(.in(far_0_563_0[1]), .out(far_0_563_1[1]));
    assign layer_0[563] = far_0_563_1[1]; 
    wire [1:0] far_0_564_0;    relay_conn far_0_564_0_a(.in(in[24]), .out(far_0_564_0[0]));    relay_conn far_0_564_0_b(.in(in[121]), .out(far_0_564_0[1]));
    wire [1:0] far_0_564_1;    relay_conn far_0_564_1_a(.in(far_0_564_0[0]), .out(far_0_564_1[0]));    relay_conn far_0_564_1_b(.in(far_0_564_0[1]), .out(far_0_564_1[1]));
    wire [1:0] far_0_564_2;    relay_conn far_0_564_2_a(.in(far_0_564_1[0]), .out(far_0_564_2[0]));    relay_conn far_0_564_2_b(.in(far_0_564_1[1]), .out(far_0_564_2[1]));
    assign layer_0[564] = ~(far_0_564_2[0] & far_0_564_2[1]); 
    wire [1:0] far_0_565_0;    relay_conn far_0_565_0_a(.in(in[215]), .out(far_0_565_0[0]));    relay_conn far_0_565_0_b(.in(in[117]), .out(far_0_565_0[1]));
    wire [1:0] far_0_565_1;    relay_conn far_0_565_1_a(.in(far_0_565_0[0]), .out(far_0_565_1[0]));    relay_conn far_0_565_1_b(.in(far_0_565_0[1]), .out(far_0_565_1[1]));
    wire [1:0] far_0_565_2;    relay_conn far_0_565_2_a(.in(far_0_565_1[0]), .out(far_0_565_2[0]));    relay_conn far_0_565_2_b(.in(far_0_565_1[1]), .out(far_0_565_2[1]));
    assign layer_0[565] = ~far_0_565_2[1]; 
    wire [1:0] far_0_566_0;    relay_conn far_0_566_0_a(.in(in[38]), .out(far_0_566_0[0]));    relay_conn far_0_566_0_b(.in(in[135]), .out(far_0_566_0[1]));
    wire [1:0] far_0_566_1;    relay_conn far_0_566_1_a(.in(far_0_566_0[0]), .out(far_0_566_1[0]));    relay_conn far_0_566_1_b(.in(far_0_566_0[1]), .out(far_0_566_1[1]));
    wire [1:0] far_0_566_2;    relay_conn far_0_566_2_a(.in(far_0_566_1[0]), .out(far_0_566_2[0]));    relay_conn far_0_566_2_b(.in(far_0_566_1[1]), .out(far_0_566_2[1]));
    assign layer_0[566] = ~far_0_566_2[0]; 
    wire [1:0] far_0_567_0;    relay_conn far_0_567_0_a(.in(in[61]), .out(far_0_567_0[0]));    relay_conn far_0_567_0_b(.in(in[111]), .out(far_0_567_0[1]));
    assign layer_0[567] = far_0_567_0[1]; 
    assign layer_0[568] = in[198]; 
    assign layer_0[569] = in[172] & ~in[198]; 
    wire [1:0] far_0_570_0;    relay_conn far_0_570_0_a(.in(in[215]), .out(far_0_570_0[0]));    relay_conn far_0_570_0_b(.in(in[117]), .out(far_0_570_0[1]));
    wire [1:0] far_0_570_1;    relay_conn far_0_570_1_a(.in(far_0_570_0[0]), .out(far_0_570_1[0]));    relay_conn far_0_570_1_b(.in(far_0_570_0[1]), .out(far_0_570_1[1]));
    wire [1:0] far_0_570_2;    relay_conn far_0_570_2_a(.in(far_0_570_1[0]), .out(far_0_570_2[0]));    relay_conn far_0_570_2_b(.in(far_0_570_1[1]), .out(far_0_570_2[1]));
    assign layer_0[570] = far_0_570_2[0] ^ far_0_570_2[1]; 
    assign layer_0[571] = ~(in[233] & in[250]); 
    wire [1:0] far_0_572_0;    relay_conn far_0_572_0_a(.in(in[179]), .out(far_0_572_0[0]));    relay_conn far_0_572_0_b(.in(in[121]), .out(far_0_572_0[1]));
    assign layer_0[572] = ~far_0_572_0[1]; 
    wire [1:0] far_0_573_0;    relay_conn far_0_573_0_a(.in(in[137]), .out(far_0_573_0[0]));    relay_conn far_0_573_0_b(.in(in[202]), .out(far_0_573_0[1]));
    wire [1:0] far_0_573_1;    relay_conn far_0_573_1_a(.in(far_0_573_0[0]), .out(far_0_573_1[0]));    relay_conn far_0_573_1_b(.in(far_0_573_0[1]), .out(far_0_573_1[1]));
    assign layer_0[573] = far_0_573_1[0]; 
    assign layer_0[574] = ~(in[171] | in[151]); 
    wire [1:0] far_0_575_0;    relay_conn far_0_575_0_a(.in(in[157]), .out(far_0_575_0[0]));    relay_conn far_0_575_0_b(.in(in[101]), .out(far_0_575_0[1]));
    assign layer_0[575] = ~(far_0_575_0[0] | far_0_575_0[1]); 
    wire [1:0] far_0_576_0;    relay_conn far_0_576_0_a(.in(in[157]), .out(far_0_576_0[0]));    relay_conn far_0_576_0_b(.in(in[97]), .out(far_0_576_0[1]));
    assign layer_0[576] = ~(far_0_576_0[0] ^ far_0_576_0[1]); 
    wire [1:0] far_0_577_0;    relay_conn far_0_577_0_a(.in(in[196]), .out(far_0_577_0[0]));    relay_conn far_0_577_0_b(.in(in[151]), .out(far_0_577_0[1]));
    assign layer_0[577] = far_0_577_0[1]; 
    wire [1:0] far_0_578_0;    relay_conn far_0_578_0_a(.in(in[182]), .out(far_0_578_0[0]));    relay_conn far_0_578_0_b(.in(in[240]), .out(far_0_578_0[1]));
    assign layer_0[578] = ~far_0_578_0[1]; 
    wire [1:0] far_0_579_0;    relay_conn far_0_579_0_a(.in(in[31]), .out(far_0_579_0[0]));    relay_conn far_0_579_0_b(.in(in[142]), .out(far_0_579_0[1]));
    wire [1:0] far_0_579_1;    relay_conn far_0_579_1_a(.in(far_0_579_0[0]), .out(far_0_579_1[0]));    relay_conn far_0_579_1_b(.in(far_0_579_0[1]), .out(far_0_579_1[1]));
    wire [1:0] far_0_579_2;    relay_conn far_0_579_2_a(.in(far_0_579_1[0]), .out(far_0_579_2[0]));    relay_conn far_0_579_2_b(.in(far_0_579_1[1]), .out(far_0_579_2[1]));
    assign layer_0[579] = far_0_579_2[0] & ~far_0_579_2[1]; 
    wire [1:0] far_0_580_0;    relay_conn far_0_580_0_a(.in(in[157]), .out(far_0_580_0[0]));    relay_conn far_0_580_0_b(.in(in[102]), .out(far_0_580_0[1]));
    assign layer_0[580] = far_0_580_0[1] & ~far_0_580_0[0]; 
    wire [1:0] far_0_581_0;    relay_conn far_0_581_0_a(.in(in[229]), .out(far_0_581_0[0]));    relay_conn far_0_581_0_b(.in(in[158]), .out(far_0_581_0[1]));
    wire [1:0] far_0_581_1;    relay_conn far_0_581_1_a(.in(far_0_581_0[0]), .out(far_0_581_1[0]));    relay_conn far_0_581_1_b(.in(far_0_581_0[1]), .out(far_0_581_1[1]));
    assign layer_0[581] = far_0_581_1[0]; 
    assign layer_0[582] = ~in[201]; 
    assign layer_0[583] = in[211] & in[238]; 
    wire [1:0] far_0_584_0;    relay_conn far_0_584_0_a(.in(in[122]), .out(far_0_584_0[0]));    relay_conn far_0_584_0_b(.in(in[15]), .out(far_0_584_0[1]));
    wire [1:0] far_0_584_1;    relay_conn far_0_584_1_a(.in(far_0_584_0[0]), .out(far_0_584_1[0]));    relay_conn far_0_584_1_b(.in(far_0_584_0[1]), .out(far_0_584_1[1]));
    wire [1:0] far_0_584_2;    relay_conn far_0_584_2_a(.in(far_0_584_1[0]), .out(far_0_584_2[0]));    relay_conn far_0_584_2_b(.in(far_0_584_1[1]), .out(far_0_584_2[1]));
    assign layer_0[584] = far_0_584_2[0]; 
    wire [1:0] far_0_585_0;    relay_conn far_0_585_0_a(.in(in[212]), .out(far_0_585_0[0]));    relay_conn far_0_585_0_b(.in(in[105]), .out(far_0_585_0[1]));
    wire [1:0] far_0_585_1;    relay_conn far_0_585_1_a(.in(far_0_585_0[0]), .out(far_0_585_1[0]));    relay_conn far_0_585_1_b(.in(far_0_585_0[1]), .out(far_0_585_1[1]));
    wire [1:0] far_0_585_2;    relay_conn far_0_585_2_a(.in(far_0_585_1[0]), .out(far_0_585_2[0]));    relay_conn far_0_585_2_b(.in(far_0_585_1[1]), .out(far_0_585_2[1]));
    assign layer_0[585] = ~far_0_585_2[0] | (far_0_585_2[0] & far_0_585_2[1]); 
    wire [1:0] far_0_586_0;    relay_conn far_0_586_0_a(.in(in[3]), .out(far_0_586_0[0]));    relay_conn far_0_586_0_b(.in(in[88]), .out(far_0_586_0[1]));
    wire [1:0] far_0_586_1;    relay_conn far_0_586_1_a(.in(far_0_586_0[0]), .out(far_0_586_1[0]));    relay_conn far_0_586_1_b(.in(far_0_586_0[1]), .out(far_0_586_1[1]));
    assign layer_0[586] = far_0_586_1[1] & ~far_0_586_1[0]; 
    assign layer_0[587] = in[211] | in[201]; 
    wire [1:0] far_0_588_0;    relay_conn far_0_588_0_a(.in(in[10]), .out(far_0_588_0[0]));    relay_conn far_0_588_0_b(.in(in[70]), .out(far_0_588_0[1]));
    assign layer_0[588] = ~(far_0_588_0[0] | far_0_588_0[1]); 
    wire [1:0] far_0_589_0;    relay_conn far_0_589_0_a(.in(in[159]), .out(far_0_589_0[0]));    relay_conn far_0_589_0_b(.in(in[37]), .out(far_0_589_0[1]));
    wire [1:0] far_0_589_1;    relay_conn far_0_589_1_a(.in(far_0_589_0[0]), .out(far_0_589_1[0]));    relay_conn far_0_589_1_b(.in(far_0_589_0[1]), .out(far_0_589_1[1]));
    wire [1:0] far_0_589_2;    relay_conn far_0_589_2_a(.in(far_0_589_1[0]), .out(far_0_589_2[0]));    relay_conn far_0_589_2_b(.in(far_0_589_1[1]), .out(far_0_589_2[1]));
    assign layer_0[589] = far_0_589_2[0] & far_0_589_2[1]; 
    wire [1:0] far_0_590_0;    relay_conn far_0_590_0_a(.in(in[208]), .out(far_0_590_0[0]));    relay_conn far_0_590_0_b(.in(in[109]), .out(far_0_590_0[1]));
    wire [1:0] far_0_590_1;    relay_conn far_0_590_1_a(.in(far_0_590_0[0]), .out(far_0_590_1[0]));    relay_conn far_0_590_1_b(.in(far_0_590_0[1]), .out(far_0_590_1[1]));
    wire [1:0] far_0_590_2;    relay_conn far_0_590_2_a(.in(far_0_590_1[0]), .out(far_0_590_2[0]));    relay_conn far_0_590_2_b(.in(far_0_590_1[1]), .out(far_0_590_2[1]));
    assign layer_0[590] = ~far_0_590_2[0] | (far_0_590_2[0] & far_0_590_2[1]); 
    wire [1:0] far_0_591_0;    relay_conn far_0_591_0_a(.in(in[151]), .out(far_0_591_0[0]));    relay_conn far_0_591_0_b(.in(in[117]), .out(far_0_591_0[1]));
    assign layer_0[591] = ~(far_0_591_0[0] ^ far_0_591_0[1]); 
    wire [1:0] far_0_592_0;    relay_conn far_0_592_0_a(.in(in[111]), .out(far_0_592_0[0]));    relay_conn far_0_592_0_b(.in(in[72]), .out(far_0_592_0[1]));
    assign layer_0[592] = ~(far_0_592_0[0] & far_0_592_0[1]); 
    wire [1:0] far_0_593_0;    relay_conn far_0_593_0_a(.in(in[132]), .out(far_0_593_0[0]));    relay_conn far_0_593_0_b(.in(in[10]), .out(far_0_593_0[1]));
    wire [1:0] far_0_593_1;    relay_conn far_0_593_1_a(.in(far_0_593_0[0]), .out(far_0_593_1[0]));    relay_conn far_0_593_1_b(.in(far_0_593_0[1]), .out(far_0_593_1[1]));
    wire [1:0] far_0_593_2;    relay_conn far_0_593_2_a(.in(far_0_593_1[0]), .out(far_0_593_2[0]));    relay_conn far_0_593_2_b(.in(far_0_593_1[1]), .out(far_0_593_2[1]));
    assign layer_0[593] = far_0_593_2[1] & ~far_0_593_2[0]; 
    wire [1:0] far_0_594_0;    relay_conn far_0_594_0_a(.in(in[136]), .out(far_0_594_0[0]));    relay_conn far_0_594_0_b(.in(in[96]), .out(far_0_594_0[1]));
    assign layer_0[594] = ~(far_0_594_0[0] & far_0_594_0[1]); 
    assign layer_0[595] = in[233] & in[239]; 
    wire [1:0] far_0_596_0;    relay_conn far_0_596_0_a(.in(in[219]), .out(far_0_596_0[0]));    relay_conn far_0_596_0_b(.in(in[125]), .out(far_0_596_0[1]));
    wire [1:0] far_0_596_1;    relay_conn far_0_596_1_a(.in(far_0_596_0[0]), .out(far_0_596_1[0]));    relay_conn far_0_596_1_b(.in(far_0_596_0[1]), .out(far_0_596_1[1]));
    assign layer_0[596] = far_0_596_1[0] & far_0_596_1[1]; 
    wire [1:0] far_0_597_0;    relay_conn far_0_597_0_a(.in(in[77]), .out(far_0_597_0[0]));    relay_conn far_0_597_0_b(.in(in[149]), .out(far_0_597_0[1]));
    wire [1:0] far_0_597_1;    relay_conn far_0_597_1_a(.in(far_0_597_0[0]), .out(far_0_597_1[0]));    relay_conn far_0_597_1_b(.in(far_0_597_0[1]), .out(far_0_597_1[1]));
    assign layer_0[597] = ~far_0_597_1[0]; 
    wire [1:0] far_0_598_0;    relay_conn far_0_598_0_a(.in(in[95]), .out(far_0_598_0[0]));    relay_conn far_0_598_0_b(.in(in[135]), .out(far_0_598_0[1]));
    assign layer_0[598] = far_0_598_0[0] & far_0_598_0[1]; 
    wire [1:0] far_0_599_0;    relay_conn far_0_599_0_a(.in(in[125]), .out(far_0_599_0[0]));    relay_conn far_0_599_0_b(.in(in[28]), .out(far_0_599_0[1]));
    wire [1:0] far_0_599_1;    relay_conn far_0_599_1_a(.in(far_0_599_0[0]), .out(far_0_599_1[0]));    relay_conn far_0_599_1_b(.in(far_0_599_0[1]), .out(far_0_599_1[1]));
    wire [1:0] far_0_599_2;    relay_conn far_0_599_2_a(.in(far_0_599_1[0]), .out(far_0_599_2[0]));    relay_conn far_0_599_2_b(.in(far_0_599_1[1]), .out(far_0_599_2[1]));
    assign layer_0[599] = ~far_0_599_2[0] | (far_0_599_2[0] & far_0_599_2[1]); 
    assign layer_0[600] = ~in[105]; 
    wire [1:0] far_0_601_0;    relay_conn far_0_601_0_a(.in(in[101]), .out(far_0_601_0[0]));    relay_conn far_0_601_0_b(.in(in[151]), .out(far_0_601_0[1]));
    assign layer_0[601] = ~(far_0_601_0[0] & far_0_601_0[1]); 
    assign layer_0[602] = ~in[132]; 
    wire [1:0] far_0_603_0;    relay_conn far_0_603_0_a(.in(in[187]), .out(far_0_603_0[0]));    relay_conn far_0_603_0_b(.in(in[155]), .out(far_0_603_0[1]));
    assign layer_0[603] = far_0_603_0[0] ^ far_0_603_0[1]; 
    assign layer_0[604] = ~(in[110] & in[115]); 
    assign layer_0[605] = in[53] ^ in[67]; 
    wire [1:0] far_0_606_0;    relay_conn far_0_606_0_a(.in(in[43]), .out(far_0_606_0[0]));    relay_conn far_0_606_0_b(.in(in[95]), .out(far_0_606_0[1]));
    assign layer_0[606] = ~far_0_606_0[0]; 
    wire [1:0] far_0_607_0;    relay_conn far_0_607_0_a(.in(in[89]), .out(far_0_607_0[0]));    relay_conn far_0_607_0_b(.in(in[0]), .out(far_0_607_0[1]));
    wire [1:0] far_0_607_1;    relay_conn far_0_607_1_a(.in(far_0_607_0[0]), .out(far_0_607_1[0]));    relay_conn far_0_607_1_b(.in(far_0_607_0[1]), .out(far_0_607_1[1]));
    assign layer_0[607] = ~far_0_607_1[1]; 
    assign layer_0[608] = ~in[181]; 
    assign layer_0[609] = ~(in[101] | in[82]); 
    wire [1:0] far_0_610_0;    relay_conn far_0_610_0_a(.in(in[202]), .out(far_0_610_0[0]));    relay_conn far_0_610_0_b(.in(in[81]), .out(far_0_610_0[1]));
    wire [1:0] far_0_610_1;    relay_conn far_0_610_1_a(.in(far_0_610_0[0]), .out(far_0_610_1[0]));    relay_conn far_0_610_1_b(.in(far_0_610_0[1]), .out(far_0_610_1[1]));
    wire [1:0] far_0_610_2;    relay_conn far_0_610_2_a(.in(far_0_610_1[0]), .out(far_0_610_2[0]));    relay_conn far_0_610_2_b(.in(far_0_610_1[1]), .out(far_0_610_2[1]));
    assign layer_0[610] = far_0_610_2[1]; 
    assign layer_0[611] = in[182]; 
    assign layer_0[612] = in[158] | in[151]; 
    wire [1:0] far_0_613_0;    relay_conn far_0_613_0_a(.in(in[181]), .out(far_0_613_0[0]));    relay_conn far_0_613_0_b(.in(in[125]), .out(far_0_613_0[1]));
    assign layer_0[613] = far_0_613_0[0] ^ far_0_613_0[1]; 
    wire [1:0] far_0_614_0;    relay_conn far_0_614_0_a(.in(in[195]), .out(far_0_614_0[0]));    relay_conn far_0_614_0_b(.in(in[102]), .out(far_0_614_0[1]));
    wire [1:0] far_0_614_1;    relay_conn far_0_614_1_a(.in(far_0_614_0[0]), .out(far_0_614_1[0]));    relay_conn far_0_614_1_b(.in(far_0_614_0[1]), .out(far_0_614_1[1]));
    assign layer_0[614] = ~(far_0_614_1[0] & far_0_614_1[1]); 
    wire [1:0] far_0_615_0;    relay_conn far_0_615_0_a(.in(in[109]), .out(far_0_615_0[0]));    relay_conn far_0_615_0_b(.in(in[195]), .out(far_0_615_0[1]));
    wire [1:0] far_0_615_1;    relay_conn far_0_615_1_a(.in(far_0_615_0[0]), .out(far_0_615_1[0]));    relay_conn far_0_615_1_b(.in(far_0_615_0[1]), .out(far_0_615_1[1]));
    assign layer_0[615] = far_0_615_1[1]; 
    wire [1:0] far_0_616_0;    relay_conn far_0_616_0_a(.in(in[113]), .out(far_0_616_0[0]));    relay_conn far_0_616_0_b(.in(in[215]), .out(far_0_616_0[1]));
    wire [1:0] far_0_616_1;    relay_conn far_0_616_1_a(.in(far_0_616_0[0]), .out(far_0_616_1[0]));    relay_conn far_0_616_1_b(.in(far_0_616_0[1]), .out(far_0_616_1[1]));
    wire [1:0] far_0_616_2;    relay_conn far_0_616_2_a(.in(far_0_616_1[0]), .out(far_0_616_2[0]));    relay_conn far_0_616_2_b(.in(far_0_616_1[1]), .out(far_0_616_2[1]));
    assign layer_0[616] = ~far_0_616_2[1]; 
    assign layer_0[617] = ~in[88] | (in[74] & in[88]); 
    wire [1:0] far_0_618_0;    relay_conn far_0_618_0_a(.in(in[145]), .out(far_0_618_0[0]));    relay_conn far_0_618_0_b(.in(in[55]), .out(far_0_618_0[1]));
    wire [1:0] far_0_618_1;    relay_conn far_0_618_1_a(.in(far_0_618_0[0]), .out(far_0_618_1[0]));    relay_conn far_0_618_1_b(.in(far_0_618_0[1]), .out(far_0_618_1[1]));
    assign layer_0[618] = ~far_0_618_1[0] | (far_0_618_1[0] & far_0_618_1[1]); 
    wire [1:0] far_0_619_0;    relay_conn far_0_619_0_a(.in(in[76]), .out(far_0_619_0[0]));    relay_conn far_0_619_0_b(.in(in[197]), .out(far_0_619_0[1]));
    wire [1:0] far_0_619_1;    relay_conn far_0_619_1_a(.in(far_0_619_0[0]), .out(far_0_619_1[0]));    relay_conn far_0_619_1_b(.in(far_0_619_0[1]), .out(far_0_619_1[1]));
    wire [1:0] far_0_619_2;    relay_conn far_0_619_2_a(.in(far_0_619_1[0]), .out(far_0_619_2[0]));    relay_conn far_0_619_2_b(.in(far_0_619_1[1]), .out(far_0_619_2[1]));
    assign layer_0[619] = far_0_619_2[0] & ~far_0_619_2[1]; 
    wire [1:0] far_0_620_0;    relay_conn far_0_620_0_a(.in(in[230]), .out(far_0_620_0[0]));    relay_conn far_0_620_0_b(.in(in[138]), .out(far_0_620_0[1]));
    wire [1:0] far_0_620_1;    relay_conn far_0_620_1_a(.in(far_0_620_0[0]), .out(far_0_620_1[0]));    relay_conn far_0_620_1_b(.in(far_0_620_0[1]), .out(far_0_620_1[1]));
    assign layer_0[620] = far_0_620_1[1]; 
    wire [1:0] far_0_621_0;    relay_conn far_0_621_0_a(.in(in[83]), .out(far_0_621_0[0]));    relay_conn far_0_621_0_b(.in(in[188]), .out(far_0_621_0[1]));
    wire [1:0] far_0_621_1;    relay_conn far_0_621_1_a(.in(far_0_621_0[0]), .out(far_0_621_1[0]));    relay_conn far_0_621_1_b(.in(far_0_621_0[1]), .out(far_0_621_1[1]));
    wire [1:0] far_0_621_2;    relay_conn far_0_621_2_a(.in(far_0_621_1[0]), .out(far_0_621_2[0]));    relay_conn far_0_621_2_b(.in(far_0_621_1[1]), .out(far_0_621_2[1]));
    assign layer_0[621] = far_0_621_2[0] & far_0_621_2[1]; 
    wire [1:0] far_0_622_0;    relay_conn far_0_622_0_a(.in(in[15]), .out(far_0_622_0[0]));    relay_conn far_0_622_0_b(.in(in[75]), .out(far_0_622_0[1]));
    assign layer_0[622] = ~(far_0_622_0[0] | far_0_622_0[1]); 
    wire [1:0] far_0_623_0;    relay_conn far_0_623_0_a(.in(in[241]), .out(far_0_623_0[0]));    relay_conn far_0_623_0_b(.in(in[149]), .out(far_0_623_0[1]));
    wire [1:0] far_0_623_1;    relay_conn far_0_623_1_a(.in(far_0_623_0[0]), .out(far_0_623_1[0]));    relay_conn far_0_623_1_b(.in(far_0_623_0[1]), .out(far_0_623_1[1]));
    assign layer_0[623] = ~(far_0_623_1[0] ^ far_0_623_1[1]); 
    wire [1:0] far_0_624_0;    relay_conn far_0_624_0_a(.in(in[157]), .out(far_0_624_0[0]));    relay_conn far_0_624_0_b(.in(in[241]), .out(far_0_624_0[1]));
    wire [1:0] far_0_624_1;    relay_conn far_0_624_1_a(.in(far_0_624_0[0]), .out(far_0_624_1[0]));    relay_conn far_0_624_1_b(.in(far_0_624_0[1]), .out(far_0_624_1[1]));
    assign layer_0[624] = ~far_0_624_1[0] | (far_0_624_1[0] & far_0_624_1[1]); 
    wire [1:0] far_0_625_0;    relay_conn far_0_625_0_a(.in(in[3]), .out(far_0_625_0[0]));    relay_conn far_0_625_0_b(.in(in[43]), .out(far_0_625_0[1]));
    assign layer_0[625] = ~far_0_625_0[1] | (far_0_625_0[0] & far_0_625_0[1]); 
    wire [1:0] far_0_626_0;    relay_conn far_0_626_0_a(.in(in[245]), .out(far_0_626_0[0]));    relay_conn far_0_626_0_b(.in(in[136]), .out(far_0_626_0[1]));
    wire [1:0] far_0_626_1;    relay_conn far_0_626_1_a(.in(far_0_626_0[0]), .out(far_0_626_1[0]));    relay_conn far_0_626_1_b(.in(far_0_626_0[1]), .out(far_0_626_1[1]));
    wire [1:0] far_0_626_2;    relay_conn far_0_626_2_a(.in(far_0_626_1[0]), .out(far_0_626_2[0]));    relay_conn far_0_626_2_b(.in(far_0_626_1[1]), .out(far_0_626_2[1]));
    assign layer_0[626] = ~(far_0_626_2[0] & far_0_626_2[1]); 
    wire [1:0] far_0_627_0;    relay_conn far_0_627_0_a(.in(in[157]), .out(far_0_627_0[0]));    relay_conn far_0_627_0_b(.in(in[125]), .out(far_0_627_0[1]));
    assign layer_0[627] = far_0_627_0[0] & ~far_0_627_0[1]; 
    wire [1:0] far_0_628_0;    relay_conn far_0_628_0_a(.in(in[135]), .out(far_0_628_0[0]));    relay_conn far_0_628_0_b(.in(in[82]), .out(far_0_628_0[1]));
    assign layer_0[628] = ~far_0_628_0[1]; 
    wire [1:0] far_0_629_0;    relay_conn far_0_629_0_a(.in(in[125]), .out(far_0_629_0[0]));    relay_conn far_0_629_0_b(.in(in[199]), .out(far_0_629_0[1]));
    wire [1:0] far_0_629_1;    relay_conn far_0_629_1_a(.in(far_0_629_0[0]), .out(far_0_629_1[0]));    relay_conn far_0_629_1_b(.in(far_0_629_0[1]), .out(far_0_629_1[1]));
    assign layer_0[629] = ~far_0_629_1[1]; 
    assign layer_0[630] = in[66] & in[76]; 
    wire [1:0] far_0_631_0;    relay_conn far_0_631_0_a(.in(in[214]), .out(far_0_631_0[0]));    relay_conn far_0_631_0_b(.in(in[139]), .out(far_0_631_0[1]));
    wire [1:0] far_0_631_1;    relay_conn far_0_631_1_a(.in(far_0_631_0[0]), .out(far_0_631_1[0]));    relay_conn far_0_631_1_b(.in(far_0_631_0[1]), .out(far_0_631_1[1]));
    assign layer_0[631] = far_0_631_1[1] & ~far_0_631_1[0]; 
    wire [1:0] far_0_632_0;    relay_conn far_0_632_0_a(.in(in[0]), .out(far_0_632_0[0]));    relay_conn far_0_632_0_b(.in(in[44]), .out(far_0_632_0[1]));
    assign layer_0[632] = far_0_632_0[0] & far_0_632_0[1]; 
    wire [1:0] far_0_633_0;    relay_conn far_0_633_0_a(.in(in[243]), .out(far_0_633_0[0]));    relay_conn far_0_633_0_b(.in(in[150]), .out(far_0_633_0[1]));
    wire [1:0] far_0_633_1;    relay_conn far_0_633_1_a(.in(far_0_633_0[0]), .out(far_0_633_1[0]));    relay_conn far_0_633_1_b(.in(far_0_633_0[1]), .out(far_0_633_1[1]));
    assign layer_0[633] = ~far_0_633_1[0] | (far_0_633_1[0] & far_0_633_1[1]); 
    wire [1:0] far_0_634_0;    relay_conn far_0_634_0_a(.in(in[0]), .out(far_0_634_0[0]));    relay_conn far_0_634_0_b(.in(in[97]), .out(far_0_634_0[1]));
    wire [1:0] far_0_634_1;    relay_conn far_0_634_1_a(.in(far_0_634_0[0]), .out(far_0_634_1[0]));    relay_conn far_0_634_1_b(.in(far_0_634_0[1]), .out(far_0_634_1[1]));
    wire [1:0] far_0_634_2;    relay_conn far_0_634_2_a(.in(far_0_634_1[0]), .out(far_0_634_2[0]));    relay_conn far_0_634_2_b(.in(far_0_634_1[1]), .out(far_0_634_2[1]));
    assign layer_0[634] = ~(far_0_634_2[0] | far_0_634_2[1]); 
    wire [1:0] far_0_635_0;    relay_conn far_0_635_0_a(.in(in[113]), .out(far_0_635_0[0]));    relay_conn far_0_635_0_b(.in(in[195]), .out(far_0_635_0[1]));
    wire [1:0] far_0_635_1;    relay_conn far_0_635_1_a(.in(far_0_635_0[0]), .out(far_0_635_1[0]));    relay_conn far_0_635_1_b(.in(far_0_635_0[1]), .out(far_0_635_1[1]));
    assign layer_0[635] = ~far_0_635_1[1] | (far_0_635_1[0] & far_0_635_1[1]); 
    wire [1:0] far_0_636_0;    relay_conn far_0_636_0_a(.in(in[66]), .out(far_0_636_0[0]));    relay_conn far_0_636_0_b(.in(in[111]), .out(far_0_636_0[1]));
    assign layer_0[636] = ~far_0_636_0[0] | (far_0_636_0[0] & far_0_636_0[1]); 
    assign layer_0[637] = ~(in[79] & in[84]); 
    assign layer_0[638] = ~(in[84] | in[98]); 
    wire [1:0] far_0_639_0;    relay_conn far_0_639_0_a(.in(in[94]), .out(far_0_639_0[0]));    relay_conn far_0_639_0_b(.in(in[181]), .out(far_0_639_0[1]));
    wire [1:0] far_0_639_1;    relay_conn far_0_639_1_a(.in(far_0_639_0[0]), .out(far_0_639_1[0]));    relay_conn far_0_639_1_b(.in(far_0_639_0[1]), .out(far_0_639_1[1]));
    assign layer_0[639] = far_0_639_1[0] ^ far_0_639_1[1]; 
    wire [1:0] far_0_640_0;    relay_conn far_0_640_0_a(.in(in[18]), .out(far_0_640_0[0]));    relay_conn far_0_640_0_b(.in(in[132]), .out(far_0_640_0[1]));
    wire [1:0] far_0_640_1;    relay_conn far_0_640_1_a(.in(far_0_640_0[0]), .out(far_0_640_1[0]));    relay_conn far_0_640_1_b(.in(far_0_640_0[1]), .out(far_0_640_1[1]));
    wire [1:0] far_0_640_2;    relay_conn far_0_640_2_a(.in(far_0_640_1[0]), .out(far_0_640_2[0]));    relay_conn far_0_640_2_b(.in(far_0_640_1[1]), .out(far_0_640_2[1]));
    assign layer_0[640] = far_0_640_2[0]; 
    assign layer_0[641] = in[181]; 
    assign layer_0[642] = ~in[187]; 
    wire [1:0] far_0_643_0;    relay_conn far_0_643_0_a(.in(in[188]), .out(far_0_643_0[0]));    relay_conn far_0_643_0_b(.in(in[71]), .out(far_0_643_0[1]));
    wire [1:0] far_0_643_1;    relay_conn far_0_643_1_a(.in(far_0_643_0[0]), .out(far_0_643_1[0]));    relay_conn far_0_643_1_b(.in(far_0_643_0[1]), .out(far_0_643_1[1]));
    wire [1:0] far_0_643_2;    relay_conn far_0_643_2_a(.in(far_0_643_1[0]), .out(far_0_643_2[0]));    relay_conn far_0_643_2_b(.in(far_0_643_1[1]), .out(far_0_643_2[1]));
    assign layer_0[643] = far_0_643_2[1]; 
    wire [1:0] far_0_644_0;    relay_conn far_0_644_0_a(.in(in[157]), .out(far_0_644_0[0]));    relay_conn far_0_644_0_b(.in(in[105]), .out(far_0_644_0[1]));
    assign layer_0[644] = ~far_0_644_0[0]; 
    assign layer_0[645] = ~in[133]; 
    wire [1:0] far_0_646_0;    relay_conn far_0_646_0_a(.in(in[79]), .out(far_0_646_0[0]));    relay_conn far_0_646_0_b(.in(in[27]), .out(far_0_646_0[1]));
    assign layer_0[646] = ~(far_0_646_0[0] ^ far_0_646_0[1]); 
    assign layer_0[647] = ~(in[117] & in[111]); 
    wire [1:0] far_0_648_0;    relay_conn far_0_648_0_a(.in(in[18]), .out(far_0_648_0[0]));    relay_conn far_0_648_0_b(.in(in[113]), .out(far_0_648_0[1]));
    wire [1:0] far_0_648_1;    relay_conn far_0_648_1_a(.in(far_0_648_0[0]), .out(far_0_648_1[0]));    relay_conn far_0_648_1_b(.in(far_0_648_0[1]), .out(far_0_648_1[1]));
    assign layer_0[648] = ~far_0_648_1[0] | (far_0_648_1[0] & far_0_648_1[1]); 
    assign layer_0[649] = in[111] & in[99]; 
    assign layer_0[650] = in[234] ^ in[215]; 
    assign layer_0[651] = ~in[219]; 
    assign layer_0[652] = in[117] | in[142]; 
    wire [1:0] far_0_653_0;    relay_conn far_0_653_0_a(.in(in[60]), .out(far_0_653_0[0]));    relay_conn far_0_653_0_b(.in(in[134]), .out(far_0_653_0[1]));
    wire [1:0] far_0_653_1;    relay_conn far_0_653_1_a(.in(far_0_653_0[0]), .out(far_0_653_1[0]));    relay_conn far_0_653_1_b(.in(far_0_653_0[1]), .out(far_0_653_1[1]));
    assign layer_0[653] = ~(far_0_653_1[0] & far_0_653_1[1]); 
    wire [1:0] far_0_654_0;    relay_conn far_0_654_0_a(.in(in[13]), .out(far_0_654_0[0]));    relay_conn far_0_654_0_b(.in(in[71]), .out(far_0_654_0[1]));
    assign layer_0[654] = far_0_654_0[0] & far_0_654_0[1]; 
    assign layer_0[655] = ~in[113]; 
    wire [1:0] far_0_656_0;    relay_conn far_0_656_0_a(.in(in[95]), .out(far_0_656_0[0]));    relay_conn far_0_656_0_b(.in(in[223]), .out(far_0_656_0[1]));
    wire [1:0] far_0_656_1;    relay_conn far_0_656_1_a(.in(far_0_656_0[0]), .out(far_0_656_1[0]));    relay_conn far_0_656_1_b(.in(far_0_656_0[1]), .out(far_0_656_1[1]));
    wire [1:0] far_0_656_2;    relay_conn far_0_656_2_a(.in(far_0_656_1[0]), .out(far_0_656_2[0]));    relay_conn far_0_656_2_b(.in(far_0_656_1[1]), .out(far_0_656_2[1]));
    wire [1:0] far_0_656_3;    relay_conn far_0_656_3_a(.in(far_0_656_2[0]), .out(far_0_656_3[0]));    relay_conn far_0_656_3_b(.in(far_0_656_2[1]), .out(far_0_656_3[1]));
    assign layer_0[656] = ~(far_0_656_3[0] & far_0_656_3[1]); 
    wire [1:0] far_0_657_0;    relay_conn far_0_657_0_a(.in(in[236]), .out(far_0_657_0[0]));    relay_conn far_0_657_0_b(.in(in[151]), .out(far_0_657_0[1]));
    wire [1:0] far_0_657_1;    relay_conn far_0_657_1_a(.in(far_0_657_0[0]), .out(far_0_657_1[0]));    relay_conn far_0_657_1_b(.in(far_0_657_0[1]), .out(far_0_657_1[1]));
    assign layer_0[657] = far_0_657_1[0] | far_0_657_1[1]; 
    wire [1:0] far_0_658_0;    relay_conn far_0_658_0_a(.in(in[82]), .out(far_0_658_0[0]));    relay_conn far_0_658_0_b(.in(in[42]), .out(far_0_658_0[1]));
    assign layer_0[658] = far_0_658_0[0] & far_0_658_0[1]; 
    assign layer_0[659] = ~in[97]; 
    wire [1:0] far_0_660_0;    relay_conn far_0_660_0_a(.in(in[76]), .out(far_0_660_0[0]));    relay_conn far_0_660_0_b(.in(in[163]), .out(far_0_660_0[1]));
    wire [1:0] far_0_660_1;    relay_conn far_0_660_1_a(.in(far_0_660_0[0]), .out(far_0_660_1[0]));    relay_conn far_0_660_1_b(.in(far_0_660_0[1]), .out(far_0_660_1[1]));
    assign layer_0[660] = ~(far_0_660_1[0] & far_0_660_1[1]); 
    wire [1:0] far_0_661_0;    relay_conn far_0_661_0_a(.in(in[187]), .out(far_0_661_0[0]));    relay_conn far_0_661_0_b(.in(in[59]), .out(far_0_661_0[1]));
    wire [1:0] far_0_661_1;    relay_conn far_0_661_1_a(.in(far_0_661_0[0]), .out(far_0_661_1[0]));    relay_conn far_0_661_1_b(.in(far_0_661_0[1]), .out(far_0_661_1[1]));
    wire [1:0] far_0_661_2;    relay_conn far_0_661_2_a(.in(far_0_661_1[0]), .out(far_0_661_2[0]));    relay_conn far_0_661_2_b(.in(far_0_661_1[1]), .out(far_0_661_2[1]));
    wire [1:0] far_0_661_3;    relay_conn far_0_661_3_a(.in(far_0_661_2[0]), .out(far_0_661_3[0]));    relay_conn far_0_661_3_b(.in(far_0_661_2[1]), .out(far_0_661_3[1]));
    assign layer_0[661] = far_0_661_3[0]; 
    assign layer_0[662] = in[215] | in[186]; 
    wire [1:0] far_0_663_0;    relay_conn far_0_663_0_a(.in(in[19]), .out(far_0_663_0[0]));    relay_conn far_0_663_0_b(.in(in[72]), .out(far_0_663_0[1]));
    assign layer_0[663] = far_0_663_0[0] & far_0_663_0[1]; 
    wire [1:0] far_0_664_0;    relay_conn far_0_664_0_a(.in(in[79]), .out(far_0_664_0[0]));    relay_conn far_0_664_0_b(.in(in[151]), .out(far_0_664_0[1]));
    wire [1:0] far_0_664_1;    relay_conn far_0_664_1_a(.in(far_0_664_0[0]), .out(far_0_664_1[0]));    relay_conn far_0_664_1_b(.in(far_0_664_0[1]), .out(far_0_664_1[1]));
    assign layer_0[664] = far_0_664_1[1] & ~far_0_664_1[0]; 
    assign layer_0[665] = in[212] | in[236]; 
    assign layer_0[666] = in[229] | in[236]; 
    assign layer_0[667] = in[202] & ~in[183]; 
    wire [1:0] far_0_668_0;    relay_conn far_0_668_0_a(.in(in[149]), .out(far_0_668_0[0]));    relay_conn far_0_668_0_b(.in(in[99]), .out(far_0_668_0[1]));
    assign layer_0[668] = ~(far_0_668_0[0] | far_0_668_0[1]); 
    wire [1:0] far_0_669_0;    relay_conn far_0_669_0_a(.in(in[82]), .out(far_0_669_0[0]));    relay_conn far_0_669_0_b(.in(in[203]), .out(far_0_669_0[1]));
    wire [1:0] far_0_669_1;    relay_conn far_0_669_1_a(.in(far_0_669_0[0]), .out(far_0_669_1[0]));    relay_conn far_0_669_1_b(.in(far_0_669_0[1]), .out(far_0_669_1[1]));
    wire [1:0] far_0_669_2;    relay_conn far_0_669_2_a(.in(far_0_669_1[0]), .out(far_0_669_2[0]));    relay_conn far_0_669_2_b(.in(far_0_669_1[1]), .out(far_0_669_2[1]));
    assign layer_0[669] = ~far_0_669_2[1]; 
    assign layer_0[670] = in[121] | in[140]; 
    wire [1:0] far_0_671_0;    relay_conn far_0_671_0_a(.in(in[109]), .out(far_0_671_0[0]));    relay_conn far_0_671_0_b(.in(in[207]), .out(far_0_671_0[1]));
    wire [1:0] far_0_671_1;    relay_conn far_0_671_1_a(.in(far_0_671_0[0]), .out(far_0_671_1[0]));    relay_conn far_0_671_1_b(.in(far_0_671_0[1]), .out(far_0_671_1[1]));
    wire [1:0] far_0_671_2;    relay_conn far_0_671_2_a(.in(far_0_671_1[0]), .out(far_0_671_2[0]));    relay_conn far_0_671_2_b(.in(far_0_671_1[1]), .out(far_0_671_2[1]));
    assign layer_0[671] = ~(far_0_671_2[0] ^ far_0_671_2[1]); 
    wire [1:0] far_0_672_0;    relay_conn far_0_672_0_a(.in(in[189]), .out(far_0_672_0[0]));    relay_conn far_0_672_0_b(.in(in[113]), .out(far_0_672_0[1]));
    wire [1:0] far_0_672_1;    relay_conn far_0_672_1_a(.in(far_0_672_0[0]), .out(far_0_672_1[0]));    relay_conn far_0_672_1_b(.in(far_0_672_0[1]), .out(far_0_672_1[1]));
    assign layer_0[672] = far_0_672_1[0] & ~far_0_672_1[1]; 
    wire [1:0] far_0_673_0;    relay_conn far_0_673_0_a(.in(in[111]), .out(far_0_673_0[0]));    relay_conn far_0_673_0_b(.in(in[151]), .out(far_0_673_0[1]));
    assign layer_0[673] = ~far_0_673_0[1]; 
    wire [1:0] far_0_674_0;    relay_conn far_0_674_0_a(.in(in[22]), .out(far_0_674_0[0]));    relay_conn far_0_674_0_b(.in(in[95]), .out(far_0_674_0[1]));
    wire [1:0] far_0_674_1;    relay_conn far_0_674_1_a(.in(far_0_674_0[0]), .out(far_0_674_1[0]));    relay_conn far_0_674_1_b(.in(far_0_674_0[1]), .out(far_0_674_1[1]));
    assign layer_0[674] = far_0_674_1[0] & far_0_674_1[1]; 
    wire [1:0] far_0_675_0;    relay_conn far_0_675_0_a(.in(in[198]), .out(far_0_675_0[0]));    relay_conn far_0_675_0_b(.in(in[90]), .out(far_0_675_0[1]));
    wire [1:0] far_0_675_1;    relay_conn far_0_675_1_a(.in(far_0_675_0[0]), .out(far_0_675_1[0]));    relay_conn far_0_675_1_b(.in(far_0_675_0[1]), .out(far_0_675_1[1]));
    wire [1:0] far_0_675_2;    relay_conn far_0_675_2_a(.in(far_0_675_1[0]), .out(far_0_675_2[0]));    relay_conn far_0_675_2_b(.in(far_0_675_1[1]), .out(far_0_675_2[1]));
    assign layer_0[675] = far_0_675_2[1]; 
    wire [1:0] far_0_676_0;    relay_conn far_0_676_0_a(.in(in[133]), .out(far_0_676_0[0]));    relay_conn far_0_676_0_b(.in(in[78]), .out(far_0_676_0[1]));
    assign layer_0[676] = ~far_0_676_0[0] | (far_0_676_0[0] & far_0_676_0[1]); 
    wire [1:0] far_0_677_0;    relay_conn far_0_677_0_a(.in(in[211]), .out(far_0_677_0[0]));    relay_conn far_0_677_0_b(.in(in[159]), .out(far_0_677_0[1]));
    assign layer_0[677] = ~(far_0_677_0[0] | far_0_677_0[1]); 
    wire [1:0] far_0_678_0;    relay_conn far_0_678_0_a(.in(in[75]), .out(far_0_678_0[0]));    relay_conn far_0_678_0_b(.in(in[182]), .out(far_0_678_0[1]));
    wire [1:0] far_0_678_1;    relay_conn far_0_678_1_a(.in(far_0_678_0[0]), .out(far_0_678_1[0]));    relay_conn far_0_678_1_b(.in(far_0_678_0[1]), .out(far_0_678_1[1]));
    wire [1:0] far_0_678_2;    relay_conn far_0_678_2_a(.in(far_0_678_1[0]), .out(far_0_678_2[0]));    relay_conn far_0_678_2_b(.in(far_0_678_1[1]), .out(far_0_678_2[1]));
    assign layer_0[678] = far_0_678_2[1] & ~far_0_678_2[0]; 
    assign layer_0[679] = in[118] & ~in[127]; 
    assign layer_0[680] = in[8] & in[3]; 
    wire [1:0] far_0_681_0;    relay_conn far_0_681_0_a(.in(in[110]), .out(far_0_681_0[0]));    relay_conn far_0_681_0_b(.in(in[157]), .out(far_0_681_0[1]));
    assign layer_0[681] = ~far_0_681_0[1]; 
    assign layer_0[682] = in[17] & in[5]; 
    assign layer_0[683] = in[109] ^ in[104]; 
    assign layer_0[684] = in[75] | in[93]; 
    assign layer_0[685] = in[138] & ~in[122]; 
    wire [1:0] far_0_686_0;    relay_conn far_0_686_0_a(.in(in[151]), .out(far_0_686_0[0]));    relay_conn far_0_686_0_b(.in(in[207]), .out(far_0_686_0[1]));
    assign layer_0[686] = ~(far_0_686_0[0] & far_0_686_0[1]); 
    wire [1:0] far_0_687_0;    relay_conn far_0_687_0_a(.in(in[73]), .out(far_0_687_0[0]));    relay_conn far_0_687_0_b(.in(in[130]), .out(far_0_687_0[1]));
    assign layer_0[687] = far_0_687_0[0]; 
    assign layer_0[688] = ~in[117]; 
    wire [1:0] far_0_689_0;    relay_conn far_0_689_0_a(.in(in[73]), .out(far_0_689_0[0]));    relay_conn far_0_689_0_b(.in(in[195]), .out(far_0_689_0[1]));
    wire [1:0] far_0_689_1;    relay_conn far_0_689_1_a(.in(far_0_689_0[0]), .out(far_0_689_1[0]));    relay_conn far_0_689_1_b(.in(far_0_689_0[1]), .out(far_0_689_1[1]));
    wire [1:0] far_0_689_2;    relay_conn far_0_689_2_a(.in(far_0_689_1[0]), .out(far_0_689_2[0]));    relay_conn far_0_689_2_b(.in(far_0_689_1[1]), .out(far_0_689_2[1]));
    assign layer_0[689] = far_0_689_2[0] | far_0_689_2[1]; 
    wire [1:0] far_0_690_0;    relay_conn far_0_690_0_a(.in(in[221]), .out(far_0_690_0[0]));    relay_conn far_0_690_0_b(.in(in[150]), .out(far_0_690_0[1]));
    wire [1:0] far_0_690_1;    relay_conn far_0_690_1_a(.in(far_0_690_0[0]), .out(far_0_690_1[0]));    relay_conn far_0_690_1_b(.in(far_0_690_0[1]), .out(far_0_690_1[1]));
    assign layer_0[690] = ~(far_0_690_1[0] & far_0_690_1[1]); 
    assign layer_0[691] = in[172]; 
    wire [1:0] far_0_692_0;    relay_conn far_0_692_0_a(.in(in[117]), .out(far_0_692_0[0]));    relay_conn far_0_692_0_b(.in(in[151]), .out(far_0_692_0[1]));
    assign layer_0[692] = ~far_0_692_0[0]; 
    wire [1:0] far_0_693_0;    relay_conn far_0_693_0_a(.in(in[197]), .out(far_0_693_0[0]));    relay_conn far_0_693_0_b(.in(in[109]), .out(far_0_693_0[1]));
    wire [1:0] far_0_693_1;    relay_conn far_0_693_1_a(.in(far_0_693_0[0]), .out(far_0_693_1[0]));    relay_conn far_0_693_1_b(.in(far_0_693_0[1]), .out(far_0_693_1[1]));
    assign layer_0[693] = ~far_0_693_1[0] | (far_0_693_1[0] & far_0_693_1[1]); 
    assign layer_0[694] = ~in[221]; 
    wire [1:0] far_0_695_0;    relay_conn far_0_695_0_a(.in(in[133]), .out(far_0_695_0[0]));    relay_conn far_0_695_0_b(.in(in[11]), .out(far_0_695_0[1]));
    wire [1:0] far_0_695_1;    relay_conn far_0_695_1_a(.in(far_0_695_0[0]), .out(far_0_695_1[0]));    relay_conn far_0_695_1_b(.in(far_0_695_0[1]), .out(far_0_695_1[1]));
    wire [1:0] far_0_695_2;    relay_conn far_0_695_2_a(.in(far_0_695_1[0]), .out(far_0_695_2[0]));    relay_conn far_0_695_2_b(.in(far_0_695_1[1]), .out(far_0_695_2[1]));
    assign layer_0[695] = far_0_695_2[1] & ~far_0_695_2[0]; 
    assign layer_0[696] = in[57] | in[63]; 
    wire [1:0] far_0_697_0;    relay_conn far_0_697_0_a(.in(in[202]), .out(far_0_697_0[0]));    relay_conn far_0_697_0_b(.in(in[89]), .out(far_0_697_0[1]));
    wire [1:0] far_0_697_1;    relay_conn far_0_697_1_a(.in(far_0_697_0[0]), .out(far_0_697_1[0]));    relay_conn far_0_697_1_b(.in(far_0_697_0[1]), .out(far_0_697_1[1]));
    wire [1:0] far_0_697_2;    relay_conn far_0_697_2_a(.in(far_0_697_1[0]), .out(far_0_697_2[0]));    relay_conn far_0_697_2_b(.in(far_0_697_1[1]), .out(far_0_697_2[1]));
    assign layer_0[697] = ~far_0_697_2[1]; 
    assign layer_0[698] = ~(in[43] | in[34]); 
    assign layer_0[699] = in[4] & ~in[25]; 
    wire [1:0] far_0_700_0;    relay_conn far_0_700_0_a(.in(in[157]), .out(far_0_700_0[0]));    relay_conn far_0_700_0_b(.in(in[250]), .out(far_0_700_0[1]));
    wire [1:0] far_0_700_1;    relay_conn far_0_700_1_a(.in(far_0_700_0[0]), .out(far_0_700_1[0]));    relay_conn far_0_700_1_b(.in(far_0_700_0[1]), .out(far_0_700_1[1]));
    assign layer_0[700] = far_0_700_1[0]; 
    wire [1:0] far_0_701_0;    relay_conn far_0_701_0_a(.in(in[39]), .out(far_0_701_0[0]));    relay_conn far_0_701_0_b(.in(in[104]), .out(far_0_701_0[1]));
    wire [1:0] far_0_701_1;    relay_conn far_0_701_1_a(.in(far_0_701_0[0]), .out(far_0_701_1[0]));    relay_conn far_0_701_1_b(.in(far_0_701_0[1]), .out(far_0_701_1[1]));
    assign layer_0[701] = far_0_701_1[0] | far_0_701_1[1]; 
    wire [1:0] far_0_702_0;    relay_conn far_0_702_0_a(.in(in[136]), .out(far_0_702_0[0]));    relay_conn far_0_702_0_b(.in(in[66]), .out(far_0_702_0[1]));
    wire [1:0] far_0_702_1;    relay_conn far_0_702_1_a(.in(far_0_702_0[0]), .out(far_0_702_1[0]));    relay_conn far_0_702_1_b(.in(far_0_702_0[1]), .out(far_0_702_1[1]));
    assign layer_0[702] = far_0_702_1[0]; 
    wire [1:0] far_0_703_0;    relay_conn far_0_703_0_a(.in(in[121]), .out(far_0_703_0[0]));    relay_conn far_0_703_0_b(.in(in[193]), .out(far_0_703_0[1]));
    wire [1:0] far_0_703_1;    relay_conn far_0_703_1_a(.in(far_0_703_0[0]), .out(far_0_703_1[0]));    relay_conn far_0_703_1_b(.in(far_0_703_0[1]), .out(far_0_703_1[1]));
    assign layer_0[703] = far_0_703_1[0] | far_0_703_1[1]; 
    wire [1:0] far_0_704_0;    relay_conn far_0_704_0_a(.in(in[59]), .out(far_0_704_0[0]));    relay_conn far_0_704_0_b(.in(in[100]), .out(far_0_704_0[1]));
    assign layer_0[704] = ~far_0_704_0[1] | (far_0_704_0[0] & far_0_704_0[1]); 
    assign layer_0[705] = ~in[187]; 
    assign layer_0[706] = in[5] & in[36]; 
    wire [1:0] far_0_707_0;    relay_conn far_0_707_0_a(.in(in[84]), .out(far_0_707_0[0]));    relay_conn far_0_707_0_b(.in(in[212]), .out(far_0_707_0[1]));
    wire [1:0] far_0_707_1;    relay_conn far_0_707_1_a(.in(far_0_707_0[0]), .out(far_0_707_1[0]));    relay_conn far_0_707_1_b(.in(far_0_707_0[1]), .out(far_0_707_1[1]));
    wire [1:0] far_0_707_2;    relay_conn far_0_707_2_a(.in(far_0_707_1[0]), .out(far_0_707_2[0]));    relay_conn far_0_707_2_b(.in(far_0_707_1[1]), .out(far_0_707_2[1]));
    wire [1:0] far_0_707_3;    relay_conn far_0_707_3_a(.in(far_0_707_2[0]), .out(far_0_707_3[0]));    relay_conn far_0_707_3_b(.in(far_0_707_2[1]), .out(far_0_707_3[1]));
    assign layer_0[707] = far_0_707_3[0] & far_0_707_3[1]; 
    assign layer_0[708] = in[67] & ~in[84]; 
    assign layer_0[709] = ~in[132] | (in[132] & in[133]); 
    wire [1:0] far_0_710_0;    relay_conn far_0_710_0_a(.in(in[197]), .out(far_0_710_0[0]));    relay_conn far_0_710_0_b(.in(in[136]), .out(far_0_710_0[1]));
    assign layer_0[710] = ~far_0_710_0[0] | (far_0_710_0[0] & far_0_710_0[1]); 
    wire [1:0] far_0_711_0;    relay_conn far_0_711_0_a(.in(in[13]), .out(far_0_711_0[0]));    relay_conn far_0_711_0_b(.in(in[107]), .out(far_0_711_0[1]));
    wire [1:0] far_0_711_1;    relay_conn far_0_711_1_a(.in(far_0_711_0[0]), .out(far_0_711_1[0]));    relay_conn far_0_711_1_b(.in(far_0_711_0[1]), .out(far_0_711_1[1]));
    assign layer_0[711] = far_0_711_1[1]; 
    assign layer_0[712] = in[113] & ~in[105]; 
    wire [1:0] far_0_713_0;    relay_conn far_0_713_0_a(.in(in[128]), .out(far_0_713_0[0]));    relay_conn far_0_713_0_b(.in(in[164]), .out(far_0_713_0[1]));
    assign layer_0[713] = ~far_0_713_0[1]; 
    wire [1:0] far_0_714_0;    relay_conn far_0_714_0_a(.in(in[63]), .out(far_0_714_0[0]));    relay_conn far_0_714_0_b(.in(in[187]), .out(far_0_714_0[1]));
    wire [1:0] far_0_714_1;    relay_conn far_0_714_1_a(.in(far_0_714_0[0]), .out(far_0_714_1[0]));    relay_conn far_0_714_1_b(.in(far_0_714_0[1]), .out(far_0_714_1[1]));
    wire [1:0] far_0_714_2;    relay_conn far_0_714_2_a(.in(far_0_714_1[0]), .out(far_0_714_2[0]));    relay_conn far_0_714_2_b(.in(far_0_714_1[1]), .out(far_0_714_2[1]));
    assign layer_0[714] = far_0_714_2[0] ^ far_0_714_2[1]; 
    wire [1:0] far_0_715_0;    relay_conn far_0_715_0_a(.in(in[94]), .out(far_0_715_0[0]));    relay_conn far_0_715_0_b(.in(in[171]), .out(far_0_715_0[1]));
    wire [1:0] far_0_715_1;    relay_conn far_0_715_1_a(.in(far_0_715_0[0]), .out(far_0_715_1[0]));    relay_conn far_0_715_1_b(.in(far_0_715_0[1]), .out(far_0_715_1[1]));
    assign layer_0[715] = far_0_715_1[0] & ~far_0_715_1[1]; 
    wire [1:0] far_0_716_0;    relay_conn far_0_716_0_a(.in(in[113]), .out(far_0_716_0[0]));    relay_conn far_0_716_0_b(.in(in[216]), .out(far_0_716_0[1]));
    wire [1:0] far_0_716_1;    relay_conn far_0_716_1_a(.in(far_0_716_0[0]), .out(far_0_716_1[0]));    relay_conn far_0_716_1_b(.in(far_0_716_0[1]), .out(far_0_716_1[1]));
    wire [1:0] far_0_716_2;    relay_conn far_0_716_2_a(.in(far_0_716_1[0]), .out(far_0_716_2[0]));    relay_conn far_0_716_2_b(.in(far_0_716_1[1]), .out(far_0_716_2[1]));
    assign layer_0[716] = ~far_0_716_2[1]; 
    wire [1:0] far_0_717_0;    relay_conn far_0_717_0_a(.in(in[83]), .out(far_0_717_0[0]));    relay_conn far_0_717_0_b(.in(in[133]), .out(far_0_717_0[1]));
    assign layer_0[717] = ~(far_0_717_0[0] ^ far_0_717_0[1]); 
    wire [1:0] far_0_718_0;    relay_conn far_0_718_0_a(.in(in[53]), .out(far_0_718_0[0]));    relay_conn far_0_718_0_b(.in(in[164]), .out(far_0_718_0[1]));
    wire [1:0] far_0_718_1;    relay_conn far_0_718_1_a(.in(far_0_718_0[0]), .out(far_0_718_1[0]));    relay_conn far_0_718_1_b(.in(far_0_718_0[1]), .out(far_0_718_1[1]));
    wire [1:0] far_0_718_2;    relay_conn far_0_718_2_a(.in(far_0_718_1[0]), .out(far_0_718_2[0]));    relay_conn far_0_718_2_b(.in(far_0_718_1[1]), .out(far_0_718_2[1]));
    assign layer_0[718] = far_0_718_2[0] ^ far_0_718_2[1]; 
    wire [1:0] far_0_719_0;    relay_conn far_0_719_0_a(.in(in[199]), .out(far_0_719_0[0]));    relay_conn far_0_719_0_b(.in(in[91]), .out(far_0_719_0[1]));
    wire [1:0] far_0_719_1;    relay_conn far_0_719_1_a(.in(far_0_719_0[0]), .out(far_0_719_1[0]));    relay_conn far_0_719_1_b(.in(far_0_719_0[1]), .out(far_0_719_1[1]));
    wire [1:0] far_0_719_2;    relay_conn far_0_719_2_a(.in(far_0_719_1[0]), .out(far_0_719_2[0]));    relay_conn far_0_719_2_b(.in(far_0_719_1[1]), .out(far_0_719_2[1]));
    assign layer_0[719] = far_0_719_2[1] & ~far_0_719_2[0]; 
    wire [1:0] far_0_720_0;    relay_conn far_0_720_0_a(.in(in[186]), .out(far_0_720_0[0]));    relay_conn far_0_720_0_b(.in(in[134]), .out(far_0_720_0[1]));
    assign layer_0[720] = far_0_720_0[0] & far_0_720_0[1]; 
    assign layer_0[721] = ~in[37]; 
    wire [1:0] far_0_722_0;    relay_conn far_0_722_0_a(.in(in[65]), .out(far_0_722_0[0]));    relay_conn far_0_722_0_b(.in(in[13]), .out(far_0_722_0[1]));
    assign layer_0[722] = far_0_722_0[0] | far_0_722_0[1]; 
    assign layer_0[723] = in[116]; 
    assign layer_0[724] = ~in[191] | (in[191] & in[167]); 
    assign layer_0[725] = ~(in[190] | in[213]); 
    wire [1:0] far_0_726_0;    relay_conn far_0_726_0_a(.in(in[117]), .out(far_0_726_0[0]));    relay_conn far_0_726_0_b(.in(in[230]), .out(far_0_726_0[1]));
    wire [1:0] far_0_726_1;    relay_conn far_0_726_1_a(.in(far_0_726_0[0]), .out(far_0_726_1[0]));    relay_conn far_0_726_1_b(.in(far_0_726_0[1]), .out(far_0_726_1[1]));
    wire [1:0] far_0_726_2;    relay_conn far_0_726_2_a(.in(far_0_726_1[0]), .out(far_0_726_2[0]));    relay_conn far_0_726_2_b(.in(far_0_726_1[1]), .out(far_0_726_2[1]));
    assign layer_0[726] = ~far_0_726_2[1] | (far_0_726_2[0] & far_0_726_2[1]); 
    wire [1:0] far_0_727_0;    relay_conn far_0_727_0_a(.in(in[172]), .out(far_0_727_0[0]));    relay_conn far_0_727_0_b(.in(in[82]), .out(far_0_727_0[1]));
    wire [1:0] far_0_727_1;    relay_conn far_0_727_1_a(.in(far_0_727_0[0]), .out(far_0_727_1[0]));    relay_conn far_0_727_1_b(.in(far_0_727_0[1]), .out(far_0_727_1[1]));
    assign layer_0[727] = far_0_727_1[0]; 
    assign layer_0[728] = in[117]; 
    wire [1:0] far_0_729_0;    relay_conn far_0_729_0_a(.in(in[22]), .out(far_0_729_0[0]));    relay_conn far_0_729_0_b(.in(in[109]), .out(far_0_729_0[1]));
    wire [1:0] far_0_729_1;    relay_conn far_0_729_1_a(.in(far_0_729_0[0]), .out(far_0_729_1[0]));    relay_conn far_0_729_1_b(.in(far_0_729_0[1]), .out(far_0_729_1[1]));
    assign layer_0[729] = ~(far_0_729_1[0] | far_0_729_1[1]); 
    wire [1:0] far_0_730_0;    relay_conn far_0_730_0_a(.in(in[52]), .out(far_0_730_0[0]));    relay_conn far_0_730_0_b(.in(in[156]), .out(far_0_730_0[1]));
    wire [1:0] far_0_730_1;    relay_conn far_0_730_1_a(.in(far_0_730_0[0]), .out(far_0_730_1[0]));    relay_conn far_0_730_1_b(.in(far_0_730_0[1]), .out(far_0_730_1[1]));
    wire [1:0] far_0_730_2;    relay_conn far_0_730_2_a(.in(far_0_730_1[0]), .out(far_0_730_2[0]));    relay_conn far_0_730_2_b(.in(far_0_730_1[1]), .out(far_0_730_2[1]));
    assign layer_0[730] = ~far_0_730_2[0]; 
    assign layer_0[731] = in[152]; 
    wire [1:0] far_0_732_0;    relay_conn far_0_732_0_a(.in(in[121]), .out(far_0_732_0[0]));    relay_conn far_0_732_0_b(.in(in[165]), .out(far_0_732_0[1]));
    assign layer_0[732] = ~far_0_732_0[0] | (far_0_732_0[0] & far_0_732_0[1]); 
    wire [1:0] far_0_733_0;    relay_conn far_0_733_0_a(.in(in[99]), .out(far_0_733_0[0]));    relay_conn far_0_733_0_b(.in(in[48]), .out(far_0_733_0[1]));
    assign layer_0[733] = ~far_0_733_0[0] | (far_0_733_0[0] & far_0_733_0[1]); 
    wire [1:0] far_0_734_0;    relay_conn far_0_734_0_a(.in(in[57]), .out(far_0_734_0[0]));    relay_conn far_0_734_0_b(.in(in[15]), .out(far_0_734_0[1]));
    assign layer_0[734] = far_0_734_0[0]; 
    wire [1:0] far_0_735_0;    relay_conn far_0_735_0_a(.in(in[41]), .out(far_0_735_0[0]));    relay_conn far_0_735_0_b(.in(in[158]), .out(far_0_735_0[1]));
    wire [1:0] far_0_735_1;    relay_conn far_0_735_1_a(.in(far_0_735_0[0]), .out(far_0_735_1[0]));    relay_conn far_0_735_1_b(.in(far_0_735_0[1]), .out(far_0_735_1[1]));
    wire [1:0] far_0_735_2;    relay_conn far_0_735_2_a(.in(far_0_735_1[0]), .out(far_0_735_2[0]));    relay_conn far_0_735_2_b(.in(far_0_735_1[1]), .out(far_0_735_2[1]));
    assign layer_0[735] = far_0_735_2[1]; 
    assign layer_0[736] = in[232] & ~in[202]; 
    wire [1:0] far_0_737_0;    relay_conn far_0_737_0_a(.in(in[113]), .out(far_0_737_0[0]));    relay_conn far_0_737_0_b(.in(in[16]), .out(far_0_737_0[1]));
    wire [1:0] far_0_737_1;    relay_conn far_0_737_1_a(.in(far_0_737_0[0]), .out(far_0_737_1[0]));    relay_conn far_0_737_1_b(.in(far_0_737_0[1]), .out(far_0_737_1[1]));
    wire [1:0] far_0_737_2;    relay_conn far_0_737_2_a(.in(far_0_737_1[0]), .out(far_0_737_2[0]));    relay_conn far_0_737_2_b(.in(far_0_737_1[1]), .out(far_0_737_2[1]));
    assign layer_0[737] = far_0_737_2[0] & ~far_0_737_2[1]; 
    wire [1:0] far_0_738_0;    relay_conn far_0_738_0_a(.in(in[119]), .out(far_0_738_0[0]));    relay_conn far_0_738_0_b(.in(in[213]), .out(far_0_738_0[1]));
    wire [1:0] far_0_738_1;    relay_conn far_0_738_1_a(.in(far_0_738_0[0]), .out(far_0_738_1[0]));    relay_conn far_0_738_1_b(.in(far_0_738_0[1]), .out(far_0_738_1[1]));
    assign layer_0[738] = far_0_738_1[0] | far_0_738_1[1]; 
    wire [1:0] far_0_739_0;    relay_conn far_0_739_0_a(.in(in[109]), .out(far_0_739_0[0]));    relay_conn far_0_739_0_b(.in(in[215]), .out(far_0_739_0[1]));
    wire [1:0] far_0_739_1;    relay_conn far_0_739_1_a(.in(far_0_739_0[0]), .out(far_0_739_1[0]));    relay_conn far_0_739_1_b(.in(far_0_739_0[1]), .out(far_0_739_1[1]));
    wire [1:0] far_0_739_2;    relay_conn far_0_739_2_a(.in(far_0_739_1[0]), .out(far_0_739_2[0]));    relay_conn far_0_739_2_b(.in(far_0_739_1[1]), .out(far_0_739_2[1]));
    assign layer_0[739] = ~(far_0_739_2[0] ^ far_0_739_2[1]); 
    wire [1:0] far_0_740_0;    relay_conn far_0_740_0_a(.in(in[195]), .out(far_0_740_0[0]));    relay_conn far_0_740_0_b(.in(in[149]), .out(far_0_740_0[1]));
    assign layer_0[740] = far_0_740_0[0] & ~far_0_740_0[1]; 
    wire [1:0] far_0_741_0;    relay_conn far_0_741_0_a(.in(in[74]), .out(far_0_741_0[0]));    relay_conn far_0_741_0_b(.in(in[151]), .out(far_0_741_0[1]));
    wire [1:0] far_0_741_1;    relay_conn far_0_741_1_a(.in(far_0_741_0[0]), .out(far_0_741_1[0]));    relay_conn far_0_741_1_b(.in(far_0_741_0[1]), .out(far_0_741_1[1]));
    assign layer_0[741] = ~(far_0_741_1[0] | far_0_741_1[1]); 
    wire [1:0] far_0_742_0;    relay_conn far_0_742_0_a(.in(in[79]), .out(far_0_742_0[0]));    relay_conn far_0_742_0_b(.in(in[113]), .out(far_0_742_0[1]));
    assign layer_0[742] = far_0_742_0[0] & ~far_0_742_0[1]; 
    wire [1:0] far_0_743_0;    relay_conn far_0_743_0_a(.in(in[10]), .out(far_0_743_0[0]));    relay_conn far_0_743_0_b(.in(in[87]), .out(far_0_743_0[1]));
    wire [1:0] far_0_743_1;    relay_conn far_0_743_1_a(.in(far_0_743_0[0]), .out(far_0_743_1[0]));    relay_conn far_0_743_1_b(.in(far_0_743_0[1]), .out(far_0_743_1[1]));
    assign layer_0[743] = far_0_743_1[0] & ~far_0_743_1[1]; 
    assign layer_0[744] = ~in[109]; 
    wire [1:0] far_0_745_0;    relay_conn far_0_745_0_a(.in(in[99]), .out(far_0_745_0[0]));    relay_conn far_0_745_0_b(.in(in[221]), .out(far_0_745_0[1]));
    wire [1:0] far_0_745_1;    relay_conn far_0_745_1_a(.in(far_0_745_0[0]), .out(far_0_745_1[0]));    relay_conn far_0_745_1_b(.in(far_0_745_0[1]), .out(far_0_745_1[1]));
    wire [1:0] far_0_745_2;    relay_conn far_0_745_2_a(.in(far_0_745_1[0]), .out(far_0_745_2[0]));    relay_conn far_0_745_2_b(.in(far_0_745_1[1]), .out(far_0_745_2[1]));
    assign layer_0[745] = far_0_745_2[0]; 
    wire [1:0] far_0_746_0;    relay_conn far_0_746_0_a(.in(in[46]), .out(far_0_746_0[0]));    relay_conn far_0_746_0_b(.in(in[134]), .out(far_0_746_0[1]));
    wire [1:0] far_0_746_1;    relay_conn far_0_746_1_a(.in(far_0_746_0[0]), .out(far_0_746_1[0]));    relay_conn far_0_746_1_b(.in(far_0_746_0[1]), .out(far_0_746_1[1]));
    assign layer_0[746] = ~(far_0_746_1[0] | far_0_746_1[1]); 
    wire [1:0] far_0_747_0;    relay_conn far_0_747_0_a(.in(in[239]), .out(far_0_747_0[0]));    relay_conn far_0_747_0_b(.in(in[197]), .out(far_0_747_0[1]));
    assign layer_0[747] = far_0_747_0[1] & ~far_0_747_0[0]; 
    assign layer_0[748] = in[203] & ~in[187]; 
    wire [1:0] far_0_749_0;    relay_conn far_0_749_0_a(.in(in[199]), .out(far_0_749_0[0]));    relay_conn far_0_749_0_b(.in(in[236]), .out(far_0_749_0[1]));
    assign layer_0[749] = ~far_0_749_0[0] | (far_0_749_0[0] & far_0_749_0[1]); 
    wire [1:0] far_0_750_0;    relay_conn far_0_750_0_a(.in(in[132]), .out(far_0_750_0[0]));    relay_conn far_0_750_0_b(.in(in[215]), .out(far_0_750_0[1]));
    wire [1:0] far_0_750_1;    relay_conn far_0_750_1_a(.in(far_0_750_0[0]), .out(far_0_750_1[0]));    relay_conn far_0_750_1_b(.in(far_0_750_0[1]), .out(far_0_750_1[1]));
    assign layer_0[750] = ~far_0_750_1[1] | (far_0_750_1[0] & far_0_750_1[1]); 
    wire [1:0] far_0_751_0;    relay_conn far_0_751_0_a(.in(in[151]), .out(far_0_751_0[0]));    relay_conn far_0_751_0_b(.in(in[74]), .out(far_0_751_0[1]));
    wire [1:0] far_0_751_1;    relay_conn far_0_751_1_a(.in(far_0_751_0[0]), .out(far_0_751_1[0]));    relay_conn far_0_751_1_b(.in(far_0_751_0[1]), .out(far_0_751_1[1]));
    assign layer_0[751] = far_0_751_1[0] & ~far_0_751_1[1]; 
    assign layer_0[752] = in[241] & ~in[211]; 
    wire [1:0] far_0_753_0;    relay_conn far_0_753_0_a(.in(in[55]), .out(far_0_753_0[0]));    relay_conn far_0_753_0_b(.in(in[87]), .out(far_0_753_0[1]));
    assign layer_0[753] = far_0_753_0[0] | far_0_753_0[1]; 
    assign layer_0[754] = ~in[34] | (in[34] & in[57]); 
    wire [1:0] far_0_755_0;    relay_conn far_0_755_0_a(.in(in[51]), .out(far_0_755_0[0]));    relay_conn far_0_755_0_b(.in(in[94]), .out(far_0_755_0[1]));
    assign layer_0[755] = far_0_755_0[0] | far_0_755_0[1]; 
    wire [1:0] far_0_756_0;    relay_conn far_0_756_0_a(.in(in[229]), .out(far_0_756_0[0]));    relay_conn far_0_756_0_b(.in(in[170]), .out(far_0_756_0[1]));
    assign layer_0[756] = far_0_756_0[0] ^ far_0_756_0[1]; 
    wire [1:0] far_0_757_0;    relay_conn far_0_757_0_a(.in(in[215]), .out(far_0_757_0[0]));    relay_conn far_0_757_0_b(.in(in[157]), .out(far_0_757_0[1]));
    assign layer_0[757] = ~far_0_757_0[1]; 
    assign layer_0[758] = in[113]; 
    assign layer_0[759] = in[212] & in[207]; 
    assign layer_0[760] = in[113] & ~in[125]; 
    wire [1:0] far_0_761_0;    relay_conn far_0_761_0_a(.in(in[157]), .out(far_0_761_0[0]));    relay_conn far_0_761_0_b(.in(in[202]), .out(far_0_761_0[1]));
    assign layer_0[761] = ~far_0_761_0[0] | (far_0_761_0[0] & far_0_761_0[1]); 
    wire [1:0] far_0_762_0;    relay_conn far_0_762_0_a(.in(in[3]), .out(far_0_762_0[0]));    relay_conn far_0_762_0_b(.in(in[113]), .out(far_0_762_0[1]));
    wire [1:0] far_0_762_1;    relay_conn far_0_762_1_a(.in(far_0_762_0[0]), .out(far_0_762_1[0]));    relay_conn far_0_762_1_b(.in(far_0_762_0[1]), .out(far_0_762_1[1]));
    wire [1:0] far_0_762_2;    relay_conn far_0_762_2_a(.in(far_0_762_1[0]), .out(far_0_762_2[0]));    relay_conn far_0_762_2_b(.in(far_0_762_1[1]), .out(far_0_762_2[1]));
    assign layer_0[762] = far_0_762_2[1] & ~far_0_762_2[0]; 
    wire [1:0] far_0_763_0;    relay_conn far_0_763_0_a(.in(in[121]), .out(far_0_763_0[0]));    relay_conn far_0_763_0_b(.in(in[187]), .out(far_0_763_0[1]));
    wire [1:0] far_0_763_1;    relay_conn far_0_763_1_a(.in(far_0_763_0[0]), .out(far_0_763_1[0]));    relay_conn far_0_763_1_b(.in(far_0_763_0[1]), .out(far_0_763_1[1]));
    assign layer_0[763] = ~far_0_763_1[0] | (far_0_763_1[0] & far_0_763_1[1]); 
    wire [1:0] far_0_764_0;    relay_conn far_0_764_0_a(.in(in[207]), .out(far_0_764_0[0]));    relay_conn far_0_764_0_b(.in(in[99]), .out(far_0_764_0[1]));
    wire [1:0] far_0_764_1;    relay_conn far_0_764_1_a(.in(far_0_764_0[0]), .out(far_0_764_1[0]));    relay_conn far_0_764_1_b(.in(far_0_764_0[1]), .out(far_0_764_1[1]));
    wire [1:0] far_0_764_2;    relay_conn far_0_764_2_a(.in(far_0_764_1[0]), .out(far_0_764_2[0]));    relay_conn far_0_764_2_b(.in(far_0_764_1[1]), .out(far_0_764_2[1]));
    assign layer_0[764] = ~(far_0_764_2[0] & far_0_764_2[1]); 
    wire [1:0] far_0_765_0;    relay_conn far_0_765_0_a(.in(in[51]), .out(far_0_765_0[0]));    relay_conn far_0_765_0_b(.in(in[161]), .out(far_0_765_0[1]));
    wire [1:0] far_0_765_1;    relay_conn far_0_765_1_a(.in(far_0_765_0[0]), .out(far_0_765_1[0]));    relay_conn far_0_765_1_b(.in(far_0_765_0[1]), .out(far_0_765_1[1]));
    wire [1:0] far_0_765_2;    relay_conn far_0_765_2_a(.in(far_0_765_1[0]), .out(far_0_765_2[0]));    relay_conn far_0_765_2_b(.in(far_0_765_1[1]), .out(far_0_765_2[1]));
    assign layer_0[765] = far_0_765_2[1] & ~far_0_765_2[0]; 
    wire [1:0] far_0_766_0;    relay_conn far_0_766_0_a(.in(in[52]), .out(far_0_766_0[0]));    relay_conn far_0_766_0_b(.in(in[107]), .out(far_0_766_0[1]));
    assign layer_0[766] = far_0_766_0[0] & ~far_0_766_0[1]; 
    wire [1:0] far_0_767_0;    relay_conn far_0_767_0_a(.in(in[165]), .out(far_0_767_0[0]));    relay_conn far_0_767_0_b(.in(in[215]), .out(far_0_767_0[1]));
    assign layer_0[767] = far_0_767_0[0] & ~far_0_767_0[1]; 
    wire [1:0] far_0_768_0;    relay_conn far_0_768_0_a(.in(in[10]), .out(far_0_768_0[0]));    relay_conn far_0_768_0_b(.in(in[84]), .out(far_0_768_0[1]));
    wire [1:0] far_0_768_1;    relay_conn far_0_768_1_a(.in(far_0_768_0[0]), .out(far_0_768_1[0]));    relay_conn far_0_768_1_b(.in(far_0_768_0[1]), .out(far_0_768_1[1]));
    assign layer_0[768] = ~far_0_768_1[0] | (far_0_768_1[0] & far_0_768_1[1]); 
    wire [1:0] far_0_769_0;    relay_conn far_0_769_0_a(.in(in[117]), .out(far_0_769_0[0]));    relay_conn far_0_769_0_b(.in(in[151]), .out(far_0_769_0[1]));
    assign layer_0[769] = far_0_769_0[0]; 
    wire [1:0] far_0_770_0;    relay_conn far_0_770_0_a(.in(in[36]), .out(far_0_770_0[0]));    relay_conn far_0_770_0_b(.in(in[157]), .out(far_0_770_0[1]));
    wire [1:0] far_0_770_1;    relay_conn far_0_770_1_a(.in(far_0_770_0[0]), .out(far_0_770_1[0]));    relay_conn far_0_770_1_b(.in(far_0_770_0[1]), .out(far_0_770_1[1]));
    wire [1:0] far_0_770_2;    relay_conn far_0_770_2_a(.in(far_0_770_1[0]), .out(far_0_770_2[0]));    relay_conn far_0_770_2_b(.in(far_0_770_1[1]), .out(far_0_770_2[1]));
    assign layer_0[770] = ~far_0_770_2[0] | (far_0_770_2[0] & far_0_770_2[1]); 
    assign layer_0[771] = ~(in[80] & in[72]); 
    wire [1:0] far_0_772_0;    relay_conn far_0_772_0_a(.in(in[93]), .out(far_0_772_0[0]));    relay_conn far_0_772_0_b(.in(in[153]), .out(far_0_772_0[1]));
    assign layer_0[772] = far_0_772_0[1]; 
    wire [1:0] far_0_773_0;    relay_conn far_0_773_0_a(.in(in[207]), .out(far_0_773_0[0]));    relay_conn far_0_773_0_b(.in(in[248]), .out(far_0_773_0[1]));
    assign layer_0[773] = far_0_773_0[1]; 
    assign layer_0[774] = in[121]; 
    assign layer_0[775] = in[181]; 
    wire [1:0] far_0_776_0;    relay_conn far_0_776_0_a(.in(in[134]), .out(far_0_776_0[0]));    relay_conn far_0_776_0_b(.in(in[37]), .out(far_0_776_0[1]));
    wire [1:0] far_0_776_1;    relay_conn far_0_776_1_a(.in(far_0_776_0[0]), .out(far_0_776_1[0]));    relay_conn far_0_776_1_b(.in(far_0_776_0[1]), .out(far_0_776_1[1]));
    wire [1:0] far_0_776_2;    relay_conn far_0_776_2_a(.in(far_0_776_1[0]), .out(far_0_776_2[0]));    relay_conn far_0_776_2_b(.in(far_0_776_1[1]), .out(far_0_776_2[1]));
    assign layer_0[776] = ~far_0_776_2[0] | (far_0_776_2[0] & far_0_776_2[1]); 
    wire [1:0] far_0_777_0;    relay_conn far_0_777_0_a(.in(in[77]), .out(far_0_777_0[0]));    relay_conn far_0_777_0_b(.in(in[30]), .out(far_0_777_0[1]));
    assign layer_0[777] = far_0_777_0[1]; 
    wire [1:0] far_0_778_0;    relay_conn far_0_778_0_a(.in(in[202]), .out(far_0_778_0[0]));    relay_conn far_0_778_0_b(.in(in[109]), .out(far_0_778_0[1]));
    wire [1:0] far_0_778_1;    relay_conn far_0_778_1_a(.in(far_0_778_0[0]), .out(far_0_778_1[0]));    relay_conn far_0_778_1_b(.in(far_0_778_0[1]), .out(far_0_778_1[1]));
    assign layer_0[778] = ~far_0_778_1[0]; 
    wire [1:0] far_0_779_0;    relay_conn far_0_779_0_a(.in(in[57]), .out(far_0_779_0[0]));    relay_conn far_0_779_0_b(.in(in[150]), .out(far_0_779_0[1]));
    wire [1:0] far_0_779_1;    relay_conn far_0_779_1_a(.in(far_0_779_0[0]), .out(far_0_779_1[0]));    relay_conn far_0_779_1_b(.in(far_0_779_0[1]), .out(far_0_779_1[1]));
    assign layer_0[779] = ~far_0_779_1[1] | (far_0_779_1[0] & far_0_779_1[1]); 
    assign layer_0[780] = ~(in[127] ^ in[97]); 
    assign layer_0[781] = in[125] & in[148]; 
    wire [1:0] far_0_782_0;    relay_conn far_0_782_0_a(.in(in[111]), .out(far_0_782_0[0]));    relay_conn far_0_782_0_b(.in(in[34]), .out(far_0_782_0[1]));
    wire [1:0] far_0_782_1;    relay_conn far_0_782_1_a(.in(far_0_782_0[0]), .out(far_0_782_1[0]));    relay_conn far_0_782_1_b(.in(far_0_782_0[1]), .out(far_0_782_1[1]));
    assign layer_0[782] = far_0_782_1[0] & far_0_782_1[1]; 
    wire [1:0] far_0_783_0;    relay_conn far_0_783_0_a(.in(in[79]), .out(far_0_783_0[0]));    relay_conn far_0_783_0_b(.in(in[33]), .out(far_0_783_0[1]));
    assign layer_0[783] = far_0_783_0[0] & ~far_0_783_0[1]; 
    wire [1:0] far_0_784_0;    relay_conn far_0_784_0_a(.in(in[241]), .out(far_0_784_0[0]));    relay_conn far_0_784_0_b(.in(in[199]), .out(far_0_784_0[1]));
    assign layer_0[784] = ~far_0_784_0[1]; 
    wire [1:0] far_0_785_0;    relay_conn far_0_785_0_a(.in(in[125]), .out(far_0_785_0[0]));    relay_conn far_0_785_0_b(.in(in[223]), .out(far_0_785_0[1]));
    wire [1:0] far_0_785_1;    relay_conn far_0_785_1_a(.in(far_0_785_0[0]), .out(far_0_785_1[0]));    relay_conn far_0_785_1_b(.in(far_0_785_0[1]), .out(far_0_785_1[1]));
    wire [1:0] far_0_785_2;    relay_conn far_0_785_2_a(.in(far_0_785_1[0]), .out(far_0_785_2[0]));    relay_conn far_0_785_2_b(.in(far_0_785_1[1]), .out(far_0_785_2[1]));
    assign layer_0[785] = ~(far_0_785_2[0] & far_0_785_2[1]); 
    wire [1:0] far_0_786_0;    relay_conn far_0_786_0_a(.in(in[121]), .out(far_0_786_0[0]));    relay_conn far_0_786_0_b(.in(in[197]), .out(far_0_786_0[1]));
    wire [1:0] far_0_786_1;    relay_conn far_0_786_1_a(.in(far_0_786_0[0]), .out(far_0_786_1[0]));    relay_conn far_0_786_1_b(.in(far_0_786_0[1]), .out(far_0_786_1[1]));
    assign layer_0[786] = far_0_786_1[0] | far_0_786_1[1]; 
    wire [1:0] far_0_787_0;    relay_conn far_0_787_0_a(.in(in[109]), .out(far_0_787_0[0]));    relay_conn far_0_787_0_b(.in(in[199]), .out(far_0_787_0[1]));
    wire [1:0] far_0_787_1;    relay_conn far_0_787_1_a(.in(far_0_787_0[0]), .out(far_0_787_1[0]));    relay_conn far_0_787_1_b(.in(far_0_787_0[1]), .out(far_0_787_1[1]));
    assign layer_0[787] = ~far_0_787_1[1] | (far_0_787_1[0] & far_0_787_1[1]); 
    wire [1:0] far_0_788_0;    relay_conn far_0_788_0_a(.in(in[34]), .out(far_0_788_0[0]));    relay_conn far_0_788_0_b(.in(in[87]), .out(far_0_788_0[1]));
    assign layer_0[788] = ~far_0_788_0[0]; 
    wire [1:0] far_0_789_0;    relay_conn far_0_789_0_a(.in(in[172]), .out(far_0_789_0[0]));    relay_conn far_0_789_0_b(.in(in[125]), .out(far_0_789_0[1]));
    assign layer_0[789] = ~far_0_789_0[1]; 
    wire [1:0] far_0_790_0;    relay_conn far_0_790_0_a(.in(in[92]), .out(far_0_790_0[0]));    relay_conn far_0_790_0_b(.in(in[150]), .out(far_0_790_0[1]));
    assign layer_0[790] = far_0_790_0[0] ^ far_0_790_0[1]; 
    wire [1:0] far_0_791_0;    relay_conn far_0_791_0_a(.in(in[104]), .out(far_0_791_0[0]));    relay_conn far_0_791_0_b(.in(in[170]), .out(far_0_791_0[1]));
    wire [1:0] far_0_791_1;    relay_conn far_0_791_1_a(.in(far_0_791_0[0]), .out(far_0_791_1[0]));    relay_conn far_0_791_1_b(.in(far_0_791_0[1]), .out(far_0_791_1[1]));
    assign layer_0[791] = far_0_791_1[0] & ~far_0_791_1[1]; 
    assign layer_0[792] = in[161] ^ in[186]; 
    wire [1:0] far_0_793_0;    relay_conn far_0_793_0_a(.in(in[187]), .out(far_0_793_0[0]));    relay_conn far_0_793_0_b(.in(in[251]), .out(far_0_793_0[1]));
    wire [1:0] far_0_793_1;    relay_conn far_0_793_1_a(.in(far_0_793_0[0]), .out(far_0_793_1[0]));    relay_conn far_0_793_1_b(.in(far_0_793_0[1]), .out(far_0_793_1[1]));
    assign layer_0[793] = ~far_0_793_1[1] | (far_0_793_1[0] & far_0_793_1[1]); 
    wire [1:0] far_0_794_0;    relay_conn far_0_794_0_a(.in(in[85]), .out(far_0_794_0[0]));    relay_conn far_0_794_0_b(.in(in[34]), .out(far_0_794_0[1]));
    assign layer_0[794] = far_0_794_0[0]; 
    wire [1:0] far_0_795_0;    relay_conn far_0_795_0_a(.in(in[113]), .out(far_0_795_0[0]));    relay_conn far_0_795_0_b(.in(in[74]), .out(far_0_795_0[1]));
    assign layer_0[795] = far_0_795_0[1]; 
    wire [1:0] far_0_796_0;    relay_conn far_0_796_0_a(.in(in[151]), .out(far_0_796_0[0]));    relay_conn far_0_796_0_b(.in(in[247]), .out(far_0_796_0[1]));
    wire [1:0] far_0_796_1;    relay_conn far_0_796_1_a(.in(far_0_796_0[0]), .out(far_0_796_1[0]));    relay_conn far_0_796_1_b(.in(far_0_796_0[1]), .out(far_0_796_1[1]));
    wire [1:0] far_0_796_2;    relay_conn far_0_796_2_a(.in(far_0_796_1[0]), .out(far_0_796_2[0]));    relay_conn far_0_796_2_b(.in(far_0_796_1[1]), .out(far_0_796_2[1]));
    assign layer_0[796] = far_0_796_2[1] & ~far_0_796_2[0]; 
    wire [1:0] far_0_797_0;    relay_conn far_0_797_0_a(.in(in[99]), .out(far_0_797_0[0]));    relay_conn far_0_797_0_b(.in(in[66]), .out(far_0_797_0[1]));
    assign layer_0[797] = far_0_797_0[0] & ~far_0_797_0[1]; 
    assign layer_0[798] = ~(in[99] & in[97]); 
    wire [1:0] far_0_799_0;    relay_conn far_0_799_0_a(.in(in[151]), .out(far_0_799_0[0]));    relay_conn far_0_799_0_b(.in(in[72]), .out(far_0_799_0[1]));
    wire [1:0] far_0_799_1;    relay_conn far_0_799_1_a(.in(far_0_799_0[0]), .out(far_0_799_1[0]));    relay_conn far_0_799_1_b(.in(far_0_799_0[1]), .out(far_0_799_1[1]));
    assign layer_0[799] = ~far_0_799_1[0] | (far_0_799_1[0] & far_0_799_1[1]); 
    wire [1:0] far_0_800_0;    relay_conn far_0_800_0_a(.in(in[243]), .out(far_0_800_0[0]));    relay_conn far_0_800_0_b(.in(in[157]), .out(far_0_800_0[1]));
    wire [1:0] far_0_800_1;    relay_conn far_0_800_1_a(.in(far_0_800_0[0]), .out(far_0_800_1[0]));    relay_conn far_0_800_1_b(.in(far_0_800_0[1]), .out(far_0_800_1[1]));
    assign layer_0[800] = ~(far_0_800_1[0] & far_0_800_1[1]); 
    assign layer_0[801] = in[130] ^ in[157]; 
    wire [1:0] far_0_802_0;    relay_conn far_0_802_0_a(.in(in[143]), .out(far_0_802_0[0]));    relay_conn far_0_802_0_b(.in(in[101]), .out(far_0_802_0[1]));
    assign layer_0[802] = far_0_802_0[0] | far_0_802_0[1]; 
    wire [1:0] far_0_803_0;    relay_conn far_0_803_0_a(.in(in[74]), .out(far_0_803_0[0]));    relay_conn far_0_803_0_b(.in(in[116]), .out(far_0_803_0[1]));
    assign layer_0[803] = far_0_803_0[0]; 
    wire [1:0] far_0_804_0;    relay_conn far_0_804_0_a(.in(in[162]), .out(far_0_804_0[0]));    relay_conn far_0_804_0_b(.in(in[110]), .out(far_0_804_0[1]));
    assign layer_0[804] = far_0_804_0[1] & ~far_0_804_0[0]; 
    assign layer_0[805] = in[121] | in[99]; 
    assign layer_0[806] = ~in[88] | (in[77] & in[88]); 
    wire [1:0] far_0_807_0;    relay_conn far_0_807_0_a(.in(in[61]), .out(far_0_807_0[0]));    relay_conn far_0_807_0_b(.in(in[165]), .out(far_0_807_0[1]));
    wire [1:0] far_0_807_1;    relay_conn far_0_807_1_a(.in(far_0_807_0[0]), .out(far_0_807_1[0]));    relay_conn far_0_807_1_b(.in(far_0_807_0[1]), .out(far_0_807_1[1]));
    wire [1:0] far_0_807_2;    relay_conn far_0_807_2_a(.in(far_0_807_1[0]), .out(far_0_807_2[0]));    relay_conn far_0_807_2_b(.in(far_0_807_1[1]), .out(far_0_807_2[1]));
    assign layer_0[807] = far_0_807_2[0] | far_0_807_2[1]; 
    wire [1:0] far_0_808_0;    relay_conn far_0_808_0_a(.in(in[53]), .out(far_0_808_0[0]));    relay_conn far_0_808_0_b(.in(in[158]), .out(far_0_808_0[1]));
    wire [1:0] far_0_808_1;    relay_conn far_0_808_1_a(.in(far_0_808_0[0]), .out(far_0_808_1[0]));    relay_conn far_0_808_1_b(.in(far_0_808_0[1]), .out(far_0_808_1[1]));
    wire [1:0] far_0_808_2;    relay_conn far_0_808_2_a(.in(far_0_808_1[0]), .out(far_0_808_2[0]));    relay_conn far_0_808_2_b(.in(far_0_808_1[1]), .out(far_0_808_2[1]));
    assign layer_0[808] = far_0_808_2[0] | far_0_808_2[1]; 
    wire [1:0] far_0_809_0;    relay_conn far_0_809_0_a(.in(in[88]), .out(far_0_809_0[0]));    relay_conn far_0_809_0_b(.in(in[48]), .out(far_0_809_0[1]));
    assign layer_0[809] = far_0_809_0[1] & ~far_0_809_0[0]; 
    assign layer_0[810] = ~(in[188] | in[213]); 
    wire [1:0] far_0_811_0;    relay_conn far_0_811_0_a(.in(in[109]), .out(far_0_811_0[0]));    relay_conn far_0_811_0_b(.in(in[34]), .out(far_0_811_0[1]));
    wire [1:0] far_0_811_1;    relay_conn far_0_811_1_a(.in(far_0_811_0[0]), .out(far_0_811_1[0]));    relay_conn far_0_811_1_b(.in(far_0_811_0[1]), .out(far_0_811_1[1]));
    assign layer_0[811] = far_0_811_1[0] & far_0_811_1[1]; 
    wire [1:0] far_0_812_0;    relay_conn far_0_812_0_a(.in(in[15]), .out(far_0_812_0[0]));    relay_conn far_0_812_0_b(.in(in[113]), .out(far_0_812_0[1]));
    wire [1:0] far_0_812_1;    relay_conn far_0_812_1_a(.in(far_0_812_0[0]), .out(far_0_812_1[0]));    relay_conn far_0_812_1_b(.in(far_0_812_0[1]), .out(far_0_812_1[1]));
    wire [1:0] far_0_812_2;    relay_conn far_0_812_2_a(.in(far_0_812_1[0]), .out(far_0_812_2[0]));    relay_conn far_0_812_2_b(.in(far_0_812_1[1]), .out(far_0_812_2[1]));
    assign layer_0[812] = far_0_812_2[0] | far_0_812_2[1]; 
    assign layer_0[813] = in[17]; 
    assign layer_0[814] = ~(in[204] ^ in[207]); 
    wire [1:0] far_0_815_0;    relay_conn far_0_815_0_a(.in(in[30]), .out(far_0_815_0[0]));    relay_conn far_0_815_0_b(.in(in[158]), .out(far_0_815_0[1]));
    wire [1:0] far_0_815_1;    relay_conn far_0_815_1_a(.in(far_0_815_0[0]), .out(far_0_815_1[0]));    relay_conn far_0_815_1_b(.in(far_0_815_0[1]), .out(far_0_815_1[1]));
    wire [1:0] far_0_815_2;    relay_conn far_0_815_2_a(.in(far_0_815_1[0]), .out(far_0_815_2[0]));    relay_conn far_0_815_2_b(.in(far_0_815_1[1]), .out(far_0_815_2[1]));
    wire [1:0] far_0_815_3;    relay_conn far_0_815_3_a(.in(far_0_815_2[0]), .out(far_0_815_3[0]));    relay_conn far_0_815_3_b(.in(far_0_815_2[1]), .out(far_0_815_3[1]));
    assign layer_0[815] = ~far_0_815_3[0] | (far_0_815_3[0] & far_0_815_3[1]); 
    assign layer_0[816] = in[87] & in[112]; 
    assign layer_0[817] = in[229]; 
    assign layer_0[818] = ~in[197] | (in[167] & in[197]); 
    wire [1:0] far_0_819_0;    relay_conn far_0_819_0_a(.in(in[30]), .out(far_0_819_0[0]));    relay_conn far_0_819_0_b(.in(in[71]), .out(far_0_819_0[1]));
    assign layer_0[819] = ~far_0_819_0[0]; 
    wire [1:0] far_0_820_0;    relay_conn far_0_820_0_a(.in(in[150]), .out(far_0_820_0[0]));    relay_conn far_0_820_0_b(.in(in[62]), .out(far_0_820_0[1]));
    wire [1:0] far_0_820_1;    relay_conn far_0_820_1_a(.in(far_0_820_0[0]), .out(far_0_820_1[0]));    relay_conn far_0_820_1_b(.in(far_0_820_0[1]), .out(far_0_820_1[1]));
    assign layer_0[820] = ~far_0_820_1[1]; 
    wire [1:0] far_0_821_0;    relay_conn far_0_821_0_a(.in(in[120]), .out(far_0_821_0[0]));    relay_conn far_0_821_0_b(.in(in[179]), .out(far_0_821_0[1]));
    assign layer_0[821] = far_0_821_0[0]; 
    assign layer_0[822] = ~in[109] | (in[95] & in[109]); 
    assign layer_0[823] = ~(in[73] ^ in[48]); 
    wire [1:0] far_0_824_0;    relay_conn far_0_824_0_a(.in(in[185]), .out(far_0_824_0[0]));    relay_conn far_0_824_0_b(.in(in[97]), .out(far_0_824_0[1]));
    wire [1:0] far_0_824_1;    relay_conn far_0_824_1_a(.in(far_0_824_0[0]), .out(far_0_824_1[0]));    relay_conn far_0_824_1_b(.in(far_0_824_0[1]), .out(far_0_824_1[1]));
    assign layer_0[824] = ~far_0_824_1[0] | (far_0_824_1[0] & far_0_824_1[1]); 
    wire [1:0] far_0_825_0;    relay_conn far_0_825_0_a(.in(in[15]), .out(far_0_825_0[0]));    relay_conn far_0_825_0_b(.in(in[132]), .out(far_0_825_0[1]));
    wire [1:0] far_0_825_1;    relay_conn far_0_825_1_a(.in(far_0_825_0[0]), .out(far_0_825_1[0]));    relay_conn far_0_825_1_b(.in(far_0_825_0[1]), .out(far_0_825_1[1]));
    wire [1:0] far_0_825_2;    relay_conn far_0_825_2_a(.in(far_0_825_1[0]), .out(far_0_825_2[0]));    relay_conn far_0_825_2_b(.in(far_0_825_1[1]), .out(far_0_825_2[1]));
    assign layer_0[825] = ~(far_0_825_2[0] & far_0_825_2[1]); 
    assign layer_0[826] = ~(in[109] | in[93]); 
    wire [1:0] far_0_827_0;    relay_conn far_0_827_0_a(.in(in[238]), .out(far_0_827_0[0]));    relay_conn far_0_827_0_b(.in(in[173]), .out(far_0_827_0[1]));
    wire [1:0] far_0_827_1;    relay_conn far_0_827_1_a(.in(far_0_827_0[0]), .out(far_0_827_1[0]));    relay_conn far_0_827_1_b(.in(far_0_827_0[1]), .out(far_0_827_1[1]));
    assign layer_0[827] = ~far_0_827_1[0]; 
    wire [1:0] far_0_828_0;    relay_conn far_0_828_0_a(.in(in[202]), .out(far_0_828_0[0]));    relay_conn far_0_828_0_b(.in(in[239]), .out(far_0_828_0[1]));
    assign layer_0[828] = far_0_828_0[1] & ~far_0_828_0[0]; 
    wire [1:0] far_0_829_0;    relay_conn far_0_829_0_a(.in(in[110]), .out(far_0_829_0[0]));    relay_conn far_0_829_0_b(.in(in[71]), .out(far_0_829_0[1]));
    assign layer_0[829] = far_0_829_0[0] & far_0_829_0[1]; 
    assign layer_0[830] = ~(in[186] ^ in[210]); 
    assign layer_0[831] = ~in[22] | (in[52] & in[22]); 
    wire [1:0] far_0_832_0;    relay_conn far_0_832_0_a(.in(in[44]), .out(far_0_832_0[0]));    relay_conn far_0_832_0_b(.in(in[125]), .out(far_0_832_0[1]));
    wire [1:0] far_0_832_1;    relay_conn far_0_832_1_a(.in(far_0_832_0[0]), .out(far_0_832_1[0]));    relay_conn far_0_832_1_b(.in(far_0_832_0[1]), .out(far_0_832_1[1]));
    assign layer_0[832] = far_0_832_1[0] | far_0_832_1[1]; 
    wire [1:0] far_0_833_0;    relay_conn far_0_833_0_a(.in(in[67]), .out(far_0_833_0[0]));    relay_conn far_0_833_0_b(.in(in[13]), .out(far_0_833_0[1]));
    assign layer_0[833] = ~(far_0_833_0[0] & far_0_833_0[1]); 
    wire [1:0] far_0_834_0;    relay_conn far_0_834_0_a(.in(in[90]), .out(far_0_834_0[0]));    relay_conn far_0_834_0_b(.in(in[213]), .out(far_0_834_0[1]));
    wire [1:0] far_0_834_1;    relay_conn far_0_834_1_a(.in(far_0_834_0[0]), .out(far_0_834_1[0]));    relay_conn far_0_834_1_b(.in(far_0_834_0[1]), .out(far_0_834_1[1]));
    wire [1:0] far_0_834_2;    relay_conn far_0_834_2_a(.in(far_0_834_1[0]), .out(far_0_834_2[0]));    relay_conn far_0_834_2_b(.in(far_0_834_1[1]), .out(far_0_834_2[1]));
    assign layer_0[834] = ~far_0_834_2[0] | (far_0_834_2[0] & far_0_834_2[1]); 
    wire [1:0] far_0_835_0;    relay_conn far_0_835_0_a(.in(in[216]), .out(far_0_835_0[0]));    relay_conn far_0_835_0_b(.in(in[134]), .out(far_0_835_0[1]));
    wire [1:0] far_0_835_1;    relay_conn far_0_835_1_a(.in(far_0_835_0[0]), .out(far_0_835_1[0]));    relay_conn far_0_835_1_b(.in(far_0_835_0[1]), .out(far_0_835_1[1]));
    assign layer_0[835] = ~far_0_835_1[1] | (far_0_835_1[0] & far_0_835_1[1]); 
    assign layer_0[836] = in[142] & ~in[122]; 
    wire [1:0] far_0_837_0;    relay_conn far_0_837_0_a(.in(in[130]), .out(far_0_837_0[0]));    relay_conn far_0_837_0_b(.in(in[89]), .out(far_0_837_0[1]));
    assign layer_0[837] = far_0_837_0[0] & far_0_837_0[1]; 
    wire [1:0] far_0_838_0;    relay_conn far_0_838_0_a(.in(in[239]), .out(far_0_838_0[0]));    relay_conn far_0_838_0_b(.in(in[117]), .out(far_0_838_0[1]));
    wire [1:0] far_0_838_1;    relay_conn far_0_838_1_a(.in(far_0_838_0[0]), .out(far_0_838_1[0]));    relay_conn far_0_838_1_b(.in(far_0_838_0[1]), .out(far_0_838_1[1]));
    wire [1:0] far_0_838_2;    relay_conn far_0_838_2_a(.in(far_0_838_1[0]), .out(far_0_838_2[0]));    relay_conn far_0_838_2_b(.in(far_0_838_1[1]), .out(far_0_838_2[1]));
    assign layer_0[838] = ~far_0_838_2[0] | (far_0_838_2[0] & far_0_838_2[1]); 
    wire [1:0] far_0_839_0;    relay_conn far_0_839_0_a(.in(in[34]), .out(far_0_839_0[0]));    relay_conn far_0_839_0_b(.in(in[151]), .out(far_0_839_0[1]));
    wire [1:0] far_0_839_1;    relay_conn far_0_839_1_a(.in(far_0_839_0[0]), .out(far_0_839_1[0]));    relay_conn far_0_839_1_b(.in(far_0_839_0[1]), .out(far_0_839_1[1]));
    wire [1:0] far_0_839_2;    relay_conn far_0_839_2_a(.in(far_0_839_1[0]), .out(far_0_839_2[0]));    relay_conn far_0_839_2_b(.in(far_0_839_1[1]), .out(far_0_839_2[1]));
    assign layer_0[839] = far_0_839_2[1] & ~far_0_839_2[0]; 
    assign layer_0[840] = in[91] & ~in[75]; 
    wire [1:0] far_0_841_0;    relay_conn far_0_841_0_a(.in(in[223]), .out(far_0_841_0[0]));    relay_conn far_0_841_0_b(.in(in[175]), .out(far_0_841_0[1]));
    assign layer_0[841] = far_0_841_0[0] & far_0_841_0[1]; 
    wire [1:0] far_0_842_0;    relay_conn far_0_842_0_a(.in(in[150]), .out(far_0_842_0[0]));    relay_conn far_0_842_0_b(.in(in[37]), .out(far_0_842_0[1]));
    wire [1:0] far_0_842_1;    relay_conn far_0_842_1_a(.in(far_0_842_0[0]), .out(far_0_842_1[0]));    relay_conn far_0_842_1_b(.in(far_0_842_0[1]), .out(far_0_842_1[1]));
    wire [1:0] far_0_842_2;    relay_conn far_0_842_2_a(.in(far_0_842_1[0]), .out(far_0_842_2[0]));    relay_conn far_0_842_2_b(.in(far_0_842_1[1]), .out(far_0_842_2[1]));
    assign layer_0[842] = far_0_842_2[0] | far_0_842_2[1]; 
    assign layer_0[843] = ~in[82]; 
    wire [1:0] far_0_844_0;    relay_conn far_0_844_0_a(.in(in[239]), .out(far_0_844_0[0]));    relay_conn far_0_844_0_b(.in(in[115]), .out(far_0_844_0[1]));
    wire [1:0] far_0_844_1;    relay_conn far_0_844_1_a(.in(far_0_844_0[0]), .out(far_0_844_1[0]));    relay_conn far_0_844_1_b(.in(far_0_844_0[1]), .out(far_0_844_1[1]));
    wire [1:0] far_0_844_2;    relay_conn far_0_844_2_a(.in(far_0_844_1[0]), .out(far_0_844_2[0]));    relay_conn far_0_844_2_b(.in(far_0_844_1[1]), .out(far_0_844_2[1]));
    assign layer_0[844] = ~far_0_844_2[1] | (far_0_844_2[0] & far_0_844_2[1]); 
    assign layer_0[845] = ~(in[72] ^ in[68]); 
    assign layer_0[846] = ~in[159]; 
    assign layer_0[847] = in[204]; 
    assign layer_0[848] = ~in[203] | (in[233] & in[203]); 
    wire [1:0] far_0_849_0;    relay_conn far_0_849_0_a(.in(in[127]), .out(far_0_849_0[0]));    relay_conn far_0_849_0_b(.in(in[51]), .out(far_0_849_0[1]));
    wire [1:0] far_0_849_1;    relay_conn far_0_849_1_a(.in(far_0_849_0[0]), .out(far_0_849_1[0]));    relay_conn far_0_849_1_b(.in(far_0_849_0[1]), .out(far_0_849_1[1]));
    assign layer_0[849] = far_0_849_1[0]; 
    wire [1:0] far_0_850_0;    relay_conn far_0_850_0_a(.in(in[76]), .out(far_0_850_0[0]));    relay_conn far_0_850_0_b(.in(in[130]), .out(far_0_850_0[1]));
    assign layer_0[850] = ~(far_0_850_0[0] & far_0_850_0[1]); 
    assign layer_0[851] = ~in[158] | (in[172] & in[158]); 
    wire [1:0] far_0_852_0;    relay_conn far_0_852_0_a(.in(in[151]), .out(far_0_852_0[0]));    relay_conn far_0_852_0_b(.in(in[215]), .out(far_0_852_0[1]));
    wire [1:0] far_0_852_1;    relay_conn far_0_852_1_a(.in(far_0_852_0[0]), .out(far_0_852_1[0]));    relay_conn far_0_852_1_b(.in(far_0_852_0[1]), .out(far_0_852_1[1]));
    assign layer_0[852] = ~(far_0_852_1[0] & far_0_852_1[1]); 
    wire [1:0] far_0_853_0;    relay_conn far_0_853_0_a(.in(in[18]), .out(far_0_853_0[0]));    relay_conn far_0_853_0_b(.in(in[111]), .out(far_0_853_0[1]));
    wire [1:0] far_0_853_1;    relay_conn far_0_853_1_a(.in(far_0_853_0[0]), .out(far_0_853_1[0]));    relay_conn far_0_853_1_b(.in(far_0_853_0[1]), .out(far_0_853_1[1]));
    assign layer_0[853] = ~(far_0_853_1[0] | far_0_853_1[1]); 
    wire [1:0] far_0_854_0;    relay_conn far_0_854_0_a(.in(in[57]), .out(far_0_854_0[0]));    relay_conn far_0_854_0_b(.in(in[175]), .out(far_0_854_0[1]));
    wire [1:0] far_0_854_1;    relay_conn far_0_854_1_a(.in(far_0_854_0[0]), .out(far_0_854_1[0]));    relay_conn far_0_854_1_b(.in(far_0_854_0[1]), .out(far_0_854_1[1]));
    wire [1:0] far_0_854_2;    relay_conn far_0_854_2_a(.in(far_0_854_1[0]), .out(far_0_854_2[0]));    relay_conn far_0_854_2_b(.in(far_0_854_1[1]), .out(far_0_854_2[1]));
    assign layer_0[854] = ~(far_0_854_2[0] ^ far_0_854_2[1]); 
    wire [1:0] far_0_855_0;    relay_conn far_0_855_0_a(.in(in[88]), .out(far_0_855_0[0]));    relay_conn far_0_855_0_b(.in(in[191]), .out(far_0_855_0[1]));
    wire [1:0] far_0_855_1;    relay_conn far_0_855_1_a(.in(far_0_855_0[0]), .out(far_0_855_1[0]));    relay_conn far_0_855_1_b(.in(far_0_855_0[1]), .out(far_0_855_1[1]));
    wire [1:0] far_0_855_2;    relay_conn far_0_855_2_a(.in(far_0_855_1[0]), .out(far_0_855_2[0]));    relay_conn far_0_855_2_b(.in(far_0_855_1[1]), .out(far_0_855_2[1]));
    assign layer_0[855] = ~far_0_855_2[0]; 
    wire [1:0] far_0_856_0;    relay_conn far_0_856_0_a(.in(in[94]), .out(far_0_856_0[0]));    relay_conn far_0_856_0_b(.in(in[133]), .out(far_0_856_0[1]));
    assign layer_0[856] = ~(far_0_856_0[0] ^ far_0_856_0[1]); 
    wire [1:0] far_0_857_0;    relay_conn far_0_857_0_a(.in(in[55]), .out(far_0_857_0[0]));    relay_conn far_0_857_0_b(.in(in[151]), .out(far_0_857_0[1]));
    wire [1:0] far_0_857_1;    relay_conn far_0_857_1_a(.in(far_0_857_0[0]), .out(far_0_857_1[0]));    relay_conn far_0_857_1_b(.in(far_0_857_0[1]), .out(far_0_857_1[1]));
    wire [1:0] far_0_857_2;    relay_conn far_0_857_2_a(.in(far_0_857_1[0]), .out(far_0_857_2[0]));    relay_conn far_0_857_2_b(.in(far_0_857_1[1]), .out(far_0_857_2[1]));
    assign layer_0[857] = ~far_0_857_2[1]; 
    wire [1:0] far_0_858_0;    relay_conn far_0_858_0_a(.in(in[63]), .out(far_0_858_0[0]));    relay_conn far_0_858_0_b(.in(in[153]), .out(far_0_858_0[1]));
    wire [1:0] far_0_858_1;    relay_conn far_0_858_1_a(.in(far_0_858_0[0]), .out(far_0_858_1[0]));    relay_conn far_0_858_1_b(.in(far_0_858_0[1]), .out(far_0_858_1[1]));
    assign layer_0[858] = ~(far_0_858_1[0] & far_0_858_1[1]); 
    wire [1:0] far_0_859_0;    relay_conn far_0_859_0_a(.in(in[79]), .out(far_0_859_0[0]));    relay_conn far_0_859_0_b(.in(in[28]), .out(far_0_859_0[1]));
    assign layer_0[859] = ~far_0_859_0[0]; 
    wire [1:0] far_0_860_0;    relay_conn far_0_860_0_a(.in(in[64]), .out(far_0_860_0[0]));    relay_conn far_0_860_0_b(.in(in[157]), .out(far_0_860_0[1]));
    wire [1:0] far_0_860_1;    relay_conn far_0_860_1_a(.in(far_0_860_0[0]), .out(far_0_860_1[0]));    relay_conn far_0_860_1_b(.in(far_0_860_0[1]), .out(far_0_860_1[1]));
    assign layer_0[860] = far_0_860_1[0]; 
    assign layer_0[861] = ~in[26]; 
    wire [1:0] far_0_862_0;    relay_conn far_0_862_0_a(.in(in[157]), .out(far_0_862_0[0]));    relay_conn far_0_862_0_b(.in(in[57]), .out(far_0_862_0[1]));
    wire [1:0] far_0_862_1;    relay_conn far_0_862_1_a(.in(far_0_862_0[0]), .out(far_0_862_1[0]));    relay_conn far_0_862_1_b(.in(far_0_862_0[1]), .out(far_0_862_1[1]));
    wire [1:0] far_0_862_2;    relay_conn far_0_862_2_a(.in(far_0_862_1[0]), .out(far_0_862_2[0]));    relay_conn far_0_862_2_b(.in(far_0_862_1[1]), .out(far_0_862_2[1]));
    assign layer_0[862] = far_0_862_2[0]; 
    assign layer_0[863] = ~(in[101] | in[90]); 
    assign layer_0[864] = ~(in[186] | in[174]); 
    wire [1:0] far_0_865_0;    relay_conn far_0_865_0_a(.in(in[132]), .out(far_0_865_0[0]));    relay_conn far_0_865_0_b(.in(in[17]), .out(far_0_865_0[1]));
    wire [1:0] far_0_865_1;    relay_conn far_0_865_1_a(.in(far_0_865_0[0]), .out(far_0_865_1[0]));    relay_conn far_0_865_1_b(.in(far_0_865_0[1]), .out(far_0_865_1[1]));
    wire [1:0] far_0_865_2;    relay_conn far_0_865_2_a(.in(far_0_865_1[0]), .out(far_0_865_2[0]));    relay_conn far_0_865_2_b(.in(far_0_865_1[1]), .out(far_0_865_2[1]));
    assign layer_0[865] = far_0_865_2[0] & far_0_865_2[1]; 
    assign layer_0[866] = in[203] & ~in[186]; 
    wire [1:0] far_0_867_0;    relay_conn far_0_867_0_a(.in(in[239]), .out(far_0_867_0[0]));    relay_conn far_0_867_0_b(.in(in[157]), .out(far_0_867_0[1]));
    wire [1:0] far_0_867_1;    relay_conn far_0_867_1_a(.in(far_0_867_0[0]), .out(far_0_867_1[0]));    relay_conn far_0_867_1_b(.in(far_0_867_0[1]), .out(far_0_867_1[1]));
    assign layer_0[867] = ~far_0_867_1[0] | (far_0_867_1[0] & far_0_867_1[1]); 
    assign layer_0[868] = in[136] | in[122]; 
    assign layer_0[869] = ~in[199]; 
    wire [1:0] far_0_870_0;    relay_conn far_0_870_0_a(.in(in[179]), .out(far_0_870_0[0]));    relay_conn far_0_870_0_b(.in(in[212]), .out(far_0_870_0[1]));
    assign layer_0[870] = far_0_870_0[0] & ~far_0_870_0[1]; 
    assign layer_0[871] = in[41] & ~in[57]; 
    wire [1:0] far_0_872_0;    relay_conn far_0_872_0_a(.in(in[164]), .out(far_0_872_0[0]));    relay_conn far_0_872_0_b(.in(in[99]), .out(far_0_872_0[1]));
    wire [1:0] far_0_872_1;    relay_conn far_0_872_1_a(.in(far_0_872_0[0]), .out(far_0_872_1[0]));    relay_conn far_0_872_1_b(.in(far_0_872_0[1]), .out(far_0_872_1[1]));
    assign layer_0[872] = ~far_0_872_1[0] | (far_0_872_1[0] & far_0_872_1[1]); 
    wire [1:0] far_0_873_0;    relay_conn far_0_873_0_a(.in(in[156]), .out(far_0_873_0[0]));    relay_conn far_0_873_0_b(.in(in[252]), .out(far_0_873_0[1]));
    wire [1:0] far_0_873_1;    relay_conn far_0_873_1_a(.in(far_0_873_0[0]), .out(far_0_873_1[0]));    relay_conn far_0_873_1_b(.in(far_0_873_0[1]), .out(far_0_873_1[1]));
    wire [1:0] far_0_873_2;    relay_conn far_0_873_2_a(.in(far_0_873_1[0]), .out(far_0_873_2[0]));    relay_conn far_0_873_2_b(.in(far_0_873_1[1]), .out(far_0_873_2[1]));
    assign layer_0[873] = far_0_873_2[1]; 
    wire [1:0] far_0_874_0;    relay_conn far_0_874_0_a(.in(in[138]), .out(far_0_874_0[0]));    relay_conn far_0_874_0_b(.in(in[187]), .out(far_0_874_0[1]));
    assign layer_0[874] = ~far_0_874_0[0]; 
    assign layer_0[875] = ~(in[82] | in[79]); 
    assign layer_0[876] = in[202] & ~in[196]; 
    wire [1:0] far_0_877_0;    relay_conn far_0_877_0_a(.in(in[117]), .out(far_0_877_0[0]));    relay_conn far_0_877_0_b(.in(in[45]), .out(far_0_877_0[1]));
    wire [1:0] far_0_877_1;    relay_conn far_0_877_1_a(.in(far_0_877_0[0]), .out(far_0_877_1[0]));    relay_conn far_0_877_1_b(.in(far_0_877_0[1]), .out(far_0_877_1[1]));
    assign layer_0[877] = far_0_877_1[1] & ~far_0_877_1[0]; 
    wire [1:0] far_0_878_0;    relay_conn far_0_878_0_a(.in(in[17]), .out(far_0_878_0[0]));    relay_conn far_0_878_0_b(.in(in[59]), .out(far_0_878_0[1]));
    assign layer_0[878] = ~far_0_878_0[0] | (far_0_878_0[0] & far_0_878_0[1]); 
    assign layer_0[879] = in[165] & in[186]; 
    wire [1:0] far_0_880_0;    relay_conn far_0_880_0_a(.in(in[95]), .out(far_0_880_0[0]));    relay_conn far_0_880_0_b(.in(in[34]), .out(far_0_880_0[1]));
    assign layer_0[880] = far_0_880_0[0] & ~far_0_880_0[1]; 
    wire [1:0] far_0_881_0;    relay_conn far_0_881_0_a(.in(in[51]), .out(far_0_881_0[0]));    relay_conn far_0_881_0_b(.in(in[112]), .out(far_0_881_0[1]));
    assign layer_0[881] = far_0_881_0[1]; 
    wire [1:0] far_0_882_0;    relay_conn far_0_882_0_a(.in(in[190]), .out(far_0_882_0[0]));    relay_conn far_0_882_0_b(.in(in[150]), .out(far_0_882_0[1]));
    assign layer_0[882] = ~far_0_882_0[0] | (far_0_882_0[0] & far_0_882_0[1]); 
    wire [1:0] far_0_883_0;    relay_conn far_0_883_0_a(.in(in[204]), .out(far_0_883_0[0]));    relay_conn far_0_883_0_b(.in(in[150]), .out(far_0_883_0[1]));
    assign layer_0[883] = far_0_883_0[0] ^ far_0_883_0[1]; 
    assign layer_0[884] = ~in[150]; 
    wire [1:0] far_0_885_0;    relay_conn far_0_885_0_a(.in(in[74]), .out(far_0_885_0[0]));    relay_conn far_0_885_0_b(.in(in[149]), .out(far_0_885_0[1]));
    wire [1:0] far_0_885_1;    relay_conn far_0_885_1_a(.in(far_0_885_0[0]), .out(far_0_885_1[0]));    relay_conn far_0_885_1_b(.in(far_0_885_0[1]), .out(far_0_885_1[1]));
    assign layer_0[885] = ~(far_0_885_1[0] ^ far_0_885_1[1]); 
    assign layer_0[886] = in[44] & ~in[17]; 
    assign layer_0[887] = ~in[197]; 
    assign layer_0[888] = in[221]; 
    wire [1:0] far_0_889_0;    relay_conn far_0_889_0_a(.in(in[68]), .out(far_0_889_0[0]));    relay_conn far_0_889_0_b(.in(in[122]), .out(far_0_889_0[1]));
    assign layer_0[889] = far_0_889_0[1] & ~far_0_889_0[0]; 
    wire [1:0] far_0_890_0;    relay_conn far_0_890_0_a(.in(in[211]), .out(far_0_890_0[0]));    relay_conn far_0_890_0_b(.in(in[134]), .out(far_0_890_0[1]));
    wire [1:0] far_0_890_1;    relay_conn far_0_890_1_a(.in(far_0_890_0[0]), .out(far_0_890_1[0]));    relay_conn far_0_890_1_b(.in(far_0_890_0[1]), .out(far_0_890_1[1]));
    assign layer_0[890] = ~(far_0_890_1[0] & far_0_890_1[1]); 
    wire [1:0] far_0_891_0;    relay_conn far_0_891_0_a(.in(in[113]), .out(far_0_891_0[0]));    relay_conn far_0_891_0_b(.in(in[241]), .out(far_0_891_0[1]));
    wire [1:0] far_0_891_1;    relay_conn far_0_891_1_a(.in(far_0_891_0[0]), .out(far_0_891_1[0]));    relay_conn far_0_891_1_b(.in(far_0_891_0[1]), .out(far_0_891_1[1]));
    wire [1:0] far_0_891_2;    relay_conn far_0_891_2_a(.in(far_0_891_1[0]), .out(far_0_891_2[0]));    relay_conn far_0_891_2_b(.in(far_0_891_1[1]), .out(far_0_891_2[1]));
    wire [1:0] far_0_891_3;    relay_conn far_0_891_3_a(.in(far_0_891_2[0]), .out(far_0_891_3[0]));    relay_conn far_0_891_3_b(.in(far_0_891_2[1]), .out(far_0_891_3[1]));
    assign layer_0[891] = ~far_0_891_3[1]; 
    assign layer_0[892] = in[88] & ~in[91]; 
    wire [1:0] far_0_893_0;    relay_conn far_0_893_0_a(.in(in[136]), .out(far_0_893_0[0]));    relay_conn far_0_893_0_b(.in(in[19]), .out(far_0_893_0[1]));
    wire [1:0] far_0_893_1;    relay_conn far_0_893_1_a(.in(far_0_893_0[0]), .out(far_0_893_1[0]));    relay_conn far_0_893_1_b(.in(far_0_893_0[1]), .out(far_0_893_1[1]));
    wire [1:0] far_0_893_2;    relay_conn far_0_893_2_a(.in(far_0_893_1[0]), .out(far_0_893_2[0]));    relay_conn far_0_893_2_b(.in(far_0_893_1[1]), .out(far_0_893_2[1]));
    assign layer_0[893] = far_0_893_2[0] & ~far_0_893_2[1]; 
    assign layer_0[894] = ~in[22] | (in[19] & in[22]); 
    wire [1:0] far_0_895_0;    relay_conn far_0_895_0_a(.in(in[239]), .out(far_0_895_0[0]));    relay_conn far_0_895_0_b(.in(in[131]), .out(far_0_895_0[1]));
    wire [1:0] far_0_895_1;    relay_conn far_0_895_1_a(.in(far_0_895_0[0]), .out(far_0_895_1[0]));    relay_conn far_0_895_1_b(.in(far_0_895_0[1]), .out(far_0_895_1[1]));
    wire [1:0] far_0_895_2;    relay_conn far_0_895_2_a(.in(far_0_895_1[0]), .out(far_0_895_2[0]));    relay_conn far_0_895_2_b(.in(far_0_895_1[1]), .out(far_0_895_2[1]));
    assign layer_0[895] = ~far_0_895_2[0]; 
    wire [1:0] far_0_896_0;    relay_conn far_0_896_0_a(.in(in[165]), .out(far_0_896_0[0]));    relay_conn far_0_896_0_b(.in(in[72]), .out(far_0_896_0[1]));
    wire [1:0] far_0_896_1;    relay_conn far_0_896_1_a(.in(far_0_896_0[0]), .out(far_0_896_1[0]));    relay_conn far_0_896_1_b(.in(far_0_896_0[1]), .out(far_0_896_1[1]));
    assign layer_0[896] = far_0_896_1[1]; 
    assign layer_0[897] = ~(in[88] | in[84]); 
    wire [1:0] far_0_898_0;    relay_conn far_0_898_0_a(.in(in[173]), .out(far_0_898_0[0]));    relay_conn far_0_898_0_b(.in(in[88]), .out(far_0_898_0[1]));
    wire [1:0] far_0_898_1;    relay_conn far_0_898_1_a(.in(far_0_898_0[0]), .out(far_0_898_1[0]));    relay_conn far_0_898_1_b(.in(far_0_898_0[1]), .out(far_0_898_1[1]));
    assign layer_0[898] = far_0_898_1[0]; 
    assign layer_0[899] = ~(in[34] & in[6]); 
    wire [1:0] far_0_900_0;    relay_conn far_0_900_0_a(.in(in[74]), .out(far_0_900_0[0]));    relay_conn far_0_900_0_b(.in(in[116]), .out(far_0_900_0[1]));
    assign layer_0[900] = far_0_900_0[0] ^ far_0_900_0[1]; 
    wire [1:0] far_0_901_0;    relay_conn far_0_901_0_a(.in(in[228]), .out(far_0_901_0[0]));    relay_conn far_0_901_0_b(.in(in[151]), .out(far_0_901_0[1]));
    wire [1:0] far_0_901_1;    relay_conn far_0_901_1_a(.in(far_0_901_0[0]), .out(far_0_901_1[0]));    relay_conn far_0_901_1_b(.in(far_0_901_0[1]), .out(far_0_901_1[1]));
    assign layer_0[901] = far_0_901_1[1] & ~far_0_901_1[0]; 
    wire [1:0] far_0_902_0;    relay_conn far_0_902_0_a(.in(in[135]), .out(far_0_902_0[0]));    relay_conn far_0_902_0_b(.in(in[103]), .out(far_0_902_0[1]));
    assign layer_0[902] = far_0_902_0[0]; 
    assign layer_0[903] = in[254] & in[238]; 
    assign layer_0[904] = ~(in[199] ^ in[187]); 
    wire [1:0] far_0_905_0;    relay_conn far_0_905_0_a(.in(in[121]), .out(far_0_905_0[0]));    relay_conn far_0_905_0_b(.in(in[241]), .out(far_0_905_0[1]));
    wire [1:0] far_0_905_1;    relay_conn far_0_905_1_a(.in(far_0_905_0[0]), .out(far_0_905_1[0]));    relay_conn far_0_905_1_b(.in(far_0_905_0[1]), .out(far_0_905_1[1]));
    wire [1:0] far_0_905_2;    relay_conn far_0_905_2_a(.in(far_0_905_1[0]), .out(far_0_905_2[0]));    relay_conn far_0_905_2_b(.in(far_0_905_1[1]), .out(far_0_905_2[1]));
    assign layer_0[905] = far_0_905_2[1] & ~far_0_905_2[0]; 
    wire [1:0] far_0_906_0;    relay_conn far_0_906_0_a(.in(in[28]), .out(far_0_906_0[0]));    relay_conn far_0_906_0_b(.in(in[94]), .out(far_0_906_0[1]));
    wire [1:0] far_0_906_1;    relay_conn far_0_906_1_a(.in(far_0_906_0[0]), .out(far_0_906_1[0]));    relay_conn far_0_906_1_b(.in(far_0_906_0[1]), .out(far_0_906_1[1]));
    assign layer_0[906] = ~far_0_906_1[1] | (far_0_906_1[0] & far_0_906_1[1]); 
    wire [1:0] far_0_907_0;    relay_conn far_0_907_0_a(.in(in[56]), .out(far_0_907_0[0]));    relay_conn far_0_907_0_b(.in(in[165]), .out(far_0_907_0[1]));
    wire [1:0] far_0_907_1;    relay_conn far_0_907_1_a(.in(far_0_907_0[0]), .out(far_0_907_1[0]));    relay_conn far_0_907_1_b(.in(far_0_907_0[1]), .out(far_0_907_1[1]));
    wire [1:0] far_0_907_2;    relay_conn far_0_907_2_a(.in(far_0_907_1[0]), .out(far_0_907_2[0]));    relay_conn far_0_907_2_b(.in(far_0_907_1[1]), .out(far_0_907_2[1]));
    assign layer_0[907] = far_0_907_2[0] | far_0_907_2[1]; 
    wire [1:0] far_0_908_0;    relay_conn far_0_908_0_a(.in(in[197]), .out(far_0_908_0[0]));    relay_conn far_0_908_0_b(.in(in[236]), .out(far_0_908_0[1]));
    assign layer_0[908] = ~far_0_908_0[0]; 
    wire [1:0] far_0_909_0;    relay_conn far_0_909_0_a(.in(in[125]), .out(far_0_909_0[0]));    relay_conn far_0_909_0_b(.in(in[0]), .out(far_0_909_0[1]));
    wire [1:0] far_0_909_1;    relay_conn far_0_909_1_a(.in(far_0_909_0[0]), .out(far_0_909_1[0]));    relay_conn far_0_909_1_b(.in(far_0_909_0[1]), .out(far_0_909_1[1]));
    wire [1:0] far_0_909_2;    relay_conn far_0_909_2_a(.in(far_0_909_1[0]), .out(far_0_909_2[0]));    relay_conn far_0_909_2_b(.in(far_0_909_1[1]), .out(far_0_909_2[1]));
    assign layer_0[909] = ~far_0_909_2[0]; 
    assign layer_0[910] = ~(in[113] | in[98]); 
    wire [1:0] far_0_911_0;    relay_conn far_0_911_0_a(.in(in[79]), .out(far_0_911_0[0]));    relay_conn far_0_911_0_b(.in(in[207]), .out(far_0_911_0[1]));
    wire [1:0] far_0_911_1;    relay_conn far_0_911_1_a(.in(far_0_911_0[0]), .out(far_0_911_1[0]));    relay_conn far_0_911_1_b(.in(far_0_911_0[1]), .out(far_0_911_1[1]));
    wire [1:0] far_0_911_2;    relay_conn far_0_911_2_a(.in(far_0_911_1[0]), .out(far_0_911_2[0]));    relay_conn far_0_911_2_b(.in(far_0_911_1[1]), .out(far_0_911_2[1]));
    wire [1:0] far_0_911_3;    relay_conn far_0_911_3_a(.in(far_0_911_2[0]), .out(far_0_911_3[0]));    relay_conn far_0_911_3_b(.in(far_0_911_2[1]), .out(far_0_911_3[1]));
    assign layer_0[911] = ~(far_0_911_3[0] | far_0_911_3[1]); 
    wire [1:0] far_0_912_0;    relay_conn far_0_912_0_a(.in(in[116]), .out(far_0_912_0[0]));    relay_conn far_0_912_0_b(.in(in[168]), .out(far_0_912_0[1]));
    assign layer_0[912] = far_0_912_0[0] ^ far_0_912_0[1]; 
    wire [1:0] far_0_913_0;    relay_conn far_0_913_0_a(.in(in[73]), .out(far_0_913_0[0]));    relay_conn far_0_913_0_b(.in(in[164]), .out(far_0_913_0[1]));
    wire [1:0] far_0_913_1;    relay_conn far_0_913_1_a(.in(far_0_913_0[0]), .out(far_0_913_1[0]));    relay_conn far_0_913_1_b(.in(far_0_913_0[1]), .out(far_0_913_1[1]));
    assign layer_0[913] = ~far_0_913_1[0] | (far_0_913_1[0] & far_0_913_1[1]); 
    assign layer_0[914] = in[137]; 
    wire [1:0] far_0_915_0;    relay_conn far_0_915_0_a(.in(in[104]), .out(far_0_915_0[0]));    relay_conn far_0_915_0_b(.in(in[8]), .out(far_0_915_0[1]));
    wire [1:0] far_0_915_1;    relay_conn far_0_915_1_a(.in(far_0_915_0[0]), .out(far_0_915_1[0]));    relay_conn far_0_915_1_b(.in(far_0_915_0[1]), .out(far_0_915_1[1]));
    wire [1:0] far_0_915_2;    relay_conn far_0_915_2_a(.in(far_0_915_1[0]), .out(far_0_915_2[0]));    relay_conn far_0_915_2_b(.in(far_0_915_1[1]), .out(far_0_915_2[1]));
    assign layer_0[915] = far_0_915_2[1]; 
    wire [1:0] far_0_916_0;    relay_conn far_0_916_0_a(.in(in[119]), .out(far_0_916_0[0]));    relay_conn far_0_916_0_b(.in(in[199]), .out(far_0_916_0[1]));
    wire [1:0] far_0_916_1;    relay_conn far_0_916_1_a(.in(far_0_916_0[0]), .out(far_0_916_1[0]));    relay_conn far_0_916_1_b(.in(far_0_916_0[1]), .out(far_0_916_1[1]));
    assign layer_0[916] = ~(far_0_916_1[0] | far_0_916_1[1]); 
    assign layer_0[917] = ~in[27]; 
    wire [1:0] far_0_918_0;    relay_conn far_0_918_0_a(.in(in[215]), .out(far_0_918_0[0]));    relay_conn far_0_918_0_b(.in(in[150]), .out(far_0_918_0[1]));
    wire [1:0] far_0_918_1;    relay_conn far_0_918_1_a(.in(far_0_918_0[0]), .out(far_0_918_1[0]));    relay_conn far_0_918_1_b(.in(far_0_918_0[1]), .out(far_0_918_1[1]));
    assign layer_0[918] = ~(far_0_918_1[0] & far_0_918_1[1]); 
    wire [1:0] far_0_919_0;    relay_conn far_0_919_0_a(.in(in[181]), .out(far_0_919_0[0]));    relay_conn far_0_919_0_b(.in(in[237]), .out(far_0_919_0[1]));
    assign layer_0[919] = ~far_0_919_0[0] | (far_0_919_0[0] & far_0_919_0[1]); 
    assign layer_0[920] = in[199] & ~in[203]; 
    wire [1:0] far_0_921_0;    relay_conn far_0_921_0_a(.in(in[175]), .out(far_0_921_0[0]));    relay_conn far_0_921_0_b(.in(in[134]), .out(far_0_921_0[1]));
    assign layer_0[921] = far_0_921_0[0] | far_0_921_0[1]; 
    assign layer_0[922] = in[164]; 
    wire [1:0] far_0_923_0;    relay_conn far_0_923_0_a(.in(in[241]), .out(far_0_923_0[0]));    relay_conn far_0_923_0_b(.in(in[170]), .out(far_0_923_0[1]));
    wire [1:0] far_0_923_1;    relay_conn far_0_923_1_a(.in(far_0_923_0[0]), .out(far_0_923_1[0]));    relay_conn far_0_923_1_b(.in(far_0_923_0[1]), .out(far_0_923_1[1]));
    assign layer_0[923] = far_0_923_1[0] & far_0_923_1[1]; 
    wire [1:0] far_0_924_0;    relay_conn far_0_924_0_a(.in(in[197]), .out(far_0_924_0[0]));    relay_conn far_0_924_0_b(.in(in[117]), .out(far_0_924_0[1]));
    wire [1:0] far_0_924_1;    relay_conn far_0_924_1_a(.in(far_0_924_0[0]), .out(far_0_924_1[0]));    relay_conn far_0_924_1_b(.in(far_0_924_0[1]), .out(far_0_924_1[1]));
    assign layer_0[924] = far_0_924_1[0] | far_0_924_1[1]; 
    wire [1:0] far_0_925_0;    relay_conn far_0_925_0_a(.in(in[190]), .out(far_0_925_0[0]));    relay_conn far_0_925_0_b(.in(in[71]), .out(far_0_925_0[1]));
    wire [1:0] far_0_925_1;    relay_conn far_0_925_1_a(.in(far_0_925_0[0]), .out(far_0_925_1[0]));    relay_conn far_0_925_1_b(.in(far_0_925_0[1]), .out(far_0_925_1[1]));
    wire [1:0] far_0_925_2;    relay_conn far_0_925_2_a(.in(far_0_925_1[0]), .out(far_0_925_2[0]));    relay_conn far_0_925_2_b(.in(far_0_925_1[1]), .out(far_0_925_2[1]));
    assign layer_0[925] = ~far_0_925_2[0] | (far_0_925_2[0] & far_0_925_2[1]); 
    wire [1:0] far_0_926_0;    relay_conn far_0_926_0_a(.in(in[93]), .out(far_0_926_0[0]));    relay_conn far_0_926_0_b(.in(in[181]), .out(far_0_926_0[1]));
    wire [1:0] far_0_926_1;    relay_conn far_0_926_1_a(.in(far_0_926_0[0]), .out(far_0_926_1[0]));    relay_conn far_0_926_1_b(.in(far_0_926_0[1]), .out(far_0_926_1[1]));
    assign layer_0[926] = far_0_926_1[0] | far_0_926_1[1]; 
    wire [1:0] far_0_927_0;    relay_conn far_0_927_0_a(.in(in[211]), .out(far_0_927_0[0]));    relay_conn far_0_927_0_b(.in(in[157]), .out(far_0_927_0[1]));
    assign layer_0[927] = ~(far_0_927_0[0] | far_0_927_0[1]); 
    assign layer_0[928] = in[186] & in[202]; 
    wire [1:0] far_0_929_0;    relay_conn far_0_929_0_a(.in(in[48]), .out(far_0_929_0[0]));    relay_conn far_0_929_0_b(.in(in[158]), .out(far_0_929_0[1]));
    wire [1:0] far_0_929_1;    relay_conn far_0_929_1_a(.in(far_0_929_0[0]), .out(far_0_929_1[0]));    relay_conn far_0_929_1_b(.in(far_0_929_0[1]), .out(far_0_929_1[1]));
    wire [1:0] far_0_929_2;    relay_conn far_0_929_2_a(.in(far_0_929_1[0]), .out(far_0_929_2[0]));    relay_conn far_0_929_2_b(.in(far_0_929_1[1]), .out(far_0_929_2[1]));
    assign layer_0[929] = far_0_929_2[0] | far_0_929_2[1]; 
    wire [1:0] far_0_930_0;    relay_conn far_0_930_0_a(.in(in[70]), .out(far_0_930_0[0]));    relay_conn far_0_930_0_b(.in(in[117]), .out(far_0_930_0[1]));
    assign layer_0[930] = ~far_0_930_0[0] | (far_0_930_0[0] & far_0_930_0[1]); 
    assign layer_0[931] = in[207] & in[186]; 
    wire [1:0] far_0_932_0;    relay_conn far_0_932_0_a(.in(in[199]), .out(far_0_932_0[0]));    relay_conn far_0_932_0_b(.in(in[132]), .out(far_0_932_0[1]));
    wire [1:0] far_0_932_1;    relay_conn far_0_932_1_a(.in(far_0_932_0[0]), .out(far_0_932_1[0]));    relay_conn far_0_932_1_b(.in(far_0_932_0[1]), .out(far_0_932_1[1]));
    assign layer_0[932] = far_0_932_1[0] & ~far_0_932_1[1]; 
    assign layer_0[933] = ~(in[207] & in[199]); 
    wire [1:0] far_0_934_0;    relay_conn far_0_934_0_a(.in(in[215]), .out(far_0_934_0[0]));    relay_conn far_0_934_0_b(.in(in[125]), .out(far_0_934_0[1]));
    wire [1:0] far_0_934_1;    relay_conn far_0_934_1_a(.in(far_0_934_0[0]), .out(far_0_934_1[0]));    relay_conn far_0_934_1_b(.in(far_0_934_0[1]), .out(far_0_934_1[1]));
    assign layer_0[934] = far_0_934_1[0] ^ far_0_934_1[1]; 
    wire [1:0] far_0_935_0;    relay_conn far_0_935_0_a(.in(in[22]), .out(far_0_935_0[0]));    relay_conn far_0_935_0_b(.in(in[142]), .out(far_0_935_0[1]));
    wire [1:0] far_0_935_1;    relay_conn far_0_935_1_a(.in(far_0_935_0[0]), .out(far_0_935_1[0]));    relay_conn far_0_935_1_b(.in(far_0_935_0[1]), .out(far_0_935_1[1]));
    wire [1:0] far_0_935_2;    relay_conn far_0_935_2_a(.in(far_0_935_1[0]), .out(far_0_935_2[0]));    relay_conn far_0_935_2_b(.in(far_0_935_1[1]), .out(far_0_935_2[1]));
    assign layer_0[935] = far_0_935_2[0] | far_0_935_2[1]; 
    assign layer_0[936] = ~(in[130] & in[133]); 
    wire [1:0] far_0_937_0;    relay_conn far_0_937_0_a(.in(in[239]), .out(far_0_937_0[0]));    relay_conn far_0_937_0_b(.in(in[139]), .out(far_0_937_0[1]));
    wire [1:0] far_0_937_1;    relay_conn far_0_937_1_a(.in(far_0_937_0[0]), .out(far_0_937_1[0]));    relay_conn far_0_937_1_b(.in(far_0_937_0[1]), .out(far_0_937_1[1]));
    wire [1:0] far_0_937_2;    relay_conn far_0_937_2_a(.in(far_0_937_1[0]), .out(far_0_937_2[0]));    relay_conn far_0_937_2_b(.in(far_0_937_1[1]), .out(far_0_937_2[1]));
    assign layer_0[937] = ~(far_0_937_2[0] & far_0_937_2[1]); 
    wire [1:0] far_0_938_0;    relay_conn far_0_938_0_a(.in(in[147]), .out(far_0_938_0[0]));    relay_conn far_0_938_0_b(.in(in[113]), .out(far_0_938_0[1]));
    assign layer_0[938] = far_0_938_0[1] & ~far_0_938_0[0]; 
    assign layer_0[939] = ~in[174]; 
    wire [1:0] far_0_940_0;    relay_conn far_0_940_0_a(.in(in[172]), .out(far_0_940_0[0]));    relay_conn far_0_940_0_b(.in(in[133]), .out(far_0_940_0[1]));
    assign layer_0[940] = far_0_940_0[0] & ~far_0_940_0[1]; 
    assign layer_0[941] = ~in[114]; 
    assign layer_0[942] = ~(in[93] | in[90]); 
    wire [1:0] far_0_943_0;    relay_conn far_0_943_0_a(.in(in[221]), .out(far_0_943_0[0]));    relay_conn far_0_943_0_b(.in(in[125]), .out(far_0_943_0[1]));
    wire [1:0] far_0_943_1;    relay_conn far_0_943_1_a(.in(far_0_943_0[0]), .out(far_0_943_1[0]));    relay_conn far_0_943_1_b(.in(far_0_943_0[1]), .out(far_0_943_1[1]));
    wire [1:0] far_0_943_2;    relay_conn far_0_943_2_a(.in(far_0_943_1[0]), .out(far_0_943_2[0]));    relay_conn far_0_943_2_b(.in(far_0_943_1[1]), .out(far_0_943_2[1]));
    assign layer_0[943] = far_0_943_2[1]; 
    wire [1:0] far_0_944_0;    relay_conn far_0_944_0_a(.in(in[154]), .out(far_0_944_0[0]));    relay_conn far_0_944_0_b(.in(in[66]), .out(far_0_944_0[1]));
    wire [1:0] far_0_944_1;    relay_conn far_0_944_1_a(.in(far_0_944_0[0]), .out(far_0_944_1[0]));    relay_conn far_0_944_1_b(.in(far_0_944_0[1]), .out(far_0_944_1[1]));
    assign layer_0[944] = ~far_0_944_1[0]; 
    wire [1:0] far_0_945_0;    relay_conn far_0_945_0_a(.in(in[101]), .out(far_0_945_0[0]));    relay_conn far_0_945_0_b(.in(in[181]), .out(far_0_945_0[1]));
    wire [1:0] far_0_945_1;    relay_conn far_0_945_1_a(.in(far_0_945_0[0]), .out(far_0_945_1[0]));    relay_conn far_0_945_1_b(.in(far_0_945_0[1]), .out(far_0_945_1[1]));
    assign layer_0[945] = far_0_945_1[0] & far_0_945_1[1]; 
    wire [1:0] far_0_946_0;    relay_conn far_0_946_0_a(.in(in[122]), .out(far_0_946_0[0]));    relay_conn far_0_946_0_b(.in(in[215]), .out(far_0_946_0[1]));
    wire [1:0] far_0_946_1;    relay_conn far_0_946_1_a(.in(far_0_946_0[0]), .out(far_0_946_1[0]));    relay_conn far_0_946_1_b(.in(far_0_946_0[1]), .out(far_0_946_1[1]));
    assign layer_0[946] = ~far_0_946_1[0] | (far_0_946_1[0] & far_0_946_1[1]); 
    wire [1:0] far_0_947_0;    relay_conn far_0_947_0_a(.in(in[190]), .out(far_0_947_0[0]));    relay_conn far_0_947_0_b(.in(in[142]), .out(far_0_947_0[1]));
    assign layer_0[947] = far_0_947_0[1] & ~far_0_947_0[0]; 
    wire [1:0] far_0_948_0;    relay_conn far_0_948_0_a(.in(in[205]), .out(far_0_948_0[0]));    relay_conn far_0_948_0_b(.in(in[143]), .out(far_0_948_0[1]));
    assign layer_0[948] = ~far_0_948_0[0] | (far_0_948_0[0] & far_0_948_0[1]); 
    wire [1:0] far_0_949_0;    relay_conn far_0_949_0_a(.in(in[136]), .out(far_0_949_0[0]));    relay_conn far_0_949_0_b(.in(in[222]), .out(far_0_949_0[1]));
    wire [1:0] far_0_949_1;    relay_conn far_0_949_1_a(.in(far_0_949_0[0]), .out(far_0_949_1[0]));    relay_conn far_0_949_1_b(.in(far_0_949_0[1]), .out(far_0_949_1[1]));
    assign layer_0[949] = ~far_0_949_1[1]; 
    wire [1:0] far_0_950_0;    relay_conn far_0_950_0_a(.in(in[132]), .out(far_0_950_0[0]));    relay_conn far_0_950_0_b(.in(in[202]), .out(far_0_950_0[1]));
    wire [1:0] far_0_950_1;    relay_conn far_0_950_1_a(.in(far_0_950_0[0]), .out(far_0_950_1[0]));    relay_conn far_0_950_1_b(.in(far_0_950_0[1]), .out(far_0_950_1[1]));
    assign layer_0[950] = far_0_950_1[0]; 
    assign layer_0[951] = ~in[19] | (in[0] & in[19]); 
    wire [1:0] far_0_952_0;    relay_conn far_0_952_0_a(.in(in[66]), .out(far_0_952_0[0]));    relay_conn far_0_952_0_b(.in(in[157]), .out(far_0_952_0[1]));
    wire [1:0] far_0_952_1;    relay_conn far_0_952_1_a(.in(far_0_952_0[0]), .out(far_0_952_1[0]));    relay_conn far_0_952_1_b(.in(far_0_952_0[1]), .out(far_0_952_1[1]));
    assign layer_0[952] = far_0_952_1[0] & far_0_952_1[1]; 
    wire [1:0] far_0_953_0;    relay_conn far_0_953_0_a(.in(in[149]), .out(far_0_953_0[0]));    relay_conn far_0_953_0_b(.in(in[48]), .out(far_0_953_0[1]));
    wire [1:0] far_0_953_1;    relay_conn far_0_953_1_a(.in(far_0_953_0[0]), .out(far_0_953_1[0]));    relay_conn far_0_953_1_b(.in(far_0_953_0[1]), .out(far_0_953_1[1]));
    wire [1:0] far_0_953_2;    relay_conn far_0_953_2_a(.in(far_0_953_1[0]), .out(far_0_953_2[0]));    relay_conn far_0_953_2_b(.in(far_0_953_1[1]), .out(far_0_953_2[1]));
    assign layer_0[953] = ~far_0_953_2[0] | (far_0_953_2[0] & far_0_953_2[1]); 
    assign layer_0[954] = in[132]; 
    assign layer_0[955] = ~(in[63] | in[78]); 
    assign layer_0[956] = in[154]; 
    assign layer_0[957] = in[111]; 
    wire [1:0] far_0_958_0;    relay_conn far_0_958_0_a(.in(in[215]), .out(far_0_958_0[0]));    relay_conn far_0_958_0_b(.in(in[132]), .out(far_0_958_0[1]));
    wire [1:0] far_0_958_1;    relay_conn far_0_958_1_a(.in(far_0_958_0[0]), .out(far_0_958_1[0]));    relay_conn far_0_958_1_b(.in(far_0_958_0[1]), .out(far_0_958_1[1]));
    assign layer_0[958] = far_0_958_1[0]; 
    wire [1:0] far_0_959_0;    relay_conn far_0_959_0_a(.in(in[125]), .out(far_0_959_0[0]));    relay_conn far_0_959_0_b(.in(in[63]), .out(far_0_959_0[1]));
    assign layer_0[959] = ~(far_0_959_0[0] & far_0_959_0[1]); 
    wire [1:0] far_0_960_0;    relay_conn far_0_960_0_a(.in(in[99]), .out(far_0_960_0[0]));    relay_conn far_0_960_0_b(.in(in[48]), .out(far_0_960_0[1]));
    assign layer_0[960] = ~(far_0_960_0[0] & far_0_960_0[1]); 
    wire [1:0] far_0_961_0;    relay_conn far_0_961_0_a(.in(in[19]), .out(far_0_961_0[0]));    relay_conn far_0_961_0_b(.in(in[133]), .out(far_0_961_0[1]));
    wire [1:0] far_0_961_1;    relay_conn far_0_961_1_a(.in(far_0_961_0[0]), .out(far_0_961_1[0]));    relay_conn far_0_961_1_b(.in(far_0_961_0[1]), .out(far_0_961_1[1]));
    wire [1:0] far_0_961_2;    relay_conn far_0_961_2_a(.in(far_0_961_1[0]), .out(far_0_961_2[0]));    relay_conn far_0_961_2_b(.in(far_0_961_1[1]), .out(far_0_961_2[1]));
    assign layer_0[961] = far_0_961_2[0] & far_0_961_2[1]; 
    wire [1:0] far_0_962_0;    relay_conn far_0_962_0_a(.in(in[13]), .out(far_0_962_0[0]));    relay_conn far_0_962_0_b(.in(in[80]), .out(far_0_962_0[1]));
    wire [1:0] far_0_962_1;    relay_conn far_0_962_1_a(.in(far_0_962_0[0]), .out(far_0_962_1[0]));    relay_conn far_0_962_1_b(.in(far_0_962_0[1]), .out(far_0_962_1[1]));
    assign layer_0[962] = far_0_962_1[0] | far_0_962_1[1]; 
    wire [1:0] far_0_963_0;    relay_conn far_0_963_0_a(.in(in[17]), .out(far_0_963_0[0]));    relay_conn far_0_963_0_b(.in(in[57]), .out(far_0_963_0[1]));
    assign layer_0[963] = ~(far_0_963_0[0] | far_0_963_0[1]); 
    assign layer_0[964] = ~in[215]; 
    wire [1:0] far_0_965_0;    relay_conn far_0_965_0_a(.in(in[24]), .out(far_0_965_0[0]));    relay_conn far_0_965_0_b(.in(in[93]), .out(far_0_965_0[1]));
    wire [1:0] far_0_965_1;    relay_conn far_0_965_1_a(.in(far_0_965_0[0]), .out(far_0_965_1[0]));    relay_conn far_0_965_1_b(.in(far_0_965_0[1]), .out(far_0_965_1[1]));
    assign layer_0[965] = ~(far_0_965_1[0] | far_0_965_1[1]); 
    wire [1:0] far_0_966_0;    relay_conn far_0_966_0_a(.in(in[141]), .out(far_0_966_0[0]));    relay_conn far_0_966_0_b(.in(in[212]), .out(far_0_966_0[1]));
    wire [1:0] far_0_966_1;    relay_conn far_0_966_1_a(.in(far_0_966_0[0]), .out(far_0_966_1[0]));    relay_conn far_0_966_1_b(.in(far_0_966_0[1]), .out(far_0_966_1[1]));
    assign layer_0[966] = far_0_966_1[0] | far_0_966_1[1]; 
    assign layer_0[967] = in[104] & ~in[113]; 
    wire [1:0] far_0_968_0;    relay_conn far_0_968_0_a(.in(in[113]), .out(far_0_968_0[0]));    relay_conn far_0_968_0_b(.in(in[210]), .out(far_0_968_0[1]));
    wire [1:0] far_0_968_1;    relay_conn far_0_968_1_a(.in(far_0_968_0[0]), .out(far_0_968_1[0]));    relay_conn far_0_968_1_b(.in(far_0_968_0[1]), .out(far_0_968_1[1]));
    wire [1:0] far_0_968_2;    relay_conn far_0_968_2_a(.in(far_0_968_1[0]), .out(far_0_968_2[0]));    relay_conn far_0_968_2_b(.in(far_0_968_1[1]), .out(far_0_968_2[1]));
    assign layer_0[968] = far_0_968_2[0]; 
    assign layer_0[969] = ~in[219] | (in[198] & in[219]); 
    wire [1:0] far_0_970_0;    relay_conn far_0_970_0_a(.in(in[43]), .out(far_0_970_0[0]));    relay_conn far_0_970_0_b(.in(in[111]), .out(far_0_970_0[1]));
    wire [1:0] far_0_970_1;    relay_conn far_0_970_1_a(.in(far_0_970_0[0]), .out(far_0_970_1[0]));    relay_conn far_0_970_1_b(.in(far_0_970_0[1]), .out(far_0_970_1[1]));
    assign layer_0[970] = far_0_970_1[1]; 
    wire [1:0] far_0_971_0;    relay_conn far_0_971_0_a(.in(in[79]), .out(far_0_971_0[0]));    relay_conn far_0_971_0_b(.in(in[179]), .out(far_0_971_0[1]));
    wire [1:0] far_0_971_1;    relay_conn far_0_971_1_a(.in(far_0_971_0[0]), .out(far_0_971_1[0]));    relay_conn far_0_971_1_b(.in(far_0_971_0[1]), .out(far_0_971_1[1]));
    wire [1:0] far_0_971_2;    relay_conn far_0_971_2_a(.in(far_0_971_1[0]), .out(far_0_971_2[0]));    relay_conn far_0_971_2_b(.in(far_0_971_1[1]), .out(far_0_971_2[1]));
    assign layer_0[971] = ~far_0_971_2[0]; 
    assign layer_0[972] = ~in[90]; 
    wire [1:0] far_0_973_0;    relay_conn far_0_973_0_a(.in(in[150]), .out(far_0_973_0[0]));    relay_conn far_0_973_0_b(.in(in[49]), .out(far_0_973_0[1]));
    wire [1:0] far_0_973_1;    relay_conn far_0_973_1_a(.in(far_0_973_0[0]), .out(far_0_973_1[0]));    relay_conn far_0_973_1_b(.in(far_0_973_0[1]), .out(far_0_973_1[1]));
    wire [1:0] far_0_973_2;    relay_conn far_0_973_2_a(.in(far_0_973_1[0]), .out(far_0_973_2[0]));    relay_conn far_0_973_2_b(.in(far_0_973_1[1]), .out(far_0_973_2[1]));
    assign layer_0[973] = ~far_0_973_2[0]; 
    wire [1:0] far_0_974_0;    relay_conn far_0_974_0_a(.in(in[44]), .out(far_0_974_0[0]));    relay_conn far_0_974_0_b(.in(in[142]), .out(far_0_974_0[1]));
    wire [1:0] far_0_974_1;    relay_conn far_0_974_1_a(.in(far_0_974_0[0]), .out(far_0_974_1[0]));    relay_conn far_0_974_1_b(.in(far_0_974_0[1]), .out(far_0_974_1[1]));
    wire [1:0] far_0_974_2;    relay_conn far_0_974_2_a(.in(far_0_974_1[0]), .out(far_0_974_2[0]));    relay_conn far_0_974_2_b(.in(far_0_974_1[1]), .out(far_0_974_2[1]));
    assign layer_0[974] = ~(far_0_974_2[0] & far_0_974_2[1]); 
    wire [1:0] far_0_975_0;    relay_conn far_0_975_0_a(.in(in[170]), .out(far_0_975_0[0]));    relay_conn far_0_975_0_b(.in(in[113]), .out(far_0_975_0[1]));
    assign layer_0[975] = far_0_975_0[0] ^ far_0_975_0[1]; 
    wire [1:0] far_0_976_0;    relay_conn far_0_976_0_a(.in(in[158]), .out(far_0_976_0[0]));    relay_conn far_0_976_0_b(.in(in[205]), .out(far_0_976_0[1]));
    assign layer_0[976] = far_0_976_0[0] & far_0_976_0[1]; 
    wire [1:0] far_0_977_0;    relay_conn far_0_977_0_a(.in(in[150]), .out(far_0_977_0[0]));    relay_conn far_0_977_0_b(.in(in[41]), .out(far_0_977_0[1]));
    wire [1:0] far_0_977_1;    relay_conn far_0_977_1_a(.in(far_0_977_0[0]), .out(far_0_977_1[0]));    relay_conn far_0_977_1_b(.in(far_0_977_0[1]), .out(far_0_977_1[1]));
    wire [1:0] far_0_977_2;    relay_conn far_0_977_2_a(.in(far_0_977_1[0]), .out(far_0_977_2[0]));    relay_conn far_0_977_2_b(.in(far_0_977_1[1]), .out(far_0_977_2[1]));
    assign layer_0[977] = far_0_977_2[0]; 
    assign layer_0[978] = in[31]; 
    assign layer_0[979] = ~(in[125] | in[132]); 
    wire [1:0] far_0_980_0;    relay_conn far_0_980_0_a(.in(in[136]), .out(far_0_980_0[0]));    relay_conn far_0_980_0_b(.in(in[233]), .out(far_0_980_0[1]));
    wire [1:0] far_0_980_1;    relay_conn far_0_980_1_a(.in(far_0_980_0[0]), .out(far_0_980_1[0]));    relay_conn far_0_980_1_b(.in(far_0_980_0[1]), .out(far_0_980_1[1]));
    wire [1:0] far_0_980_2;    relay_conn far_0_980_2_a(.in(far_0_980_1[0]), .out(far_0_980_2[0]));    relay_conn far_0_980_2_b(.in(far_0_980_1[1]), .out(far_0_980_2[1]));
    assign layer_0[980] = ~(far_0_980_2[0] & far_0_980_2[1]); 
    assign layer_0[981] = in[99]; 
    wire [1:0] far_0_982_0;    relay_conn far_0_982_0_a(.in(in[151]), .out(far_0_982_0[0]));    relay_conn far_0_982_0_b(.in(in[207]), .out(far_0_982_0[1]));
    assign layer_0[982] = far_0_982_0[1] & ~far_0_982_0[0]; 
    wire [1:0] far_0_983_0;    relay_conn far_0_983_0_a(.in(in[73]), .out(far_0_983_0[0]));    relay_conn far_0_983_0_b(.in(in[199]), .out(far_0_983_0[1]));
    wire [1:0] far_0_983_1;    relay_conn far_0_983_1_a(.in(far_0_983_0[0]), .out(far_0_983_1[0]));    relay_conn far_0_983_1_b(.in(far_0_983_0[1]), .out(far_0_983_1[1]));
    wire [1:0] far_0_983_2;    relay_conn far_0_983_2_a(.in(far_0_983_1[0]), .out(far_0_983_2[0]));    relay_conn far_0_983_2_b(.in(far_0_983_1[1]), .out(far_0_983_2[1]));
    assign layer_0[983] = ~(far_0_983_2[0] & far_0_983_2[1]); 
    wire [1:0] far_0_984_0;    relay_conn far_0_984_0_a(.in(in[92]), .out(far_0_984_0[0]));    relay_conn far_0_984_0_b(.in(in[215]), .out(far_0_984_0[1]));
    wire [1:0] far_0_984_1;    relay_conn far_0_984_1_a(.in(far_0_984_0[0]), .out(far_0_984_1[0]));    relay_conn far_0_984_1_b(.in(far_0_984_0[1]), .out(far_0_984_1[1]));
    wire [1:0] far_0_984_2;    relay_conn far_0_984_2_a(.in(far_0_984_1[0]), .out(far_0_984_2[0]));    relay_conn far_0_984_2_b(.in(far_0_984_1[1]), .out(far_0_984_2[1]));
    assign layer_0[984] = far_0_984_2[0] & far_0_984_2[1]; 
    assign layer_0[985] = ~(in[174] | in[165]); 
    wire [1:0] far_0_986_0;    relay_conn far_0_986_0_a(.in(in[121]), .out(far_0_986_0[0]));    relay_conn far_0_986_0_b(.in(in[232]), .out(far_0_986_0[1]));
    wire [1:0] far_0_986_1;    relay_conn far_0_986_1_a(.in(far_0_986_0[0]), .out(far_0_986_1[0]));    relay_conn far_0_986_1_b(.in(far_0_986_0[1]), .out(far_0_986_1[1]));
    wire [1:0] far_0_986_2;    relay_conn far_0_986_2_a(.in(far_0_986_1[0]), .out(far_0_986_2[0]));    relay_conn far_0_986_2_b(.in(far_0_986_1[1]), .out(far_0_986_2[1]));
    assign layer_0[986] = ~far_0_986_2[0]; 
    wire [1:0] far_0_987_0;    relay_conn far_0_987_0_a(.in(in[247]), .out(far_0_987_0[0]));    relay_conn far_0_987_0_b(.in(in[188]), .out(far_0_987_0[1]));
    assign layer_0[987] = ~far_0_987_0[1]; 
    wire [1:0] far_0_988_0;    relay_conn far_0_988_0_a(.in(in[199]), .out(far_0_988_0[0]));    relay_conn far_0_988_0_b(.in(in[121]), .out(far_0_988_0[1]));
    wire [1:0] far_0_988_1;    relay_conn far_0_988_1_a(.in(far_0_988_0[0]), .out(far_0_988_1[0]));    relay_conn far_0_988_1_b(.in(far_0_988_0[1]), .out(far_0_988_1[1]));
    assign layer_0[988] = far_0_988_1[0]; 
    wire [1:0] far_0_989_0;    relay_conn far_0_989_0_a(.in(in[130]), .out(far_0_989_0[0]));    relay_conn far_0_989_0_b(.in(in[18]), .out(far_0_989_0[1]));
    wire [1:0] far_0_989_1;    relay_conn far_0_989_1_a(.in(far_0_989_0[0]), .out(far_0_989_1[0]));    relay_conn far_0_989_1_b(.in(far_0_989_0[1]), .out(far_0_989_1[1]));
    wire [1:0] far_0_989_2;    relay_conn far_0_989_2_a(.in(far_0_989_1[0]), .out(far_0_989_2[0]));    relay_conn far_0_989_2_b(.in(far_0_989_1[1]), .out(far_0_989_2[1]));
    assign layer_0[989] = ~far_0_989_2[1] | (far_0_989_2[0] & far_0_989_2[1]); 
    assign layer_0[990] = ~in[82] | (in[104] & in[82]); 
    assign layer_0[991] = in[193] & ~in[211]; 
    wire [1:0] far_0_992_0;    relay_conn far_0_992_0_a(.in(in[87]), .out(far_0_992_0[0]));    relay_conn far_0_992_0_b(.in(in[52]), .out(far_0_992_0[1]));
    assign layer_0[992] = ~far_0_992_0[0]; 
    assign layer_0[993] = in[212] & ~in[233]; 
    assign layer_0[994] = in[147]; 
    wire [1:0] far_0_995_0;    relay_conn far_0_995_0_a(.in(in[101]), .out(far_0_995_0[0]));    relay_conn far_0_995_0_b(.in(in[189]), .out(far_0_995_0[1]));
    wire [1:0] far_0_995_1;    relay_conn far_0_995_1_a(.in(far_0_995_0[0]), .out(far_0_995_1[0]));    relay_conn far_0_995_1_b(.in(far_0_995_0[1]), .out(far_0_995_1[1]));
    assign layer_0[995] = ~far_0_995_1[0]; 
    wire [1:0] far_0_996_0;    relay_conn far_0_996_0_a(.in(in[133]), .out(far_0_996_0[0]));    relay_conn far_0_996_0_b(.in(in[238]), .out(far_0_996_0[1]));
    wire [1:0] far_0_996_1;    relay_conn far_0_996_1_a(.in(far_0_996_0[0]), .out(far_0_996_1[0]));    relay_conn far_0_996_1_b(.in(far_0_996_0[1]), .out(far_0_996_1[1]));
    wire [1:0] far_0_996_2;    relay_conn far_0_996_2_a(.in(far_0_996_1[0]), .out(far_0_996_2[0]));    relay_conn far_0_996_2_b(.in(far_0_996_1[1]), .out(far_0_996_2[1]));
    assign layer_0[996] = far_0_996_2[0] | far_0_996_2[1]; 
    wire [1:0] far_0_997_0;    relay_conn far_0_997_0_a(.in(in[255]), .out(far_0_997_0[0]));    relay_conn far_0_997_0_b(.in(in[165]), .out(far_0_997_0[1]));
    wire [1:0] far_0_997_1;    relay_conn far_0_997_1_a(.in(far_0_997_0[0]), .out(far_0_997_1[0]));    relay_conn far_0_997_1_b(.in(far_0_997_0[1]), .out(far_0_997_1[1]));
    assign layer_0[997] = far_0_997_1[0] | far_0_997_1[1]; 
    wire [1:0] far_0_998_0;    relay_conn far_0_998_0_a(.in(in[3]), .out(far_0_998_0[0]));    relay_conn far_0_998_0_b(.in(in[93]), .out(far_0_998_0[1]));
    wire [1:0] far_0_998_1;    relay_conn far_0_998_1_a(.in(far_0_998_0[0]), .out(far_0_998_1[0]));    relay_conn far_0_998_1_b(.in(far_0_998_0[1]), .out(far_0_998_1[1]));
    assign layer_0[998] = far_0_998_1[0] & far_0_998_1[1]; 
    wire [1:0] far_0_999_0;    relay_conn far_0_999_0_a(.in(in[197]), .out(far_0_999_0[0]));    relay_conn far_0_999_0_b(.in(in[151]), .out(far_0_999_0[1]));
    assign layer_0[999] = ~far_0_999_0[1] | (far_0_999_0[0] & far_0_999_0[1]); 
    wire [1:0] far_0_1000_0;    relay_conn far_0_1000_0_a(.in(in[186]), .out(far_0_1000_0[0]));    relay_conn far_0_1000_0_b(.in(in[75]), .out(far_0_1000_0[1]));
    wire [1:0] far_0_1000_1;    relay_conn far_0_1000_1_a(.in(far_0_1000_0[0]), .out(far_0_1000_1[0]));    relay_conn far_0_1000_1_b(.in(far_0_1000_0[1]), .out(far_0_1000_1[1]));
    wire [1:0] far_0_1000_2;    relay_conn far_0_1000_2_a(.in(far_0_1000_1[0]), .out(far_0_1000_2[0]));    relay_conn far_0_1000_2_b(.in(far_0_1000_1[1]), .out(far_0_1000_2[1]));
    assign layer_0[1000] = ~far_0_1000_2[1]; 
    wire [1:0] far_0_1001_0;    relay_conn far_0_1001_0_a(.in(in[151]), .out(far_0_1001_0[0]));    relay_conn far_0_1001_0_b(.in(in[116]), .out(far_0_1001_0[1]));
    assign layer_0[1001] = far_0_1001_0[1] & ~far_0_1001_0[0]; 
    assign layer_0[1002] = ~in[44] | (in[44] & in[56]); 
    wire [1:0] far_0_1003_0;    relay_conn far_0_1003_0_a(.in(in[185]), .out(far_0_1003_0[0]));    relay_conn far_0_1003_0_b(.in(in[79]), .out(far_0_1003_0[1]));
    wire [1:0] far_0_1003_1;    relay_conn far_0_1003_1_a(.in(far_0_1003_0[0]), .out(far_0_1003_1[0]));    relay_conn far_0_1003_1_b(.in(far_0_1003_0[1]), .out(far_0_1003_1[1]));
    wire [1:0] far_0_1003_2;    relay_conn far_0_1003_2_a(.in(far_0_1003_1[0]), .out(far_0_1003_2[0]));    relay_conn far_0_1003_2_b(.in(far_0_1003_1[1]), .out(far_0_1003_2[1]));
    assign layer_0[1003] = ~far_0_1003_2[0]; 
    wire [1:0] far_0_1004_0;    relay_conn far_0_1004_0_a(.in(in[233]), .out(far_0_1004_0[0]));    relay_conn far_0_1004_0_b(.in(in[188]), .out(far_0_1004_0[1]));
    assign layer_0[1004] = far_0_1004_0[1]; 
    wire [1:0] far_0_1005_0;    relay_conn far_0_1005_0_a(.in(in[138]), .out(far_0_1005_0[0]));    relay_conn far_0_1005_0_b(.in(in[204]), .out(far_0_1005_0[1]));
    wire [1:0] far_0_1005_1;    relay_conn far_0_1005_1_a(.in(far_0_1005_0[0]), .out(far_0_1005_1[0]));    relay_conn far_0_1005_1_b(.in(far_0_1005_0[1]), .out(far_0_1005_1[1]));
    assign layer_0[1005] = far_0_1005_1[0] ^ far_0_1005_1[1]; 
    wire [1:0] far_0_1006_0;    relay_conn far_0_1006_0_a(.in(in[23]), .out(far_0_1006_0[0]));    relay_conn far_0_1006_0_b(.in(in[135]), .out(far_0_1006_0[1]));
    wire [1:0] far_0_1006_1;    relay_conn far_0_1006_1_a(.in(far_0_1006_0[0]), .out(far_0_1006_1[0]));    relay_conn far_0_1006_1_b(.in(far_0_1006_0[1]), .out(far_0_1006_1[1]));
    wire [1:0] far_0_1006_2;    relay_conn far_0_1006_2_a(.in(far_0_1006_1[0]), .out(far_0_1006_2[0]));    relay_conn far_0_1006_2_b(.in(far_0_1006_1[1]), .out(far_0_1006_2[1]));
    assign layer_0[1006] = far_0_1006_2[0] & ~far_0_1006_2[1]; 
    wire [1:0] far_0_1007_0;    relay_conn far_0_1007_0_a(.in(in[250]), .out(far_0_1007_0[0]));    relay_conn far_0_1007_0_b(.in(in[175]), .out(far_0_1007_0[1]));
    wire [1:0] far_0_1007_1;    relay_conn far_0_1007_1_a(.in(far_0_1007_0[0]), .out(far_0_1007_1[0]));    relay_conn far_0_1007_1_b(.in(far_0_1007_0[1]), .out(far_0_1007_1[1]));
    assign layer_0[1007] = far_0_1007_1[0] ^ far_0_1007_1[1]; 
    wire [1:0] far_0_1008_0;    relay_conn far_0_1008_0_a(.in(in[57]), .out(far_0_1008_0[0]));    relay_conn far_0_1008_0_b(.in(in[25]), .out(far_0_1008_0[1]));
    assign layer_0[1008] = ~far_0_1008_0[1] | (far_0_1008_0[0] & far_0_1008_0[1]); 
    wire [1:0] far_0_1009_0;    relay_conn far_0_1009_0_a(.in(in[71]), .out(far_0_1009_0[0]));    relay_conn far_0_1009_0_b(.in(in[187]), .out(far_0_1009_0[1]));
    wire [1:0] far_0_1009_1;    relay_conn far_0_1009_1_a(.in(far_0_1009_0[0]), .out(far_0_1009_1[0]));    relay_conn far_0_1009_1_b(.in(far_0_1009_0[1]), .out(far_0_1009_1[1]));
    wire [1:0] far_0_1009_2;    relay_conn far_0_1009_2_a(.in(far_0_1009_1[0]), .out(far_0_1009_2[0]));    relay_conn far_0_1009_2_b(.in(far_0_1009_1[1]), .out(far_0_1009_2[1]));
    assign layer_0[1009] = far_0_1009_2[0] ^ far_0_1009_2[1]; 
    wire [1:0] far_0_1010_0;    relay_conn far_0_1010_0_a(.in(in[111]), .out(far_0_1010_0[0]));    relay_conn far_0_1010_0_b(.in(in[71]), .out(far_0_1010_0[1]));
    assign layer_0[1010] = far_0_1010_0[0] ^ far_0_1010_0[1]; 
    assign layer_0[1011] = in[199] & ~in[204]; 
    wire [1:0] far_0_1012_0;    relay_conn far_0_1012_0_a(.in(in[134]), .out(far_0_1012_0[0]));    relay_conn far_0_1012_0_b(.in(in[67]), .out(far_0_1012_0[1]));
    wire [1:0] far_0_1012_1;    relay_conn far_0_1012_1_a(.in(far_0_1012_0[0]), .out(far_0_1012_1[0]));    relay_conn far_0_1012_1_b(.in(far_0_1012_0[1]), .out(far_0_1012_1[1]));
    assign layer_0[1012] = ~far_0_1012_1[1]; 
    assign layer_0[1013] = ~in[88] | (in[88] & in[99]); 
    assign layer_0[1014] = in[157] | in[187]; 
    wire [1:0] far_0_1015_0;    relay_conn far_0_1015_0_a(.in(in[175]), .out(far_0_1015_0[0]));    relay_conn far_0_1015_0_b(.in(in[241]), .out(far_0_1015_0[1]));
    wire [1:0] far_0_1015_1;    relay_conn far_0_1015_1_a(.in(far_0_1015_0[0]), .out(far_0_1015_1[0]));    relay_conn far_0_1015_1_b(.in(far_0_1015_0[1]), .out(far_0_1015_1[1]));
    assign layer_0[1015] = far_0_1015_1[0] ^ far_0_1015_1[1]; 
    wire [1:0] far_0_1016_0;    relay_conn far_0_1016_0_a(.in(in[239]), .out(far_0_1016_0[0]));    relay_conn far_0_1016_0_b(.in(in[139]), .out(far_0_1016_0[1]));
    wire [1:0] far_0_1016_1;    relay_conn far_0_1016_1_a(.in(far_0_1016_0[0]), .out(far_0_1016_1[0]));    relay_conn far_0_1016_1_b(.in(far_0_1016_0[1]), .out(far_0_1016_1[1]));
    wire [1:0] far_0_1016_2;    relay_conn far_0_1016_2_a(.in(far_0_1016_1[0]), .out(far_0_1016_2[0]));    relay_conn far_0_1016_2_b(.in(far_0_1016_1[1]), .out(far_0_1016_2[1]));
    assign layer_0[1016] = ~(far_0_1016_2[0] | far_0_1016_2[1]); 
    wire [1:0] far_0_1017_0;    relay_conn far_0_1017_0_a(.in(in[27]), .out(far_0_1017_0[0]));    relay_conn far_0_1017_0_b(.in(in[133]), .out(far_0_1017_0[1]));
    wire [1:0] far_0_1017_1;    relay_conn far_0_1017_1_a(.in(far_0_1017_0[0]), .out(far_0_1017_1[0]));    relay_conn far_0_1017_1_b(.in(far_0_1017_0[1]), .out(far_0_1017_1[1]));
    wire [1:0] far_0_1017_2;    relay_conn far_0_1017_2_a(.in(far_0_1017_1[0]), .out(far_0_1017_2[0]));    relay_conn far_0_1017_2_b(.in(far_0_1017_1[1]), .out(far_0_1017_2[1]));
    assign layer_0[1017] = far_0_1017_2[0] ^ far_0_1017_2[1]; 
    wire [1:0] far_0_1018_0;    relay_conn far_0_1018_0_a(.in(in[215]), .out(far_0_1018_0[0]));    relay_conn far_0_1018_0_b(.in(in[142]), .out(far_0_1018_0[1]));
    wire [1:0] far_0_1018_1;    relay_conn far_0_1018_1_a(.in(far_0_1018_0[0]), .out(far_0_1018_1[0]));    relay_conn far_0_1018_1_b(.in(far_0_1018_0[1]), .out(far_0_1018_1[1]));
    assign layer_0[1018] = far_0_1018_1[0]; 
    wire [1:0] far_0_1019_0;    relay_conn far_0_1019_0_a(.in(in[12]), .out(far_0_1019_0[0]));    relay_conn far_0_1019_0_b(.in(in[128]), .out(far_0_1019_0[1]));
    wire [1:0] far_0_1019_1;    relay_conn far_0_1019_1_a(.in(far_0_1019_0[0]), .out(far_0_1019_1[0]));    relay_conn far_0_1019_1_b(.in(far_0_1019_0[1]), .out(far_0_1019_1[1]));
    wire [1:0] far_0_1019_2;    relay_conn far_0_1019_2_a(.in(far_0_1019_1[0]), .out(far_0_1019_2[0]));    relay_conn far_0_1019_2_b(.in(far_0_1019_1[1]), .out(far_0_1019_2[1]));
    assign layer_0[1019] = far_0_1019_2[0] & far_0_1019_2[1]; 
    // Layer 1 ============================================================
    assign layer_1[0] = layer_0[409]; 
    assign layer_1[1] = layer_0[711] & ~layer_0[700]; 
    wire [1:0] far_1_1022_0;    relay_conn far_1_1022_0_a(.in(layer_0[86]), .out(far_1_1022_0[0]));    relay_conn far_1_1022_0_b(.in(layer_0[146]), .out(far_1_1022_0[1]));
    assign layer_1[2] = far_1_1022_0[1]; 
    wire [1:0] far_1_1023_0;    relay_conn far_1_1023_0_a(.in(layer_0[45]), .out(far_1_1023_0[0]));    relay_conn far_1_1023_0_b(.in(layer_0[106]), .out(far_1_1023_0[1]));
    assign layer_1[3] = ~(far_1_1023_0[0] | far_1_1023_0[1]); 
    wire [1:0] far_1_1024_0;    relay_conn far_1_1024_0_a(.in(layer_0[562]), .out(far_1_1024_0[0]));    relay_conn far_1_1024_0_b(.in(layer_0[442]), .out(far_1_1024_0[1]));
    wire [1:0] far_1_1024_1;    relay_conn far_1_1024_1_a(.in(far_1_1024_0[0]), .out(far_1_1024_1[0]));    relay_conn far_1_1024_1_b(.in(far_1_1024_0[1]), .out(far_1_1024_1[1]));
    wire [1:0] far_1_1024_2;    relay_conn far_1_1024_2_a(.in(far_1_1024_1[0]), .out(far_1_1024_2[0]));    relay_conn far_1_1024_2_b(.in(far_1_1024_1[1]), .out(far_1_1024_2[1]));
    assign layer_1[4] = far_1_1024_2[0] | far_1_1024_2[1]; 
    wire [1:0] far_1_1025_0;    relay_conn far_1_1025_0_a(.in(layer_0[480]), .out(far_1_1025_0[0]));    relay_conn far_1_1025_0_b(.in(layer_0[543]), .out(far_1_1025_0[1]));
    assign layer_1[5] = ~far_1_1025_0[0] | (far_1_1025_0[0] & far_1_1025_0[1]); 
    wire [1:0] far_1_1026_0;    relay_conn far_1_1026_0_a(.in(layer_0[419]), .out(far_1_1026_0[0]));    relay_conn far_1_1026_0_b(.in(layer_0[319]), .out(far_1_1026_0[1]));
    wire [1:0] far_1_1026_1;    relay_conn far_1_1026_1_a(.in(far_1_1026_0[0]), .out(far_1_1026_1[0]));    relay_conn far_1_1026_1_b(.in(far_1_1026_0[1]), .out(far_1_1026_1[1]));
    wire [1:0] far_1_1026_2;    relay_conn far_1_1026_2_a(.in(far_1_1026_1[0]), .out(far_1_1026_2[0]));    relay_conn far_1_1026_2_b(.in(far_1_1026_1[1]), .out(far_1_1026_2[1]));
    assign layer_1[6] = ~(far_1_1026_2[0] | far_1_1026_2[1]); 
    wire [1:0] far_1_1027_0;    relay_conn far_1_1027_0_a(.in(layer_0[819]), .out(far_1_1027_0[0]));    relay_conn far_1_1027_0_b(.in(layer_0[861]), .out(far_1_1027_0[1]));
    assign layer_1[7] = ~(far_1_1027_0[0] | far_1_1027_0[1]); 
    wire [1:0] far_1_1028_0;    relay_conn far_1_1028_0_a(.in(layer_0[855]), .out(far_1_1028_0[0]));    relay_conn far_1_1028_0_b(.in(layer_0[795]), .out(far_1_1028_0[1]));
    assign layer_1[8] = ~far_1_1028_0[0] | (far_1_1028_0[0] & far_1_1028_0[1]); 
    wire [1:0] far_1_1029_0;    relay_conn far_1_1029_0_a(.in(layer_0[40]), .out(far_1_1029_0[0]));    relay_conn far_1_1029_0_b(.in(layer_0[125]), .out(far_1_1029_0[1]));
    wire [1:0] far_1_1029_1;    relay_conn far_1_1029_1_a(.in(far_1_1029_0[0]), .out(far_1_1029_1[0]));    relay_conn far_1_1029_1_b(.in(far_1_1029_0[1]), .out(far_1_1029_1[1]));
    assign layer_1[9] = far_1_1029_1[1]; 
    wire [1:0] far_1_1030_0;    relay_conn far_1_1030_0_a(.in(layer_0[419]), .out(far_1_1030_0[0]));    relay_conn far_1_1030_0_b(.in(layer_0[454]), .out(far_1_1030_0[1]));
    assign layer_1[10] = ~far_1_1030_0[1] | (far_1_1030_0[0] & far_1_1030_0[1]); 
    wire [1:0] far_1_1031_0;    relay_conn far_1_1031_0_a(.in(layer_0[512]), .out(far_1_1031_0[0]));    relay_conn far_1_1031_0_b(.in(layer_0[573]), .out(far_1_1031_0[1]));
    assign layer_1[11] = far_1_1031_0[0] & ~far_1_1031_0[1]; 
    wire [1:0] far_1_1032_0;    relay_conn far_1_1032_0_a(.in(layer_0[623]), .out(far_1_1032_0[0]));    relay_conn far_1_1032_0_b(.in(layer_0[675]), .out(far_1_1032_0[1]));
    assign layer_1[12] = far_1_1032_0[0] | far_1_1032_0[1]; 
    wire [1:0] far_1_1033_0;    relay_conn far_1_1033_0_a(.in(layer_0[896]), .out(far_1_1033_0[0]));    relay_conn far_1_1033_0_b(.in(layer_0[786]), .out(far_1_1033_0[1]));
    wire [1:0] far_1_1033_1;    relay_conn far_1_1033_1_a(.in(far_1_1033_0[0]), .out(far_1_1033_1[0]));    relay_conn far_1_1033_1_b(.in(far_1_1033_0[1]), .out(far_1_1033_1[1]));
    wire [1:0] far_1_1033_2;    relay_conn far_1_1033_2_a(.in(far_1_1033_1[0]), .out(far_1_1033_2[0]));    relay_conn far_1_1033_2_b(.in(far_1_1033_1[1]), .out(far_1_1033_2[1]));
    assign layer_1[13] = ~far_1_1033_2[1] | (far_1_1033_2[0] & far_1_1033_2[1]); 
    wire [1:0] far_1_1034_0;    relay_conn far_1_1034_0_a(.in(layer_0[649]), .out(far_1_1034_0[0]));    relay_conn far_1_1034_0_b(.in(layer_0[530]), .out(far_1_1034_0[1]));
    wire [1:0] far_1_1034_1;    relay_conn far_1_1034_1_a(.in(far_1_1034_0[0]), .out(far_1_1034_1[0]));    relay_conn far_1_1034_1_b(.in(far_1_1034_0[1]), .out(far_1_1034_1[1]));
    wire [1:0] far_1_1034_2;    relay_conn far_1_1034_2_a(.in(far_1_1034_1[0]), .out(far_1_1034_2[0]));    relay_conn far_1_1034_2_b(.in(far_1_1034_1[1]), .out(far_1_1034_2[1]));
    assign layer_1[14] = ~(far_1_1034_2[0] | far_1_1034_2[1]); 
    wire [1:0] far_1_1035_0;    relay_conn far_1_1035_0_a(.in(layer_0[356]), .out(far_1_1035_0[0]));    relay_conn far_1_1035_0_b(.in(layer_0[421]), .out(far_1_1035_0[1]));
    wire [1:0] far_1_1035_1;    relay_conn far_1_1035_1_a(.in(far_1_1035_0[0]), .out(far_1_1035_1[0]));    relay_conn far_1_1035_1_b(.in(far_1_1035_0[1]), .out(far_1_1035_1[1]));
    assign layer_1[15] = ~far_1_1035_1[0]; 
    wire [1:0] far_1_1036_0;    relay_conn far_1_1036_0_a(.in(layer_0[666]), .out(far_1_1036_0[0]));    relay_conn far_1_1036_0_b(.in(layer_0[559]), .out(far_1_1036_0[1]));
    wire [1:0] far_1_1036_1;    relay_conn far_1_1036_1_a(.in(far_1_1036_0[0]), .out(far_1_1036_1[0]));    relay_conn far_1_1036_1_b(.in(far_1_1036_0[1]), .out(far_1_1036_1[1]));
    wire [1:0] far_1_1036_2;    relay_conn far_1_1036_2_a(.in(far_1_1036_1[0]), .out(far_1_1036_2[0]));    relay_conn far_1_1036_2_b(.in(far_1_1036_1[1]), .out(far_1_1036_2[1]));
    assign layer_1[16] = far_1_1036_2[1]; 
    wire [1:0] far_1_1037_0;    relay_conn far_1_1037_0_a(.in(layer_0[40]), .out(far_1_1037_0[0]));    relay_conn far_1_1037_0_b(.in(layer_0[76]), .out(far_1_1037_0[1]));
    assign layer_1[17] = ~(far_1_1037_0[0] ^ far_1_1037_0[1]); 
    assign layer_1[18] = layer_0[400] ^ layer_0[395]; 
    assign layer_1[19] = ~(layer_0[770] ^ layer_0[748]); 
    assign layer_1[20] = ~(layer_0[289] ^ layer_0[314]); 
    wire [1:0] far_1_1041_0;    relay_conn far_1_1041_0_a(.in(layer_0[286]), .out(far_1_1041_0[0]));    relay_conn far_1_1041_0_b(.in(layer_0[368]), .out(far_1_1041_0[1]));
    wire [1:0] far_1_1041_1;    relay_conn far_1_1041_1_a(.in(far_1_1041_0[0]), .out(far_1_1041_1[0]));    relay_conn far_1_1041_1_b(.in(far_1_1041_0[1]), .out(far_1_1041_1[1]));
    assign layer_1[21] = far_1_1041_1[0]; 
    wire [1:0] far_1_1042_0;    relay_conn far_1_1042_0_a(.in(layer_0[245]), .out(far_1_1042_0[0]));    relay_conn far_1_1042_0_b(.in(layer_0[339]), .out(far_1_1042_0[1]));
    wire [1:0] far_1_1042_1;    relay_conn far_1_1042_1_a(.in(far_1_1042_0[0]), .out(far_1_1042_1[0]));    relay_conn far_1_1042_1_b(.in(far_1_1042_0[1]), .out(far_1_1042_1[1]));
    assign layer_1[22] = ~far_1_1042_1[1]; 
    assign layer_1[23] = layer_0[891] & ~layer_0[908]; 
    wire [1:0] far_1_1044_0;    relay_conn far_1_1044_0_a(.in(layer_0[544]), .out(far_1_1044_0[0]));    relay_conn far_1_1044_0_b(.in(layer_0[419]), .out(far_1_1044_0[1]));
    wire [1:0] far_1_1044_1;    relay_conn far_1_1044_1_a(.in(far_1_1044_0[0]), .out(far_1_1044_1[0]));    relay_conn far_1_1044_1_b(.in(far_1_1044_0[1]), .out(far_1_1044_1[1]));
    wire [1:0] far_1_1044_2;    relay_conn far_1_1044_2_a(.in(far_1_1044_1[0]), .out(far_1_1044_2[0]));    relay_conn far_1_1044_2_b(.in(far_1_1044_1[1]), .out(far_1_1044_2[1]));
    assign layer_1[24] = ~(far_1_1044_2[0] & far_1_1044_2[1]); 
    wire [1:0] far_1_1045_0;    relay_conn far_1_1045_0_a(.in(layer_0[157]), .out(far_1_1045_0[0]));    relay_conn far_1_1045_0_b(.in(layer_0[95]), .out(far_1_1045_0[1]));
    assign layer_1[25] = ~(far_1_1045_0[0] ^ far_1_1045_0[1]); 
    assign layer_1[26] = layer_0[449] & layer_0[438]; 
    assign layer_1[27] = layer_0[70] & ~layer_0[91]; 
    wire [1:0] far_1_1048_0;    relay_conn far_1_1048_0_a(.in(layer_0[116]), .out(far_1_1048_0[0]));    relay_conn far_1_1048_0_b(.in(layer_0[8]), .out(far_1_1048_0[1]));
    wire [1:0] far_1_1048_1;    relay_conn far_1_1048_1_a(.in(far_1_1048_0[0]), .out(far_1_1048_1[0]));    relay_conn far_1_1048_1_b(.in(far_1_1048_0[1]), .out(far_1_1048_1[1]));
    wire [1:0] far_1_1048_2;    relay_conn far_1_1048_2_a(.in(far_1_1048_1[0]), .out(far_1_1048_2[0]));    relay_conn far_1_1048_2_b(.in(far_1_1048_1[1]), .out(far_1_1048_2[1]));
    assign layer_1[28] = far_1_1048_2[0] ^ far_1_1048_2[1]; 
    wire [1:0] far_1_1049_0;    relay_conn far_1_1049_0_a(.in(layer_0[923]), .out(far_1_1049_0[0]));    relay_conn far_1_1049_0_b(.in(layer_0[821]), .out(far_1_1049_0[1]));
    wire [1:0] far_1_1049_1;    relay_conn far_1_1049_1_a(.in(far_1_1049_0[0]), .out(far_1_1049_1[0]));    relay_conn far_1_1049_1_b(.in(far_1_1049_0[1]), .out(far_1_1049_1[1]));
    wire [1:0] far_1_1049_2;    relay_conn far_1_1049_2_a(.in(far_1_1049_1[0]), .out(far_1_1049_2[0]));    relay_conn far_1_1049_2_b(.in(far_1_1049_1[1]), .out(far_1_1049_2[1]));
    assign layer_1[29] = far_1_1049_2[0] & ~far_1_1049_2[1]; 
    wire [1:0] far_1_1050_0;    relay_conn far_1_1050_0_a(.in(layer_0[898]), .out(far_1_1050_0[0]));    relay_conn far_1_1050_0_b(.in(layer_0[1000]), .out(far_1_1050_0[1]));
    wire [1:0] far_1_1050_1;    relay_conn far_1_1050_1_a(.in(far_1_1050_0[0]), .out(far_1_1050_1[0]));    relay_conn far_1_1050_1_b(.in(far_1_1050_0[1]), .out(far_1_1050_1[1]));
    wire [1:0] far_1_1050_2;    relay_conn far_1_1050_2_a(.in(far_1_1050_1[0]), .out(far_1_1050_2[0]));    relay_conn far_1_1050_2_b(.in(far_1_1050_1[1]), .out(far_1_1050_2[1]));
    assign layer_1[30] = far_1_1050_2[0]; 
    assign layer_1[31] = ~layer_0[511] | (layer_0[488] & layer_0[511]); 
    wire [1:0] far_1_1052_0;    relay_conn far_1_1052_0_a(.in(layer_0[580]), .out(far_1_1052_0[0]));    relay_conn far_1_1052_0_b(.in(layer_0[457]), .out(far_1_1052_0[1]));
    wire [1:0] far_1_1052_1;    relay_conn far_1_1052_1_a(.in(far_1_1052_0[0]), .out(far_1_1052_1[0]));    relay_conn far_1_1052_1_b(.in(far_1_1052_0[1]), .out(far_1_1052_1[1]));
    wire [1:0] far_1_1052_2;    relay_conn far_1_1052_2_a(.in(far_1_1052_1[0]), .out(far_1_1052_2[0]));    relay_conn far_1_1052_2_b(.in(far_1_1052_1[1]), .out(far_1_1052_2[1]));
    assign layer_1[32] = ~(far_1_1052_2[0] & far_1_1052_2[1]); 
    wire [1:0] far_1_1053_0;    relay_conn far_1_1053_0_a(.in(layer_0[477]), .out(far_1_1053_0[0]));    relay_conn far_1_1053_0_b(.in(layer_0[381]), .out(far_1_1053_0[1]));
    wire [1:0] far_1_1053_1;    relay_conn far_1_1053_1_a(.in(far_1_1053_0[0]), .out(far_1_1053_1[0]));    relay_conn far_1_1053_1_b(.in(far_1_1053_0[1]), .out(far_1_1053_1[1]));
    wire [1:0] far_1_1053_2;    relay_conn far_1_1053_2_a(.in(far_1_1053_1[0]), .out(far_1_1053_2[0]));    relay_conn far_1_1053_2_b(.in(far_1_1053_1[1]), .out(far_1_1053_2[1]));
    assign layer_1[33] = ~(far_1_1053_2[0] | far_1_1053_2[1]); 
    wire [1:0] far_1_1054_0;    relay_conn far_1_1054_0_a(.in(layer_0[28]), .out(far_1_1054_0[0]));    relay_conn far_1_1054_0_b(.in(layer_0[129]), .out(far_1_1054_0[1]));
    wire [1:0] far_1_1054_1;    relay_conn far_1_1054_1_a(.in(far_1_1054_0[0]), .out(far_1_1054_1[0]));    relay_conn far_1_1054_1_b(.in(far_1_1054_0[1]), .out(far_1_1054_1[1]));
    wire [1:0] far_1_1054_2;    relay_conn far_1_1054_2_a(.in(far_1_1054_1[0]), .out(far_1_1054_2[0]));    relay_conn far_1_1054_2_b(.in(far_1_1054_1[1]), .out(far_1_1054_2[1]));
    assign layer_1[34] = far_1_1054_2[0] & far_1_1054_2[1]; 
    wire [1:0] far_1_1055_0;    relay_conn far_1_1055_0_a(.in(layer_0[208]), .out(far_1_1055_0[0]));    relay_conn far_1_1055_0_b(.in(layer_0[160]), .out(far_1_1055_0[1]));
    assign layer_1[35] = ~far_1_1055_0[0]; 
    wire [1:0] far_1_1056_0;    relay_conn far_1_1056_0_a(.in(layer_0[178]), .out(far_1_1056_0[0]));    relay_conn far_1_1056_0_b(.in(layer_0[263]), .out(far_1_1056_0[1]));
    wire [1:0] far_1_1056_1;    relay_conn far_1_1056_1_a(.in(far_1_1056_0[0]), .out(far_1_1056_1[0]));    relay_conn far_1_1056_1_b(.in(far_1_1056_0[1]), .out(far_1_1056_1[1]));
    assign layer_1[36] = far_1_1056_1[1] & ~far_1_1056_1[0]; 
    wire [1:0] far_1_1057_0;    relay_conn far_1_1057_0_a(.in(layer_0[126]), .out(far_1_1057_0[0]));    relay_conn far_1_1057_0_b(.in(layer_0[186]), .out(far_1_1057_0[1]));
    assign layer_1[37] = far_1_1057_0[0] & far_1_1057_0[1]; 
    wire [1:0] far_1_1058_0;    relay_conn far_1_1058_0_a(.in(layer_0[438]), .out(far_1_1058_0[0]));    relay_conn far_1_1058_0_b(.in(layer_0[380]), .out(far_1_1058_0[1]));
    assign layer_1[38] = far_1_1058_0[1]; 
    wire [1:0] far_1_1059_0;    relay_conn far_1_1059_0_a(.in(layer_0[877]), .out(far_1_1059_0[0]));    relay_conn far_1_1059_0_b(.in(layer_0[843]), .out(far_1_1059_0[1]));
    assign layer_1[39] = far_1_1059_0[0] & ~far_1_1059_0[1]; 
    wire [1:0] far_1_1060_0;    relay_conn far_1_1060_0_a(.in(layer_0[924]), .out(far_1_1060_0[0]));    relay_conn far_1_1060_0_b(.in(layer_0[826]), .out(far_1_1060_0[1]));
    wire [1:0] far_1_1060_1;    relay_conn far_1_1060_1_a(.in(far_1_1060_0[0]), .out(far_1_1060_1[0]));    relay_conn far_1_1060_1_b(.in(far_1_1060_0[1]), .out(far_1_1060_1[1]));
    wire [1:0] far_1_1060_2;    relay_conn far_1_1060_2_a(.in(far_1_1060_1[0]), .out(far_1_1060_2[0]));    relay_conn far_1_1060_2_b(.in(far_1_1060_1[1]), .out(far_1_1060_2[1]));
    assign layer_1[40] = far_1_1060_2[0]; 
    wire [1:0] far_1_1061_0;    relay_conn far_1_1061_0_a(.in(layer_0[111]), .out(far_1_1061_0[0]));    relay_conn far_1_1061_0_b(.in(layer_0[172]), .out(far_1_1061_0[1]));
    assign layer_1[41] = ~(far_1_1061_0[0] | far_1_1061_0[1]); 
    wire [1:0] far_1_1062_0;    relay_conn far_1_1062_0_a(.in(layer_0[853]), .out(far_1_1062_0[0]));    relay_conn far_1_1062_0_b(.in(layer_0[793]), .out(far_1_1062_0[1]));
    assign layer_1[42] = ~(far_1_1062_0[0] ^ far_1_1062_0[1]); 
    wire [1:0] far_1_1063_0;    relay_conn far_1_1063_0_a(.in(layer_0[1016]), .out(far_1_1063_0[0]));    relay_conn far_1_1063_0_b(.in(layer_0[901]), .out(far_1_1063_0[1]));
    wire [1:0] far_1_1063_1;    relay_conn far_1_1063_1_a(.in(far_1_1063_0[0]), .out(far_1_1063_1[0]));    relay_conn far_1_1063_1_b(.in(far_1_1063_0[1]), .out(far_1_1063_1[1]));
    wire [1:0] far_1_1063_2;    relay_conn far_1_1063_2_a(.in(far_1_1063_1[0]), .out(far_1_1063_2[0]));    relay_conn far_1_1063_2_b(.in(far_1_1063_1[1]), .out(far_1_1063_2[1]));
    assign layer_1[43] = far_1_1063_2[0] | far_1_1063_2[1]; 
    wire [1:0] far_1_1064_0;    relay_conn far_1_1064_0_a(.in(layer_0[773]), .out(far_1_1064_0[0]));    relay_conn far_1_1064_0_b(.in(layer_0[694]), .out(far_1_1064_0[1]));
    wire [1:0] far_1_1064_1;    relay_conn far_1_1064_1_a(.in(far_1_1064_0[0]), .out(far_1_1064_1[0]));    relay_conn far_1_1064_1_b(.in(far_1_1064_0[1]), .out(far_1_1064_1[1]));
    assign layer_1[44] = far_1_1064_1[0] ^ far_1_1064_1[1]; 
    assign layer_1[45] = ~layer_0[966] | (layer_0[966] & layer_0[973]); 
    wire [1:0] far_1_1066_0;    relay_conn far_1_1066_0_a(.in(layer_0[798]), .out(far_1_1066_0[0]));    relay_conn far_1_1066_0_b(.in(layer_0[710]), .out(far_1_1066_0[1]));
    wire [1:0] far_1_1066_1;    relay_conn far_1_1066_1_a(.in(far_1_1066_0[0]), .out(far_1_1066_1[0]));    relay_conn far_1_1066_1_b(.in(far_1_1066_0[1]), .out(far_1_1066_1[1]));
    assign layer_1[46] = ~far_1_1066_1[1] | (far_1_1066_1[0] & far_1_1066_1[1]); 
    wire [1:0] far_1_1067_0;    relay_conn far_1_1067_0_a(.in(layer_0[43]), .out(far_1_1067_0[0]));    relay_conn far_1_1067_0_b(.in(layer_0[148]), .out(far_1_1067_0[1]));
    wire [1:0] far_1_1067_1;    relay_conn far_1_1067_1_a(.in(far_1_1067_0[0]), .out(far_1_1067_1[0]));    relay_conn far_1_1067_1_b(.in(far_1_1067_0[1]), .out(far_1_1067_1[1]));
    wire [1:0] far_1_1067_2;    relay_conn far_1_1067_2_a(.in(far_1_1067_1[0]), .out(far_1_1067_2[0]));    relay_conn far_1_1067_2_b(.in(far_1_1067_1[1]), .out(far_1_1067_2[1]));
    assign layer_1[47] = far_1_1067_2[1] & ~far_1_1067_2[0]; 
    wire [1:0] far_1_1068_0;    relay_conn far_1_1068_0_a(.in(layer_0[495]), .out(far_1_1068_0[0]));    relay_conn far_1_1068_0_b(.in(layer_0[385]), .out(far_1_1068_0[1]));
    wire [1:0] far_1_1068_1;    relay_conn far_1_1068_1_a(.in(far_1_1068_0[0]), .out(far_1_1068_1[0]));    relay_conn far_1_1068_1_b(.in(far_1_1068_0[1]), .out(far_1_1068_1[1]));
    wire [1:0] far_1_1068_2;    relay_conn far_1_1068_2_a(.in(far_1_1068_1[0]), .out(far_1_1068_2[0]));    relay_conn far_1_1068_2_b(.in(far_1_1068_1[1]), .out(far_1_1068_2[1]));
    assign layer_1[48] = far_1_1068_2[0] ^ far_1_1068_2[1]; 
    assign layer_1[49] = layer_0[436] | layer_0[461]; 
    wire [1:0] far_1_1070_0;    relay_conn far_1_1070_0_a(.in(layer_0[277]), .out(far_1_1070_0[0]));    relay_conn far_1_1070_0_b(.in(layer_0[226]), .out(far_1_1070_0[1]));
    assign layer_1[50] = far_1_1070_0[0] & far_1_1070_0[1]; 
    wire [1:0] far_1_1071_0;    relay_conn far_1_1071_0_a(.in(layer_0[741]), .out(far_1_1071_0[0]));    relay_conn far_1_1071_0_b(.in(layer_0[708]), .out(far_1_1071_0[1]));
    assign layer_1[51] = ~(far_1_1071_0[0] & far_1_1071_0[1]); 
    assign layer_1[52] = ~(layer_0[127] | layer_0[109]); 
    wire [1:0] far_1_1073_0;    relay_conn far_1_1073_0_a(.in(layer_0[137]), .out(far_1_1073_0[0]));    relay_conn far_1_1073_0_b(.in(layer_0[187]), .out(far_1_1073_0[1]));
    assign layer_1[53] = far_1_1073_0[0] | far_1_1073_0[1]; 
    wire [1:0] far_1_1074_0;    relay_conn far_1_1074_0_a(.in(layer_0[614]), .out(far_1_1074_0[0]));    relay_conn far_1_1074_0_b(.in(layer_0[493]), .out(far_1_1074_0[1]));
    wire [1:0] far_1_1074_1;    relay_conn far_1_1074_1_a(.in(far_1_1074_0[0]), .out(far_1_1074_1[0]));    relay_conn far_1_1074_1_b(.in(far_1_1074_0[1]), .out(far_1_1074_1[1]));
    wire [1:0] far_1_1074_2;    relay_conn far_1_1074_2_a(.in(far_1_1074_1[0]), .out(far_1_1074_2[0]));    relay_conn far_1_1074_2_b(.in(far_1_1074_1[1]), .out(far_1_1074_2[1]));
    assign layer_1[54] = far_1_1074_2[0]; 
    wire [1:0] far_1_1075_0;    relay_conn far_1_1075_0_a(.in(layer_0[144]), .out(far_1_1075_0[0]));    relay_conn far_1_1075_0_b(.in(layer_0[56]), .out(far_1_1075_0[1]));
    wire [1:0] far_1_1075_1;    relay_conn far_1_1075_1_a(.in(far_1_1075_0[0]), .out(far_1_1075_1[0]));    relay_conn far_1_1075_1_b(.in(far_1_1075_0[1]), .out(far_1_1075_1[1]));
    assign layer_1[55] = ~(far_1_1075_1[0] & far_1_1075_1[1]); 
    wire [1:0] far_1_1076_0;    relay_conn far_1_1076_0_a(.in(layer_0[954]), .out(far_1_1076_0[0]));    relay_conn far_1_1076_0_b(.in(layer_0[997]), .out(far_1_1076_0[1]));
    assign layer_1[56] = ~(far_1_1076_0[0] ^ far_1_1076_0[1]); 
    wire [1:0] far_1_1077_0;    relay_conn far_1_1077_0_a(.in(layer_0[279]), .out(far_1_1077_0[0]));    relay_conn far_1_1077_0_b(.in(layer_0[407]), .out(far_1_1077_0[1]));
    wire [1:0] far_1_1077_1;    relay_conn far_1_1077_1_a(.in(far_1_1077_0[0]), .out(far_1_1077_1[0]));    relay_conn far_1_1077_1_b(.in(far_1_1077_0[1]), .out(far_1_1077_1[1]));
    wire [1:0] far_1_1077_2;    relay_conn far_1_1077_2_a(.in(far_1_1077_1[0]), .out(far_1_1077_2[0]));    relay_conn far_1_1077_2_b(.in(far_1_1077_1[1]), .out(far_1_1077_2[1]));
    wire [1:0] far_1_1077_3;    relay_conn far_1_1077_3_a(.in(far_1_1077_2[0]), .out(far_1_1077_3[0]));    relay_conn far_1_1077_3_b(.in(far_1_1077_2[1]), .out(far_1_1077_3[1]));
    assign layer_1[57] = ~(far_1_1077_3[0] | far_1_1077_3[1]); 
    assign layer_1[58] = layer_0[612] | layer_0[630]; 
    assign layer_1[59] = layer_0[28] & layer_0[1]; 
    assign layer_1[60] = layer_0[57] & ~layer_0[84]; 
    wire [1:0] far_1_1081_0;    relay_conn far_1_1081_0_a(.in(layer_0[867]), .out(far_1_1081_0[0]));    relay_conn far_1_1081_0_b(.in(layer_0[819]), .out(far_1_1081_0[1]));
    assign layer_1[61] = ~far_1_1081_0[0] | (far_1_1081_0[0] & far_1_1081_0[1]); 
    assign layer_1[62] = ~(layer_0[220] & layer_0[212]); 
    wire [1:0] far_1_1083_0;    relay_conn far_1_1083_0_a(.in(layer_0[211]), .out(far_1_1083_0[0]));    relay_conn far_1_1083_0_b(.in(layer_0[330]), .out(far_1_1083_0[1]));
    wire [1:0] far_1_1083_1;    relay_conn far_1_1083_1_a(.in(far_1_1083_0[0]), .out(far_1_1083_1[0]));    relay_conn far_1_1083_1_b(.in(far_1_1083_0[1]), .out(far_1_1083_1[1]));
    wire [1:0] far_1_1083_2;    relay_conn far_1_1083_2_a(.in(far_1_1083_1[0]), .out(far_1_1083_2[0]));    relay_conn far_1_1083_2_b(.in(far_1_1083_1[1]), .out(far_1_1083_2[1]));
    assign layer_1[63] = ~far_1_1083_2[0]; 
    wire [1:0] far_1_1084_0;    relay_conn far_1_1084_0_a(.in(layer_0[452]), .out(far_1_1084_0[0]));    relay_conn far_1_1084_0_b(.in(layer_0[565]), .out(far_1_1084_0[1]));
    wire [1:0] far_1_1084_1;    relay_conn far_1_1084_1_a(.in(far_1_1084_0[0]), .out(far_1_1084_1[0]));    relay_conn far_1_1084_1_b(.in(far_1_1084_0[1]), .out(far_1_1084_1[1]));
    wire [1:0] far_1_1084_2;    relay_conn far_1_1084_2_a(.in(far_1_1084_1[0]), .out(far_1_1084_2[0]));    relay_conn far_1_1084_2_b(.in(far_1_1084_1[1]), .out(far_1_1084_2[1]));
    assign layer_1[64] = far_1_1084_2[1]; 
    assign layer_1[65] = layer_0[380] & ~layer_0[384]; 
    wire [1:0] far_1_1086_0;    relay_conn far_1_1086_0_a(.in(layer_0[346]), .out(far_1_1086_0[0]));    relay_conn far_1_1086_0_b(.in(layer_0[284]), .out(far_1_1086_0[1]));
    assign layer_1[66] = far_1_1086_0[0] & ~far_1_1086_0[1]; 
    assign layer_1[67] = ~layer_0[789] | (layer_0[789] & layer_0[770]); 
    assign layer_1[68] = ~(layer_0[70] | layer_0[42]); 
    assign layer_1[69] = ~layer_0[56]; 
    wire [1:0] far_1_1090_0;    relay_conn far_1_1090_0_a(.in(layer_0[34]), .out(far_1_1090_0[0]));    relay_conn far_1_1090_0_b(.in(layer_0[93]), .out(far_1_1090_0[1]));
    assign layer_1[70] = ~far_1_1090_0[0]; 
    wire [1:0] far_1_1091_0;    relay_conn far_1_1091_0_a(.in(layer_0[348]), .out(far_1_1091_0[0]));    relay_conn far_1_1091_0_b(.in(layer_0[419]), .out(far_1_1091_0[1]));
    wire [1:0] far_1_1091_1;    relay_conn far_1_1091_1_a(.in(far_1_1091_0[0]), .out(far_1_1091_1[0]));    relay_conn far_1_1091_1_b(.in(far_1_1091_0[1]), .out(far_1_1091_1[1]));
    assign layer_1[71] = ~far_1_1091_1[1] | (far_1_1091_1[0] & far_1_1091_1[1]); 
    wire [1:0] far_1_1092_0;    relay_conn far_1_1092_0_a(.in(layer_0[35]), .out(far_1_1092_0[0]));    relay_conn far_1_1092_0_b(.in(layer_0[68]), .out(far_1_1092_0[1]));
    assign layer_1[72] = ~(far_1_1092_0[0] & far_1_1092_0[1]); 
    assign layer_1[73] = ~(layer_0[124] & layer_0[108]); 
    wire [1:0] far_1_1094_0;    relay_conn far_1_1094_0_a(.in(layer_0[219]), .out(far_1_1094_0[0]));    relay_conn far_1_1094_0_b(.in(layer_0[336]), .out(far_1_1094_0[1]));
    wire [1:0] far_1_1094_1;    relay_conn far_1_1094_1_a(.in(far_1_1094_0[0]), .out(far_1_1094_1[0]));    relay_conn far_1_1094_1_b(.in(far_1_1094_0[1]), .out(far_1_1094_1[1]));
    wire [1:0] far_1_1094_2;    relay_conn far_1_1094_2_a(.in(far_1_1094_1[0]), .out(far_1_1094_2[0]));    relay_conn far_1_1094_2_b(.in(far_1_1094_1[1]), .out(far_1_1094_2[1]));
    assign layer_1[74] = far_1_1094_2[0] | far_1_1094_2[1]; 
    wire [1:0] far_1_1095_0;    relay_conn far_1_1095_0_a(.in(layer_0[231]), .out(far_1_1095_0[0]));    relay_conn far_1_1095_0_b(.in(layer_0[345]), .out(far_1_1095_0[1]));
    wire [1:0] far_1_1095_1;    relay_conn far_1_1095_1_a(.in(far_1_1095_0[0]), .out(far_1_1095_1[0]));    relay_conn far_1_1095_1_b(.in(far_1_1095_0[1]), .out(far_1_1095_1[1]));
    wire [1:0] far_1_1095_2;    relay_conn far_1_1095_2_a(.in(far_1_1095_1[0]), .out(far_1_1095_2[0]));    relay_conn far_1_1095_2_b(.in(far_1_1095_1[1]), .out(far_1_1095_2[1]));
    assign layer_1[75] = far_1_1095_2[1]; 
    assign layer_1[76] = layer_0[307]; 
    wire [1:0] far_1_1097_0;    relay_conn far_1_1097_0_a(.in(layer_0[272]), .out(far_1_1097_0[0]));    relay_conn far_1_1097_0_b(.in(layer_0[384]), .out(far_1_1097_0[1]));
    wire [1:0] far_1_1097_1;    relay_conn far_1_1097_1_a(.in(far_1_1097_0[0]), .out(far_1_1097_1[0]));    relay_conn far_1_1097_1_b(.in(far_1_1097_0[1]), .out(far_1_1097_1[1]));
    wire [1:0] far_1_1097_2;    relay_conn far_1_1097_2_a(.in(far_1_1097_1[0]), .out(far_1_1097_2[0]));    relay_conn far_1_1097_2_b(.in(far_1_1097_1[1]), .out(far_1_1097_2[1]));
    assign layer_1[77] = far_1_1097_2[1]; 
    wire [1:0] far_1_1098_0;    relay_conn far_1_1098_0_a(.in(layer_0[741]), .out(far_1_1098_0[0]));    relay_conn far_1_1098_0_b(.in(layer_0[786]), .out(far_1_1098_0[1]));
    assign layer_1[78] = ~(far_1_1098_0[0] & far_1_1098_0[1]); 
    wire [1:0] far_1_1099_0;    relay_conn far_1_1099_0_a(.in(layer_0[710]), .out(far_1_1099_0[0]));    relay_conn far_1_1099_0_b(.in(layer_0[770]), .out(far_1_1099_0[1]));
    assign layer_1[79] = ~far_1_1099_0[1]; 
    wire [1:0] far_1_1100_0;    relay_conn far_1_1100_0_a(.in(layer_0[404]), .out(far_1_1100_0[0]));    relay_conn far_1_1100_0_b(.in(layer_0[461]), .out(far_1_1100_0[1]));
    assign layer_1[80] = ~far_1_1100_0[0]; 
    wire [1:0] far_1_1101_0;    relay_conn far_1_1101_0_a(.in(layer_0[504]), .out(far_1_1101_0[0]));    relay_conn far_1_1101_0_b(.in(layer_0[617]), .out(far_1_1101_0[1]));
    wire [1:0] far_1_1101_1;    relay_conn far_1_1101_1_a(.in(far_1_1101_0[0]), .out(far_1_1101_1[0]));    relay_conn far_1_1101_1_b(.in(far_1_1101_0[1]), .out(far_1_1101_1[1]));
    wire [1:0] far_1_1101_2;    relay_conn far_1_1101_2_a(.in(far_1_1101_1[0]), .out(far_1_1101_2[0]));    relay_conn far_1_1101_2_b(.in(far_1_1101_1[1]), .out(far_1_1101_2[1]));
    assign layer_1[81] = ~far_1_1101_2[0] | (far_1_1101_2[0] & far_1_1101_2[1]); 
    assign layer_1[82] = ~layer_0[265]; 
    wire [1:0] far_1_1103_0;    relay_conn far_1_1103_0_a(.in(layer_0[774]), .out(far_1_1103_0[0]));    relay_conn far_1_1103_0_b(.in(layer_0[816]), .out(far_1_1103_0[1]));
    assign layer_1[83] = far_1_1103_0[0] | far_1_1103_0[1]; 
    wire [1:0] far_1_1104_0;    relay_conn far_1_1104_0_a(.in(layer_0[361]), .out(far_1_1104_0[0]));    relay_conn far_1_1104_0_b(.in(layer_0[474]), .out(far_1_1104_0[1]));
    wire [1:0] far_1_1104_1;    relay_conn far_1_1104_1_a(.in(far_1_1104_0[0]), .out(far_1_1104_1[0]));    relay_conn far_1_1104_1_b(.in(far_1_1104_0[1]), .out(far_1_1104_1[1]));
    wire [1:0] far_1_1104_2;    relay_conn far_1_1104_2_a(.in(far_1_1104_1[0]), .out(far_1_1104_2[0]));    relay_conn far_1_1104_2_b(.in(far_1_1104_1[1]), .out(far_1_1104_2[1]));
    assign layer_1[84] = ~(far_1_1104_2[0] | far_1_1104_2[1]); 
    assign layer_1[85] = layer_0[886]; 
    wire [1:0] far_1_1106_0;    relay_conn far_1_1106_0_a(.in(layer_0[496]), .out(far_1_1106_0[0]));    relay_conn far_1_1106_0_b(.in(layer_0[456]), .out(far_1_1106_0[1]));
    assign layer_1[86] = ~far_1_1106_0[1] | (far_1_1106_0[0] & far_1_1106_0[1]); 
    wire [1:0] far_1_1107_0;    relay_conn far_1_1107_0_a(.in(layer_0[735]), .out(far_1_1107_0[0]));    relay_conn far_1_1107_0_b(.in(layer_0[768]), .out(far_1_1107_0[1]));
    assign layer_1[87] = ~far_1_1107_0[1]; 
    wire [1:0] far_1_1108_0;    relay_conn far_1_1108_0_a(.in(layer_0[928]), .out(far_1_1108_0[0]));    relay_conn far_1_1108_0_b(.in(layer_0[1019]), .out(far_1_1108_0[1]));
    wire [1:0] far_1_1108_1;    relay_conn far_1_1108_1_a(.in(far_1_1108_0[0]), .out(far_1_1108_1[0]));    relay_conn far_1_1108_1_b(.in(far_1_1108_0[1]), .out(far_1_1108_1[1]));
    assign layer_1[88] = ~far_1_1108_1[0]; 
    assign layer_1[89] = ~layer_0[908]; 
    wire [1:0] far_1_1110_0;    relay_conn far_1_1110_0_a(.in(layer_0[272]), .out(far_1_1110_0[0]));    relay_conn far_1_1110_0_b(.in(layer_0[369]), .out(far_1_1110_0[1]));
    wire [1:0] far_1_1110_1;    relay_conn far_1_1110_1_a(.in(far_1_1110_0[0]), .out(far_1_1110_1[0]));    relay_conn far_1_1110_1_b(.in(far_1_1110_0[1]), .out(far_1_1110_1[1]));
    wire [1:0] far_1_1110_2;    relay_conn far_1_1110_2_a(.in(far_1_1110_1[0]), .out(far_1_1110_2[0]));    relay_conn far_1_1110_2_b(.in(far_1_1110_1[1]), .out(far_1_1110_2[1]));
    assign layer_1[90] = ~(far_1_1110_2[0] & far_1_1110_2[1]); 
    assign layer_1[91] = ~layer_0[855]; 
    assign layer_1[92] = ~layer_0[11]; 
    wire [1:0] far_1_1113_0;    relay_conn far_1_1113_0_a(.in(layer_0[513]), .out(far_1_1113_0[0]));    relay_conn far_1_1113_0_b(.in(layer_0[400]), .out(far_1_1113_0[1]));
    wire [1:0] far_1_1113_1;    relay_conn far_1_1113_1_a(.in(far_1_1113_0[0]), .out(far_1_1113_1[0]));    relay_conn far_1_1113_1_b(.in(far_1_1113_0[1]), .out(far_1_1113_1[1]));
    wire [1:0] far_1_1113_2;    relay_conn far_1_1113_2_a(.in(far_1_1113_1[0]), .out(far_1_1113_2[0]));    relay_conn far_1_1113_2_b(.in(far_1_1113_1[1]), .out(far_1_1113_2[1]));
    assign layer_1[93] = ~far_1_1113_2[0] | (far_1_1113_2[0] & far_1_1113_2[1]); 
    wire [1:0] far_1_1114_0;    relay_conn far_1_1114_0_a(.in(layer_0[983]), .out(far_1_1114_0[0]));    relay_conn far_1_1114_0_b(.in(layer_0[886]), .out(far_1_1114_0[1]));
    wire [1:0] far_1_1114_1;    relay_conn far_1_1114_1_a(.in(far_1_1114_0[0]), .out(far_1_1114_1[0]));    relay_conn far_1_1114_1_b(.in(far_1_1114_0[1]), .out(far_1_1114_1[1]));
    wire [1:0] far_1_1114_2;    relay_conn far_1_1114_2_a(.in(far_1_1114_1[0]), .out(far_1_1114_2[0]));    relay_conn far_1_1114_2_b(.in(far_1_1114_1[1]), .out(far_1_1114_2[1]));
    assign layer_1[94] = ~(far_1_1114_2[0] & far_1_1114_2[1]); 
    assign layer_1[95] = ~layer_0[322] | (layer_0[322] & layer_0[339]); 
    assign layer_1[96] = ~layer_0[839]; 
    wire [1:0] far_1_1117_0;    relay_conn far_1_1117_0_a(.in(layer_0[544]), .out(far_1_1117_0[0]));    relay_conn far_1_1117_0_b(.in(layer_0[461]), .out(far_1_1117_0[1]));
    wire [1:0] far_1_1117_1;    relay_conn far_1_1117_1_a(.in(far_1_1117_0[0]), .out(far_1_1117_1[0]));    relay_conn far_1_1117_1_b(.in(far_1_1117_0[1]), .out(far_1_1117_1[1]));
    assign layer_1[97] = ~(far_1_1117_1[0] & far_1_1117_1[1]); 
    wire [1:0] far_1_1118_0;    relay_conn far_1_1118_0_a(.in(layer_0[898]), .out(far_1_1118_0[0]));    relay_conn far_1_1118_0_b(.in(layer_0[1004]), .out(far_1_1118_0[1]));
    wire [1:0] far_1_1118_1;    relay_conn far_1_1118_1_a(.in(far_1_1118_0[0]), .out(far_1_1118_1[0]));    relay_conn far_1_1118_1_b(.in(far_1_1118_0[1]), .out(far_1_1118_1[1]));
    wire [1:0] far_1_1118_2;    relay_conn far_1_1118_2_a(.in(far_1_1118_1[0]), .out(far_1_1118_2[0]));    relay_conn far_1_1118_2_b(.in(far_1_1118_1[1]), .out(far_1_1118_2[1]));
    assign layer_1[98] = far_1_1118_2[0] & far_1_1118_2[1]; 
    assign layer_1[99] = ~layer_0[565]; 
    wire [1:0] far_1_1120_0;    relay_conn far_1_1120_0_a(.in(layer_0[639]), .out(far_1_1120_0[0]));    relay_conn far_1_1120_0_b(.in(layer_0[579]), .out(far_1_1120_0[1]));
    assign layer_1[100] = far_1_1120_0[0] & far_1_1120_0[1]; 
    wire [1:0] far_1_1121_0;    relay_conn far_1_1121_0_a(.in(layer_0[914]), .out(far_1_1121_0[0]));    relay_conn far_1_1121_0_b(.in(layer_0[978]), .out(far_1_1121_0[1]));
    wire [1:0] far_1_1121_1;    relay_conn far_1_1121_1_a(.in(far_1_1121_0[0]), .out(far_1_1121_1[0]));    relay_conn far_1_1121_1_b(.in(far_1_1121_0[1]), .out(far_1_1121_1[1]));
    assign layer_1[101] = far_1_1121_1[0]; 
    wire [1:0] far_1_1122_0;    relay_conn far_1_1122_0_a(.in(layer_0[468]), .out(far_1_1122_0[0]));    relay_conn far_1_1122_0_b(.in(layer_0[587]), .out(far_1_1122_0[1]));
    wire [1:0] far_1_1122_1;    relay_conn far_1_1122_1_a(.in(far_1_1122_0[0]), .out(far_1_1122_1[0]));    relay_conn far_1_1122_1_b(.in(far_1_1122_0[1]), .out(far_1_1122_1[1]));
    wire [1:0] far_1_1122_2;    relay_conn far_1_1122_2_a(.in(far_1_1122_1[0]), .out(far_1_1122_2[0]));    relay_conn far_1_1122_2_b(.in(far_1_1122_1[1]), .out(far_1_1122_2[1]));
    assign layer_1[102] = far_1_1122_2[1]; 
    wire [1:0] far_1_1123_0;    relay_conn far_1_1123_0_a(.in(layer_0[591]), .out(far_1_1123_0[0]));    relay_conn far_1_1123_0_b(.in(layer_0[478]), .out(far_1_1123_0[1]));
    wire [1:0] far_1_1123_1;    relay_conn far_1_1123_1_a(.in(far_1_1123_0[0]), .out(far_1_1123_1[0]));    relay_conn far_1_1123_1_b(.in(far_1_1123_0[1]), .out(far_1_1123_1[1]));
    wire [1:0] far_1_1123_2;    relay_conn far_1_1123_2_a(.in(far_1_1123_1[0]), .out(far_1_1123_2[0]));    relay_conn far_1_1123_2_b(.in(far_1_1123_1[1]), .out(far_1_1123_2[1]));
    assign layer_1[103] = far_1_1123_2[0] & ~far_1_1123_2[1]; 
    wire [1:0] far_1_1124_0;    relay_conn far_1_1124_0_a(.in(layer_0[230]), .out(far_1_1124_0[0]));    relay_conn far_1_1124_0_b(.in(layer_0[193]), .out(far_1_1124_0[1]));
    assign layer_1[104] = far_1_1124_0[0]; 
    wire [1:0] far_1_1125_0;    relay_conn far_1_1125_0_a(.in(layer_0[117]), .out(far_1_1125_0[0]));    relay_conn far_1_1125_0_b(.in(layer_0[27]), .out(far_1_1125_0[1]));
    wire [1:0] far_1_1125_1;    relay_conn far_1_1125_1_a(.in(far_1_1125_0[0]), .out(far_1_1125_1[0]));    relay_conn far_1_1125_1_b(.in(far_1_1125_0[1]), .out(far_1_1125_1[1]));
    assign layer_1[105] = far_1_1125_1[0] | far_1_1125_1[1]; 
    wire [1:0] far_1_1126_0;    relay_conn far_1_1126_0_a(.in(layer_0[620]), .out(far_1_1126_0[0]));    relay_conn far_1_1126_0_b(.in(layer_0[540]), .out(far_1_1126_0[1]));
    wire [1:0] far_1_1126_1;    relay_conn far_1_1126_1_a(.in(far_1_1126_0[0]), .out(far_1_1126_1[0]));    relay_conn far_1_1126_1_b(.in(far_1_1126_0[1]), .out(far_1_1126_1[1]));
    assign layer_1[106] = ~far_1_1126_1[0] | (far_1_1126_1[0] & far_1_1126_1[1]); 
    wire [1:0] far_1_1127_0;    relay_conn far_1_1127_0_a(.in(layer_0[1002]), .out(far_1_1127_0[0]));    relay_conn far_1_1127_0_b(.in(layer_0[915]), .out(far_1_1127_0[1]));
    wire [1:0] far_1_1127_1;    relay_conn far_1_1127_1_a(.in(far_1_1127_0[0]), .out(far_1_1127_1[0]));    relay_conn far_1_1127_1_b(.in(far_1_1127_0[1]), .out(far_1_1127_1[1]));
    assign layer_1[107] = ~(far_1_1127_1[0] & far_1_1127_1[1]); 
    wire [1:0] far_1_1128_0;    relay_conn far_1_1128_0_a(.in(layer_0[338]), .out(far_1_1128_0[0]));    relay_conn far_1_1128_0_b(.in(layer_0[405]), .out(far_1_1128_0[1]));
    wire [1:0] far_1_1128_1;    relay_conn far_1_1128_1_a(.in(far_1_1128_0[0]), .out(far_1_1128_1[0]));    relay_conn far_1_1128_1_b(.in(far_1_1128_0[1]), .out(far_1_1128_1[1]));
    assign layer_1[108] = ~far_1_1128_1[1] | (far_1_1128_1[0] & far_1_1128_1[1]); 
    wire [1:0] far_1_1129_0;    relay_conn far_1_1129_0_a(.in(layer_0[475]), .out(far_1_1129_0[0]));    relay_conn far_1_1129_0_b(.in(layer_0[374]), .out(far_1_1129_0[1]));
    wire [1:0] far_1_1129_1;    relay_conn far_1_1129_1_a(.in(far_1_1129_0[0]), .out(far_1_1129_1[0]));    relay_conn far_1_1129_1_b(.in(far_1_1129_0[1]), .out(far_1_1129_1[1]));
    wire [1:0] far_1_1129_2;    relay_conn far_1_1129_2_a(.in(far_1_1129_1[0]), .out(far_1_1129_2[0]));    relay_conn far_1_1129_2_b(.in(far_1_1129_1[1]), .out(far_1_1129_2[1]));
    assign layer_1[109] = ~(far_1_1129_2[0] ^ far_1_1129_2[1]); 
    wire [1:0] far_1_1130_0;    relay_conn far_1_1130_0_a(.in(layer_0[463]), .out(far_1_1130_0[0]));    relay_conn far_1_1130_0_b(.in(layer_0[360]), .out(far_1_1130_0[1]));
    wire [1:0] far_1_1130_1;    relay_conn far_1_1130_1_a(.in(far_1_1130_0[0]), .out(far_1_1130_1[0]));    relay_conn far_1_1130_1_b(.in(far_1_1130_0[1]), .out(far_1_1130_1[1]));
    wire [1:0] far_1_1130_2;    relay_conn far_1_1130_2_a(.in(far_1_1130_1[0]), .out(far_1_1130_2[0]));    relay_conn far_1_1130_2_b(.in(far_1_1130_1[1]), .out(far_1_1130_2[1]));
    assign layer_1[110] = far_1_1130_2[0] & far_1_1130_2[1]; 
    wire [1:0] far_1_1131_0;    relay_conn far_1_1131_0_a(.in(layer_0[970]), .out(far_1_1131_0[0]));    relay_conn far_1_1131_0_b(.in(layer_0[915]), .out(far_1_1131_0[1]));
    assign layer_1[111] = ~far_1_1131_0[0]; 
    wire [1:0] far_1_1132_0;    relay_conn far_1_1132_0_a(.in(layer_0[681]), .out(far_1_1132_0[0]));    relay_conn far_1_1132_0_b(.in(layer_0[578]), .out(far_1_1132_0[1]));
    wire [1:0] far_1_1132_1;    relay_conn far_1_1132_1_a(.in(far_1_1132_0[0]), .out(far_1_1132_1[0]));    relay_conn far_1_1132_1_b(.in(far_1_1132_0[1]), .out(far_1_1132_1[1]));
    wire [1:0] far_1_1132_2;    relay_conn far_1_1132_2_a(.in(far_1_1132_1[0]), .out(far_1_1132_2[0]));    relay_conn far_1_1132_2_b(.in(far_1_1132_1[1]), .out(far_1_1132_2[1]));
    assign layer_1[112] = ~far_1_1132_2[1] | (far_1_1132_2[0] & far_1_1132_2[1]); 
    wire [1:0] far_1_1133_0;    relay_conn far_1_1133_0_a(.in(layer_0[158]), .out(far_1_1133_0[0]));    relay_conn far_1_1133_0_b(.in(layer_0[117]), .out(far_1_1133_0[1]));
    assign layer_1[113] = far_1_1133_0[0] & far_1_1133_0[1]; 
    wire [1:0] far_1_1134_0;    relay_conn far_1_1134_0_a(.in(layer_0[829]), .out(far_1_1134_0[0]));    relay_conn far_1_1134_0_b(.in(layer_0[762]), .out(far_1_1134_0[1]));
    wire [1:0] far_1_1134_1;    relay_conn far_1_1134_1_a(.in(far_1_1134_0[0]), .out(far_1_1134_1[0]));    relay_conn far_1_1134_1_b(.in(far_1_1134_0[1]), .out(far_1_1134_1[1]));
    assign layer_1[114] = ~far_1_1134_1[1] | (far_1_1134_1[0] & far_1_1134_1[1]); 
    wire [1:0] far_1_1135_0;    relay_conn far_1_1135_0_a(.in(layer_0[615]), .out(far_1_1135_0[0]));    relay_conn far_1_1135_0_b(.in(layer_0[723]), .out(far_1_1135_0[1]));
    wire [1:0] far_1_1135_1;    relay_conn far_1_1135_1_a(.in(far_1_1135_0[0]), .out(far_1_1135_1[0]));    relay_conn far_1_1135_1_b(.in(far_1_1135_0[1]), .out(far_1_1135_1[1]));
    wire [1:0] far_1_1135_2;    relay_conn far_1_1135_2_a(.in(far_1_1135_1[0]), .out(far_1_1135_2[0]));    relay_conn far_1_1135_2_b(.in(far_1_1135_1[1]), .out(far_1_1135_2[1]));
    assign layer_1[115] = far_1_1135_2[1]; 
    wire [1:0] far_1_1136_0;    relay_conn far_1_1136_0_a(.in(layer_0[607]), .out(far_1_1136_0[0]));    relay_conn far_1_1136_0_b(.in(layer_0[707]), .out(far_1_1136_0[1]));
    wire [1:0] far_1_1136_1;    relay_conn far_1_1136_1_a(.in(far_1_1136_0[0]), .out(far_1_1136_1[0]));    relay_conn far_1_1136_1_b(.in(far_1_1136_0[1]), .out(far_1_1136_1[1]));
    wire [1:0] far_1_1136_2;    relay_conn far_1_1136_2_a(.in(far_1_1136_1[0]), .out(far_1_1136_2[0]));    relay_conn far_1_1136_2_b(.in(far_1_1136_1[1]), .out(far_1_1136_2[1]));
    assign layer_1[116] = ~far_1_1136_2[0]; 
    wire [1:0] far_1_1137_0;    relay_conn far_1_1137_0_a(.in(layer_0[628]), .out(far_1_1137_0[0]));    relay_conn far_1_1137_0_b(.in(layer_0[514]), .out(far_1_1137_0[1]));
    wire [1:0] far_1_1137_1;    relay_conn far_1_1137_1_a(.in(far_1_1137_0[0]), .out(far_1_1137_1[0]));    relay_conn far_1_1137_1_b(.in(far_1_1137_0[1]), .out(far_1_1137_1[1]));
    wire [1:0] far_1_1137_2;    relay_conn far_1_1137_2_a(.in(far_1_1137_1[0]), .out(far_1_1137_2[0]));    relay_conn far_1_1137_2_b(.in(far_1_1137_1[1]), .out(far_1_1137_2[1]));
    assign layer_1[117] = far_1_1137_2[0]; 
    wire [1:0] far_1_1138_0;    relay_conn far_1_1138_0_a(.in(layer_0[560]), .out(far_1_1138_0[0]));    relay_conn far_1_1138_0_b(.in(layer_0[471]), .out(far_1_1138_0[1]));
    wire [1:0] far_1_1138_1;    relay_conn far_1_1138_1_a(.in(far_1_1138_0[0]), .out(far_1_1138_1[0]));    relay_conn far_1_1138_1_b(.in(far_1_1138_0[1]), .out(far_1_1138_1[1]));
    assign layer_1[118] = far_1_1138_1[0] & ~far_1_1138_1[1]; 
    wire [1:0] far_1_1139_0;    relay_conn far_1_1139_0_a(.in(layer_0[997]), .out(far_1_1139_0[0]));    relay_conn far_1_1139_0_b(.in(layer_0[914]), .out(far_1_1139_0[1]));
    wire [1:0] far_1_1139_1;    relay_conn far_1_1139_1_a(.in(far_1_1139_0[0]), .out(far_1_1139_1[0]));    relay_conn far_1_1139_1_b(.in(far_1_1139_0[1]), .out(far_1_1139_1[1]));
    assign layer_1[119] = far_1_1139_1[0] & ~far_1_1139_1[1]; 
    wire [1:0] far_1_1140_0;    relay_conn far_1_1140_0_a(.in(layer_0[367]), .out(far_1_1140_0[0]));    relay_conn far_1_1140_0_b(.in(layer_0[272]), .out(far_1_1140_0[1]));
    wire [1:0] far_1_1140_1;    relay_conn far_1_1140_1_a(.in(far_1_1140_0[0]), .out(far_1_1140_1[0]));    relay_conn far_1_1140_1_b(.in(far_1_1140_0[1]), .out(far_1_1140_1[1]));
    assign layer_1[120] = ~far_1_1140_1[0]; 
    wire [1:0] far_1_1141_0;    relay_conn far_1_1141_0_a(.in(layer_0[354]), .out(far_1_1141_0[0]));    relay_conn far_1_1141_0_b(.in(layer_0[397]), .out(far_1_1141_0[1]));
    assign layer_1[121] = far_1_1141_0[0] | far_1_1141_0[1]; 
    wire [1:0] far_1_1142_0;    relay_conn far_1_1142_0_a(.in(layer_0[2]), .out(far_1_1142_0[0]));    relay_conn far_1_1142_0_b(.in(layer_0[70]), .out(far_1_1142_0[1]));
    wire [1:0] far_1_1142_1;    relay_conn far_1_1142_1_a(.in(far_1_1142_0[0]), .out(far_1_1142_1[0]));    relay_conn far_1_1142_1_b(.in(far_1_1142_0[1]), .out(far_1_1142_1[1]));
    assign layer_1[122] = ~(far_1_1142_1[0] ^ far_1_1142_1[1]); 
    wire [1:0] far_1_1143_0;    relay_conn far_1_1143_0_a(.in(layer_0[316]), .out(far_1_1143_0[0]));    relay_conn far_1_1143_0_b(.in(layer_0[272]), .out(far_1_1143_0[1]));
    assign layer_1[123] = ~far_1_1143_0[1] | (far_1_1143_0[0] & far_1_1143_0[1]); 
    wire [1:0] far_1_1144_0;    relay_conn far_1_1144_0_a(.in(layer_0[1004]), .out(far_1_1144_0[0]));    relay_conn far_1_1144_0_b(.in(layer_0[938]), .out(far_1_1144_0[1]));
    wire [1:0] far_1_1144_1;    relay_conn far_1_1144_1_a(.in(far_1_1144_0[0]), .out(far_1_1144_1[0]));    relay_conn far_1_1144_1_b(.in(far_1_1144_0[1]), .out(far_1_1144_1[1]));
    assign layer_1[124] = far_1_1144_1[0] & far_1_1144_1[1]; 
    wire [1:0] far_1_1145_0;    relay_conn far_1_1145_0_a(.in(layer_0[821]), .out(far_1_1145_0[0]));    relay_conn far_1_1145_0_b(.in(layer_0[716]), .out(far_1_1145_0[1]));
    wire [1:0] far_1_1145_1;    relay_conn far_1_1145_1_a(.in(far_1_1145_0[0]), .out(far_1_1145_1[0]));    relay_conn far_1_1145_1_b(.in(far_1_1145_0[1]), .out(far_1_1145_1[1]));
    wire [1:0] far_1_1145_2;    relay_conn far_1_1145_2_a(.in(far_1_1145_1[0]), .out(far_1_1145_2[0]));    relay_conn far_1_1145_2_b(.in(far_1_1145_1[1]), .out(far_1_1145_2[1]));
    assign layer_1[125] = ~far_1_1145_2[1]; 
    wire [1:0] far_1_1146_0;    relay_conn far_1_1146_0_a(.in(layer_0[850]), .out(far_1_1146_0[0]));    relay_conn far_1_1146_0_b(.in(layer_0[915]), .out(far_1_1146_0[1]));
    wire [1:0] far_1_1146_1;    relay_conn far_1_1146_1_a(.in(far_1_1146_0[0]), .out(far_1_1146_1[0]));    relay_conn far_1_1146_1_b(.in(far_1_1146_0[1]), .out(far_1_1146_1[1]));
    assign layer_1[126] = ~(far_1_1146_1[0] | far_1_1146_1[1]); 
    assign layer_1[127] = ~layer_0[549] | (layer_0[549] & layer_0[580]); 
    assign layer_1[128] = layer_0[35] | layer_0[41]; 
    wire [1:0] far_1_1149_0;    relay_conn far_1_1149_0_a(.in(layer_0[218]), .out(far_1_1149_0[0]));    relay_conn far_1_1149_0_b(.in(layer_0[131]), .out(far_1_1149_0[1]));
    wire [1:0] far_1_1149_1;    relay_conn far_1_1149_1_a(.in(far_1_1149_0[0]), .out(far_1_1149_1[0]));    relay_conn far_1_1149_1_b(.in(far_1_1149_0[1]), .out(far_1_1149_1[1]));
    assign layer_1[129] = ~(far_1_1149_1[0] & far_1_1149_1[1]); 
    wire [1:0] far_1_1150_0;    relay_conn far_1_1150_0_a(.in(layer_0[789]), .out(far_1_1150_0[0]));    relay_conn far_1_1150_0_b(.in(layer_0[858]), .out(far_1_1150_0[1]));
    wire [1:0] far_1_1150_1;    relay_conn far_1_1150_1_a(.in(far_1_1150_0[0]), .out(far_1_1150_1[0]));    relay_conn far_1_1150_1_b(.in(far_1_1150_0[1]), .out(far_1_1150_1[1]));
    assign layer_1[130] = ~(far_1_1150_1[0] ^ far_1_1150_1[1]); 
    wire [1:0] far_1_1151_0;    relay_conn far_1_1151_0_a(.in(layer_0[353]), .out(far_1_1151_0[0]));    relay_conn far_1_1151_0_b(.in(layer_0[314]), .out(far_1_1151_0[1]));
    assign layer_1[131] = far_1_1151_0[1] & ~far_1_1151_0[0]; 
    assign layer_1[132] = ~(layer_0[46] | layer_0[57]); 
    wire [1:0] far_1_1153_0;    relay_conn far_1_1153_0_a(.in(layer_0[997]), .out(far_1_1153_0[0]));    relay_conn far_1_1153_0_b(.in(layer_0[915]), .out(far_1_1153_0[1]));
    wire [1:0] far_1_1153_1;    relay_conn far_1_1153_1_a(.in(far_1_1153_0[0]), .out(far_1_1153_1[0]));    relay_conn far_1_1153_1_b(.in(far_1_1153_0[1]), .out(far_1_1153_1[1]));
    assign layer_1[133] = ~far_1_1153_1[1] | (far_1_1153_1[0] & far_1_1153_1[1]); 
    assign layer_1[134] = ~(layer_0[795] ^ layer_0[816]); 
    assign layer_1[135] = layer_0[99] & ~layer_0[71]; 
    wire [1:0] far_1_1156_0;    relay_conn far_1_1156_0_a(.in(layer_0[151]), .out(far_1_1156_0[0]));    relay_conn far_1_1156_0_b(.in(layer_0[24]), .out(far_1_1156_0[1]));
    wire [1:0] far_1_1156_1;    relay_conn far_1_1156_1_a(.in(far_1_1156_0[0]), .out(far_1_1156_1[0]));    relay_conn far_1_1156_1_b(.in(far_1_1156_0[1]), .out(far_1_1156_1[1]));
    wire [1:0] far_1_1156_2;    relay_conn far_1_1156_2_a(.in(far_1_1156_1[0]), .out(far_1_1156_2[0]));    relay_conn far_1_1156_2_b(.in(far_1_1156_1[1]), .out(far_1_1156_2[1]));
    assign layer_1[136] = far_1_1156_2[0] | far_1_1156_2[1]; 
    wire [1:0] far_1_1157_0;    relay_conn far_1_1157_0_a(.in(layer_0[304]), .out(far_1_1157_0[0]));    relay_conn far_1_1157_0_b(.in(layer_0[261]), .out(far_1_1157_0[1]));
    assign layer_1[137] = ~far_1_1157_0[1]; 
    wire [1:0] far_1_1158_0;    relay_conn far_1_1158_0_a(.in(layer_0[23]), .out(far_1_1158_0[0]));    relay_conn far_1_1158_0_b(.in(layer_0[68]), .out(far_1_1158_0[1]));
    assign layer_1[138] = far_1_1158_0[0] & far_1_1158_0[1]; 
    assign layer_1[139] = layer_0[991]; 
    wire [1:0] far_1_1160_0;    relay_conn far_1_1160_0_a(.in(layer_0[824]), .out(far_1_1160_0[0]));    relay_conn far_1_1160_0_b(.in(layer_0[738]), .out(far_1_1160_0[1]));
    wire [1:0] far_1_1160_1;    relay_conn far_1_1160_1_a(.in(far_1_1160_0[0]), .out(far_1_1160_1[0]));    relay_conn far_1_1160_1_b(.in(far_1_1160_0[1]), .out(far_1_1160_1[1]));
    assign layer_1[140] = far_1_1160_1[0] & far_1_1160_1[1]; 
    assign layer_1[141] = ~(layer_0[696] & layer_0[723]); 
    wire [1:0] far_1_1162_0;    relay_conn far_1_1162_0_a(.in(layer_0[293]), .out(far_1_1162_0[0]));    relay_conn far_1_1162_0_b(.in(layer_0[395]), .out(far_1_1162_0[1]));
    wire [1:0] far_1_1162_1;    relay_conn far_1_1162_1_a(.in(far_1_1162_0[0]), .out(far_1_1162_1[0]));    relay_conn far_1_1162_1_b(.in(far_1_1162_0[1]), .out(far_1_1162_1[1]));
    wire [1:0] far_1_1162_2;    relay_conn far_1_1162_2_a(.in(far_1_1162_1[0]), .out(far_1_1162_2[0]));    relay_conn far_1_1162_2_b(.in(far_1_1162_1[1]), .out(far_1_1162_2[1]));
    assign layer_1[142] = far_1_1162_2[1] & ~far_1_1162_2[0]; 
    assign layer_1[143] = ~(layer_0[40] | layer_0[62]); 
    wire [1:0] far_1_1164_0;    relay_conn far_1_1164_0_a(.in(layer_0[868]), .out(far_1_1164_0[0]));    relay_conn far_1_1164_0_b(.in(layer_0[834]), .out(far_1_1164_0[1]));
    assign layer_1[144] = ~far_1_1164_0[1] | (far_1_1164_0[0] & far_1_1164_0[1]); 
    wire [1:0] far_1_1165_0;    relay_conn far_1_1165_0_a(.in(layer_0[199]), .out(far_1_1165_0[0]));    relay_conn far_1_1165_0_b(.in(layer_0[246]), .out(far_1_1165_0[1]));
    assign layer_1[145] = far_1_1165_0[1] & ~far_1_1165_0[0]; 
    wire [1:0] far_1_1166_0;    relay_conn far_1_1166_0_a(.in(layer_0[185]), .out(far_1_1166_0[0]));    relay_conn far_1_1166_0_b(.in(layer_0[272]), .out(far_1_1166_0[1]));
    wire [1:0] far_1_1166_1;    relay_conn far_1_1166_1_a(.in(far_1_1166_0[0]), .out(far_1_1166_1[0]));    relay_conn far_1_1166_1_b(.in(far_1_1166_0[1]), .out(far_1_1166_1[1]));
    assign layer_1[146] = ~far_1_1166_1[1]; 
    assign layer_1[147] = layer_0[265]; 
    wire [1:0] far_1_1168_0;    relay_conn far_1_1168_0_a(.in(layer_0[546]), .out(far_1_1168_0[0]));    relay_conn far_1_1168_0_b(.in(layer_0[476]), .out(far_1_1168_0[1]));
    wire [1:0] far_1_1168_1;    relay_conn far_1_1168_1_a(.in(far_1_1168_0[0]), .out(far_1_1168_1[0]));    relay_conn far_1_1168_1_b(.in(far_1_1168_0[1]), .out(far_1_1168_1[1]));
    assign layer_1[148] = ~(far_1_1168_1[0] ^ far_1_1168_1[1]); 
    wire [1:0] far_1_1169_0;    relay_conn far_1_1169_0_a(.in(layer_0[327]), .out(far_1_1169_0[0]));    relay_conn far_1_1169_0_b(.in(layer_0[422]), .out(far_1_1169_0[1]));
    wire [1:0] far_1_1169_1;    relay_conn far_1_1169_1_a(.in(far_1_1169_0[0]), .out(far_1_1169_1[0]));    relay_conn far_1_1169_1_b(.in(far_1_1169_0[1]), .out(far_1_1169_1[1]));
    assign layer_1[149] = far_1_1169_1[1]; 
    wire [1:0] far_1_1170_0;    relay_conn far_1_1170_0_a(.in(layer_0[19]), .out(far_1_1170_0[0]));    relay_conn far_1_1170_0_b(.in(layer_0[140]), .out(far_1_1170_0[1]));
    wire [1:0] far_1_1170_1;    relay_conn far_1_1170_1_a(.in(far_1_1170_0[0]), .out(far_1_1170_1[0]));    relay_conn far_1_1170_1_b(.in(far_1_1170_0[1]), .out(far_1_1170_1[1]));
    wire [1:0] far_1_1170_2;    relay_conn far_1_1170_2_a(.in(far_1_1170_1[0]), .out(far_1_1170_2[0]));    relay_conn far_1_1170_2_b(.in(far_1_1170_1[1]), .out(far_1_1170_2[1]));
    assign layer_1[150] = ~(far_1_1170_2[0] ^ far_1_1170_2[1]); 
    wire [1:0] far_1_1171_0;    relay_conn far_1_1171_0_a(.in(layer_0[287]), .out(far_1_1171_0[0]));    relay_conn far_1_1171_0_b(.in(layer_0[404]), .out(far_1_1171_0[1]));
    wire [1:0] far_1_1171_1;    relay_conn far_1_1171_1_a(.in(far_1_1171_0[0]), .out(far_1_1171_1[0]));    relay_conn far_1_1171_1_b(.in(far_1_1171_0[1]), .out(far_1_1171_1[1]));
    wire [1:0] far_1_1171_2;    relay_conn far_1_1171_2_a(.in(far_1_1171_1[0]), .out(far_1_1171_2[0]));    relay_conn far_1_1171_2_b(.in(far_1_1171_1[1]), .out(far_1_1171_2[1]));
    assign layer_1[151] = far_1_1171_2[0] | far_1_1171_2[1]; 
    wire [1:0] far_1_1172_0;    relay_conn far_1_1172_0_a(.in(layer_0[607]), .out(far_1_1172_0[0]));    relay_conn far_1_1172_0_b(.in(layer_0[735]), .out(far_1_1172_0[1]));
    wire [1:0] far_1_1172_1;    relay_conn far_1_1172_1_a(.in(far_1_1172_0[0]), .out(far_1_1172_1[0]));    relay_conn far_1_1172_1_b(.in(far_1_1172_0[1]), .out(far_1_1172_1[1]));
    wire [1:0] far_1_1172_2;    relay_conn far_1_1172_2_a(.in(far_1_1172_1[0]), .out(far_1_1172_2[0]));    relay_conn far_1_1172_2_b(.in(far_1_1172_1[1]), .out(far_1_1172_2[1]));
    wire [1:0] far_1_1172_3;    relay_conn far_1_1172_3_a(.in(far_1_1172_2[0]), .out(far_1_1172_3[0]));    relay_conn far_1_1172_3_b(.in(far_1_1172_2[1]), .out(far_1_1172_3[1]));
    assign layer_1[152] = ~(far_1_1172_3[0] ^ far_1_1172_3[1]); 
    wire [1:0] far_1_1173_0;    relay_conn far_1_1173_0_a(.in(layer_0[35]), .out(far_1_1173_0[0]));    relay_conn far_1_1173_0_b(.in(layer_0[148]), .out(far_1_1173_0[1]));
    wire [1:0] far_1_1173_1;    relay_conn far_1_1173_1_a(.in(far_1_1173_0[0]), .out(far_1_1173_1[0]));    relay_conn far_1_1173_1_b(.in(far_1_1173_0[1]), .out(far_1_1173_1[1]));
    wire [1:0] far_1_1173_2;    relay_conn far_1_1173_2_a(.in(far_1_1173_1[0]), .out(far_1_1173_2[0]));    relay_conn far_1_1173_2_b(.in(far_1_1173_1[1]), .out(far_1_1173_2[1]));
    assign layer_1[153] = far_1_1173_2[1]; 
    wire [1:0] far_1_1174_0;    relay_conn far_1_1174_0_a(.in(layer_0[55]), .out(far_1_1174_0[0]));    relay_conn far_1_1174_0_b(.in(layer_0[177]), .out(far_1_1174_0[1]));
    wire [1:0] far_1_1174_1;    relay_conn far_1_1174_1_a(.in(far_1_1174_0[0]), .out(far_1_1174_1[0]));    relay_conn far_1_1174_1_b(.in(far_1_1174_0[1]), .out(far_1_1174_1[1]));
    wire [1:0] far_1_1174_2;    relay_conn far_1_1174_2_a(.in(far_1_1174_1[0]), .out(far_1_1174_2[0]));    relay_conn far_1_1174_2_b(.in(far_1_1174_1[1]), .out(far_1_1174_2[1]));
    assign layer_1[154] = far_1_1174_2[0] & far_1_1174_2[1]; 
    assign layer_1[155] = ~layer_0[580]; 
    wire [1:0] far_1_1176_0;    relay_conn far_1_1176_0_a(.in(layer_0[73]), .out(far_1_1176_0[0]));    relay_conn far_1_1176_0_b(.in(layer_0[148]), .out(far_1_1176_0[1]));
    wire [1:0] far_1_1176_1;    relay_conn far_1_1176_1_a(.in(far_1_1176_0[0]), .out(far_1_1176_1[0]));    relay_conn far_1_1176_1_b(.in(far_1_1176_0[1]), .out(far_1_1176_1[1]));
    assign layer_1[156] = far_1_1176_1[0] ^ far_1_1176_1[1]; 
    wire [1:0] far_1_1177_0;    relay_conn far_1_1177_0_a(.in(layer_0[272]), .out(far_1_1177_0[0]));    relay_conn far_1_1177_0_b(.in(layer_0[216]), .out(far_1_1177_0[1]));
    assign layer_1[157] = far_1_1177_0[0]; 
    wire [1:0] far_1_1178_0;    relay_conn far_1_1178_0_a(.in(layer_0[635]), .out(far_1_1178_0[0]));    relay_conn far_1_1178_0_b(.in(layer_0[579]), .out(far_1_1178_0[1]));
    assign layer_1[158] = far_1_1178_0[0]; 
    assign layer_1[159] = ~layer_0[377] | (layer_0[377] & layer_0[379]); 
    wire [1:0] far_1_1180_0;    relay_conn far_1_1180_0_a(.in(layer_0[391]), .out(far_1_1180_0[0]));    relay_conn far_1_1180_0_b(.in(layer_0[441]), .out(far_1_1180_0[1]));
    assign layer_1[160] = ~(far_1_1180_0[0] & far_1_1180_0[1]); 
    assign layer_1[161] = ~layer_0[377]; 
    wire [1:0] far_1_1182_0;    relay_conn far_1_1182_0_a(.in(layer_0[459]), .out(far_1_1182_0[0]));    relay_conn far_1_1182_0_b(.in(layer_0[411]), .out(far_1_1182_0[1]));
    assign layer_1[162] = far_1_1182_0[0] & ~far_1_1182_0[1]; 
    wire [1:0] far_1_1183_0;    relay_conn far_1_1183_0_a(.in(layer_0[252]), .out(far_1_1183_0[0]));    relay_conn far_1_1183_0_b(.in(layer_0[349]), .out(far_1_1183_0[1]));
    wire [1:0] far_1_1183_1;    relay_conn far_1_1183_1_a(.in(far_1_1183_0[0]), .out(far_1_1183_1[0]));    relay_conn far_1_1183_1_b(.in(far_1_1183_0[1]), .out(far_1_1183_1[1]));
    wire [1:0] far_1_1183_2;    relay_conn far_1_1183_2_a(.in(far_1_1183_1[0]), .out(far_1_1183_2[0]));    relay_conn far_1_1183_2_b(.in(far_1_1183_1[1]), .out(far_1_1183_2[1]));
    assign layer_1[163] = ~far_1_1183_2[0] | (far_1_1183_2[0] & far_1_1183_2[1]); 
    wire [1:0] far_1_1184_0;    relay_conn far_1_1184_0_a(.in(layer_0[710]), .out(far_1_1184_0[0]));    relay_conn far_1_1184_0_b(.in(layer_0[678]), .out(far_1_1184_0[1]));
    assign layer_1[164] = ~far_1_1184_0[0] | (far_1_1184_0[0] & far_1_1184_0[1]); 
    wire [1:0] far_1_1185_0;    relay_conn far_1_1185_0_a(.in(layer_0[467]), .out(far_1_1185_0[0]));    relay_conn far_1_1185_0_b(.in(layer_0[432]), .out(far_1_1185_0[1]));
    assign layer_1[165] = ~far_1_1185_0[0]; 
    wire [1:0] far_1_1186_0;    relay_conn far_1_1186_0_a(.in(layer_0[810]), .out(far_1_1186_0[0]));    relay_conn far_1_1186_0_b(.in(layer_0[884]), .out(far_1_1186_0[1]));
    wire [1:0] far_1_1186_1;    relay_conn far_1_1186_1_a(.in(far_1_1186_0[0]), .out(far_1_1186_1[0]));    relay_conn far_1_1186_1_b(.in(far_1_1186_0[1]), .out(far_1_1186_1[1]));
    assign layer_1[166] = far_1_1186_1[1] & ~far_1_1186_1[0]; 
    wire [1:0] far_1_1187_0;    relay_conn far_1_1187_0_a(.in(layer_0[319]), .out(far_1_1187_0[0]));    relay_conn far_1_1187_0_b(.in(layer_0[377]), .out(far_1_1187_0[1]));
    assign layer_1[167] = far_1_1187_0[0] & ~far_1_1187_0[1]; 
    wire [1:0] far_1_1188_0;    relay_conn far_1_1188_0_a(.in(layer_0[261]), .out(far_1_1188_0[0]));    relay_conn far_1_1188_0_b(.in(layer_0[310]), .out(far_1_1188_0[1]));
    assign layer_1[168] = ~(far_1_1188_0[0] & far_1_1188_0[1]); 
    wire [1:0] far_1_1189_0;    relay_conn far_1_1189_0_a(.in(layer_0[71]), .out(far_1_1189_0[0]));    relay_conn far_1_1189_0_b(.in(layer_0[108]), .out(far_1_1189_0[1]));
    assign layer_1[169] = far_1_1189_0[1]; 
    assign layer_1[170] = layer_0[949]; 
    wire [1:0] far_1_1191_0;    relay_conn far_1_1191_0_a(.in(layer_0[360]), .out(far_1_1191_0[0]));    relay_conn far_1_1191_0_b(.in(layer_0[297]), .out(far_1_1191_0[1]));
    assign layer_1[171] = ~far_1_1191_0[1] | (far_1_1191_0[0] & far_1_1191_0[1]); 
    wire [1:0] far_1_1192_0;    relay_conn far_1_1192_0_a(.in(layer_0[116]), .out(far_1_1192_0[0]));    relay_conn far_1_1192_0_b(.in(layer_0[57]), .out(far_1_1192_0[1]));
    assign layer_1[172] = ~far_1_1192_0[0]; 
    wire [1:0] far_1_1193_0;    relay_conn far_1_1193_0_a(.in(layer_0[173]), .out(far_1_1193_0[0]));    relay_conn far_1_1193_0_b(.in(layer_0[218]), .out(far_1_1193_0[1]));
    assign layer_1[173] = far_1_1193_0[0] ^ far_1_1193_0[1]; 
    wire [1:0] far_1_1194_0;    relay_conn far_1_1194_0_a(.in(layer_0[638]), .out(far_1_1194_0[0]));    relay_conn far_1_1194_0_b(.in(layer_0[696]), .out(far_1_1194_0[1]));
    assign layer_1[174] = far_1_1194_0[0] & far_1_1194_0[1]; 
    wire [1:0] far_1_1195_0;    relay_conn far_1_1195_0_a(.in(layer_0[961]), .out(far_1_1195_0[0]));    relay_conn far_1_1195_0_b(.in(layer_0[891]), .out(far_1_1195_0[1]));
    wire [1:0] far_1_1195_1;    relay_conn far_1_1195_1_a(.in(far_1_1195_0[0]), .out(far_1_1195_1[0]));    relay_conn far_1_1195_1_b(.in(far_1_1195_0[1]), .out(far_1_1195_1[1]));
    assign layer_1[175] = far_1_1195_1[0]; 
    wire [1:0] far_1_1196_0;    relay_conn far_1_1196_0_a(.in(layer_0[310]), .out(far_1_1196_0[0]));    relay_conn far_1_1196_0_b(.in(layer_0[194]), .out(far_1_1196_0[1]));
    wire [1:0] far_1_1196_1;    relay_conn far_1_1196_1_a(.in(far_1_1196_0[0]), .out(far_1_1196_1[0]));    relay_conn far_1_1196_1_b(.in(far_1_1196_0[1]), .out(far_1_1196_1[1]));
    wire [1:0] far_1_1196_2;    relay_conn far_1_1196_2_a(.in(far_1_1196_1[0]), .out(far_1_1196_2[0]));    relay_conn far_1_1196_2_b(.in(far_1_1196_1[1]), .out(far_1_1196_2[1]));
    assign layer_1[176] = far_1_1196_2[0] | far_1_1196_2[1]; 
    wire [1:0] far_1_1197_0;    relay_conn far_1_1197_0_a(.in(layer_0[909]), .out(far_1_1197_0[0]));    relay_conn far_1_1197_0_b(.in(layer_0[954]), .out(far_1_1197_0[1]));
    assign layer_1[177] = far_1_1197_0[1] & ~far_1_1197_0[0]; 
    assign layer_1[178] = layer_0[580] & ~layer_0[607]; 
    wire [1:0] far_1_1199_0;    relay_conn far_1_1199_0_a(.in(layer_0[400]), .out(far_1_1199_0[0]));    relay_conn far_1_1199_0_b(.in(layer_0[494]), .out(far_1_1199_0[1]));
    wire [1:0] far_1_1199_1;    relay_conn far_1_1199_1_a(.in(far_1_1199_0[0]), .out(far_1_1199_1[0]));    relay_conn far_1_1199_1_b(.in(far_1_1199_0[1]), .out(far_1_1199_1[1]));
    assign layer_1[179] = far_1_1199_1[1] & ~far_1_1199_1[0]; 
    wire [1:0] far_1_1200_0;    relay_conn far_1_1200_0_a(.in(layer_0[352]), .out(far_1_1200_0[0]));    relay_conn far_1_1200_0_b(.in(layer_0[253]), .out(far_1_1200_0[1]));
    wire [1:0] far_1_1200_1;    relay_conn far_1_1200_1_a(.in(far_1_1200_0[0]), .out(far_1_1200_1[0]));    relay_conn far_1_1200_1_b(.in(far_1_1200_0[1]), .out(far_1_1200_1[1]));
    wire [1:0] far_1_1200_2;    relay_conn far_1_1200_2_a(.in(far_1_1200_1[0]), .out(far_1_1200_2[0]));    relay_conn far_1_1200_2_b(.in(far_1_1200_1[1]), .out(far_1_1200_2[1]));
    assign layer_1[180] = far_1_1200_2[0] & ~far_1_1200_2[1]; 
    wire [1:0] far_1_1201_0;    relay_conn far_1_1201_0_a(.in(layer_0[341]), .out(far_1_1201_0[0]));    relay_conn far_1_1201_0_b(.in(layer_0[448]), .out(far_1_1201_0[1]));
    wire [1:0] far_1_1201_1;    relay_conn far_1_1201_1_a(.in(far_1_1201_0[0]), .out(far_1_1201_1[0]));    relay_conn far_1_1201_1_b(.in(far_1_1201_0[1]), .out(far_1_1201_1[1]));
    wire [1:0] far_1_1201_2;    relay_conn far_1_1201_2_a(.in(far_1_1201_1[0]), .out(far_1_1201_2[0]));    relay_conn far_1_1201_2_b(.in(far_1_1201_1[1]), .out(far_1_1201_2[1]));
    assign layer_1[181] = far_1_1201_2[1] & ~far_1_1201_2[0]; 
    wire [1:0] far_1_1202_0;    relay_conn far_1_1202_0_a(.in(layer_0[204]), .out(far_1_1202_0[0]));    relay_conn far_1_1202_0_b(.in(layer_0[253]), .out(far_1_1202_0[1]));
    assign layer_1[182] = ~(far_1_1202_0[0] & far_1_1202_0[1]); 
    wire [1:0] far_1_1203_0;    relay_conn far_1_1203_0_a(.in(layer_0[57]), .out(far_1_1203_0[0]));    relay_conn far_1_1203_0_b(.in(layer_0[121]), .out(far_1_1203_0[1]));
    wire [1:0] far_1_1203_1;    relay_conn far_1_1203_1_a(.in(far_1_1203_0[0]), .out(far_1_1203_1[0]));    relay_conn far_1_1203_1_b(.in(far_1_1203_0[1]), .out(far_1_1203_1[1]));
    assign layer_1[183] = far_1_1203_1[0] | far_1_1203_1[1]; 
    wire [1:0] far_1_1204_0;    relay_conn far_1_1204_0_a(.in(layer_0[625]), .out(far_1_1204_0[0]));    relay_conn far_1_1204_0_b(.in(layer_0[748]), .out(far_1_1204_0[1]));
    wire [1:0] far_1_1204_1;    relay_conn far_1_1204_1_a(.in(far_1_1204_0[0]), .out(far_1_1204_1[0]));    relay_conn far_1_1204_1_b(.in(far_1_1204_0[1]), .out(far_1_1204_1[1]));
    wire [1:0] far_1_1204_2;    relay_conn far_1_1204_2_a(.in(far_1_1204_1[0]), .out(far_1_1204_2[0]));    relay_conn far_1_1204_2_b(.in(far_1_1204_1[1]), .out(far_1_1204_2[1]));
    assign layer_1[184] = far_1_1204_2[0] & far_1_1204_2[1]; 
    wire [1:0] far_1_1205_0;    relay_conn far_1_1205_0_a(.in(layer_0[867]), .out(far_1_1205_0[0]));    relay_conn far_1_1205_0_b(.in(layer_0[748]), .out(far_1_1205_0[1]));
    wire [1:0] far_1_1205_1;    relay_conn far_1_1205_1_a(.in(far_1_1205_0[0]), .out(far_1_1205_1[0]));    relay_conn far_1_1205_1_b(.in(far_1_1205_0[1]), .out(far_1_1205_1[1]));
    wire [1:0] far_1_1205_2;    relay_conn far_1_1205_2_a(.in(far_1_1205_1[0]), .out(far_1_1205_2[0]));    relay_conn far_1_1205_2_b(.in(far_1_1205_1[1]), .out(far_1_1205_2[1]));
    assign layer_1[185] = ~far_1_1205_2[1] | (far_1_1205_2[0] & far_1_1205_2[1]); 
    wire [1:0] far_1_1206_0;    relay_conn far_1_1206_0_a(.in(layer_0[997]), .out(far_1_1206_0[0]));    relay_conn far_1_1206_0_b(.in(layer_0[909]), .out(far_1_1206_0[1]));
    wire [1:0] far_1_1206_1;    relay_conn far_1_1206_1_a(.in(far_1_1206_0[0]), .out(far_1_1206_1[0]));    relay_conn far_1_1206_1_b(.in(far_1_1206_0[1]), .out(far_1_1206_1[1]));
    assign layer_1[186] = ~far_1_1206_1[0]; 
    wire [1:0] far_1_1207_0;    relay_conn far_1_1207_0_a(.in(layer_0[185]), .out(far_1_1207_0[0]));    relay_conn far_1_1207_0_b(.in(layer_0[271]), .out(far_1_1207_0[1]));
    wire [1:0] far_1_1207_1;    relay_conn far_1_1207_1_a(.in(far_1_1207_0[0]), .out(far_1_1207_1[0]));    relay_conn far_1_1207_1_b(.in(far_1_1207_0[1]), .out(far_1_1207_1[1]));
    assign layer_1[187] = far_1_1207_1[0] & ~far_1_1207_1[1]; 
    wire [1:0] far_1_1208_0;    relay_conn far_1_1208_0_a(.in(layer_0[456]), .out(far_1_1208_0[0]));    relay_conn far_1_1208_0_b(.in(layer_0[336]), .out(far_1_1208_0[1]));
    wire [1:0] far_1_1208_1;    relay_conn far_1_1208_1_a(.in(far_1_1208_0[0]), .out(far_1_1208_1[0]));    relay_conn far_1_1208_1_b(.in(far_1_1208_0[1]), .out(far_1_1208_1[1]));
    wire [1:0] far_1_1208_2;    relay_conn far_1_1208_2_a(.in(far_1_1208_1[0]), .out(far_1_1208_2[0]));    relay_conn far_1_1208_2_b(.in(far_1_1208_1[1]), .out(far_1_1208_2[1]));
    assign layer_1[188] = far_1_1208_2[0] & ~far_1_1208_2[1]; 
    assign layer_1[189] = ~(layer_0[485] | layer_0[489]); 
    wire [1:0] far_1_1210_0;    relay_conn far_1_1210_0_a(.in(layer_0[902]), .out(far_1_1210_0[0]));    relay_conn far_1_1210_0_b(.in(layer_0[808]), .out(far_1_1210_0[1]));
    wire [1:0] far_1_1210_1;    relay_conn far_1_1210_1_a(.in(far_1_1210_0[0]), .out(far_1_1210_1[0]));    relay_conn far_1_1210_1_b(.in(far_1_1210_0[1]), .out(far_1_1210_1[1]));
    assign layer_1[190] = far_1_1210_1[1]; 
    wire [1:0] far_1_1211_0;    relay_conn far_1_1211_0_a(.in(layer_0[676]), .out(far_1_1211_0[0]));    relay_conn far_1_1211_0_b(.in(layer_0[773]), .out(far_1_1211_0[1]));
    wire [1:0] far_1_1211_1;    relay_conn far_1_1211_1_a(.in(far_1_1211_0[0]), .out(far_1_1211_1[0]));    relay_conn far_1_1211_1_b(.in(far_1_1211_0[1]), .out(far_1_1211_1[1]));
    wire [1:0] far_1_1211_2;    relay_conn far_1_1211_2_a(.in(far_1_1211_1[0]), .out(far_1_1211_2[0]));    relay_conn far_1_1211_2_b(.in(far_1_1211_1[1]), .out(far_1_1211_2[1]));
    assign layer_1[191] = ~far_1_1211_2[1]; 
    wire [1:0] far_1_1212_0;    relay_conn far_1_1212_0_a(.in(layer_0[626]), .out(far_1_1212_0[0]));    relay_conn far_1_1212_0_b(.in(layer_0[704]), .out(far_1_1212_0[1]));
    wire [1:0] far_1_1212_1;    relay_conn far_1_1212_1_a(.in(far_1_1212_0[0]), .out(far_1_1212_1[0]));    relay_conn far_1_1212_1_b(.in(far_1_1212_0[1]), .out(far_1_1212_1[1]));
    assign layer_1[192] = ~(far_1_1212_1[0] & far_1_1212_1[1]); 
    wire [1:0] far_1_1213_0;    relay_conn far_1_1213_0_a(.in(layer_0[9]), .out(far_1_1213_0[0]));    relay_conn far_1_1213_0_b(.in(layer_0[56]), .out(far_1_1213_0[1]));
    assign layer_1[193] = far_1_1213_0[0] | far_1_1213_0[1]; 
    wire [1:0] far_1_1214_0;    relay_conn far_1_1214_0_a(.in(layer_0[431]), .out(far_1_1214_0[0]));    relay_conn far_1_1214_0_b(.in(layer_0[339]), .out(far_1_1214_0[1]));
    wire [1:0] far_1_1214_1;    relay_conn far_1_1214_1_a(.in(far_1_1214_0[0]), .out(far_1_1214_1[0]));    relay_conn far_1_1214_1_b(.in(far_1_1214_0[1]), .out(far_1_1214_1[1]));
    assign layer_1[194] = ~(far_1_1214_1[0] | far_1_1214_1[1]); 
    wire [1:0] far_1_1215_0;    relay_conn far_1_1215_0_a(.in(layer_0[386]), .out(far_1_1215_0[0]));    relay_conn far_1_1215_0_b(.in(layer_0[261]), .out(far_1_1215_0[1]));
    wire [1:0] far_1_1215_1;    relay_conn far_1_1215_1_a(.in(far_1_1215_0[0]), .out(far_1_1215_1[0]));    relay_conn far_1_1215_1_b(.in(far_1_1215_0[1]), .out(far_1_1215_1[1]));
    wire [1:0] far_1_1215_2;    relay_conn far_1_1215_2_a(.in(far_1_1215_1[0]), .out(far_1_1215_2[0]));    relay_conn far_1_1215_2_b(.in(far_1_1215_1[1]), .out(far_1_1215_2[1]));
    assign layer_1[195] = ~far_1_1215_2[1] | (far_1_1215_2[0] & far_1_1215_2[1]); 
    assign layer_1[196] = layer_0[638]; 
    wire [1:0] far_1_1217_0;    relay_conn far_1_1217_0_a(.in(layer_0[277]), .out(far_1_1217_0[0]));    relay_conn far_1_1217_0_b(.in(layer_0[152]), .out(far_1_1217_0[1]));
    wire [1:0] far_1_1217_1;    relay_conn far_1_1217_1_a(.in(far_1_1217_0[0]), .out(far_1_1217_1[0]));    relay_conn far_1_1217_1_b(.in(far_1_1217_0[1]), .out(far_1_1217_1[1]));
    wire [1:0] far_1_1217_2;    relay_conn far_1_1217_2_a(.in(far_1_1217_1[0]), .out(far_1_1217_2[0]));    relay_conn far_1_1217_2_b(.in(far_1_1217_1[1]), .out(far_1_1217_2[1]));
    assign layer_1[197] = far_1_1217_2[0] ^ far_1_1217_2[1]; 
    wire [1:0] far_1_1218_0;    relay_conn far_1_1218_0_a(.in(layer_0[841]), .out(far_1_1218_0[0]));    relay_conn far_1_1218_0_b(.in(layer_0[894]), .out(far_1_1218_0[1]));
    assign layer_1[198] = far_1_1218_0[0] ^ far_1_1218_0[1]; 
    assign layer_1[199] = layer_0[512] & layer_0[484]; 
    wire [1:0] far_1_1220_0;    relay_conn far_1_1220_0_a(.in(layer_0[559]), .out(far_1_1220_0[0]));    relay_conn far_1_1220_0_b(.in(layer_0[661]), .out(far_1_1220_0[1]));
    wire [1:0] far_1_1220_1;    relay_conn far_1_1220_1_a(.in(far_1_1220_0[0]), .out(far_1_1220_1[0]));    relay_conn far_1_1220_1_b(.in(far_1_1220_0[1]), .out(far_1_1220_1[1]));
    wire [1:0] far_1_1220_2;    relay_conn far_1_1220_2_a(.in(far_1_1220_1[0]), .out(far_1_1220_2[0]));    relay_conn far_1_1220_2_b(.in(far_1_1220_1[1]), .out(far_1_1220_2[1]));
    assign layer_1[200] = ~(far_1_1220_2[0] & far_1_1220_2[1]); 
    wire [1:0] far_1_1221_0;    relay_conn far_1_1221_0_a(.in(layer_0[365]), .out(far_1_1221_0[0]));    relay_conn far_1_1221_0_b(.in(layer_0[419]), .out(far_1_1221_0[1]));
    assign layer_1[201] = ~(far_1_1221_0[0] ^ far_1_1221_0[1]); 
    wire [1:0] far_1_1222_0;    relay_conn far_1_1222_0_a(.in(layer_0[443]), .out(far_1_1222_0[0]));    relay_conn far_1_1222_0_b(.in(layer_0[319]), .out(far_1_1222_0[1]));
    wire [1:0] far_1_1222_1;    relay_conn far_1_1222_1_a(.in(far_1_1222_0[0]), .out(far_1_1222_1[0]));    relay_conn far_1_1222_1_b(.in(far_1_1222_0[1]), .out(far_1_1222_1[1]));
    wire [1:0] far_1_1222_2;    relay_conn far_1_1222_2_a(.in(far_1_1222_1[0]), .out(far_1_1222_2[0]));    relay_conn far_1_1222_2_b(.in(far_1_1222_1[1]), .out(far_1_1222_2[1]));
    assign layer_1[202] = far_1_1222_2[0] | far_1_1222_2[1]; 
    wire [1:0] far_1_1223_0;    relay_conn far_1_1223_0_a(.in(layer_0[506]), .out(far_1_1223_0[0]));    relay_conn far_1_1223_0_b(.in(layer_0[621]), .out(far_1_1223_0[1]));
    wire [1:0] far_1_1223_1;    relay_conn far_1_1223_1_a(.in(far_1_1223_0[0]), .out(far_1_1223_1[0]));    relay_conn far_1_1223_1_b(.in(far_1_1223_0[1]), .out(far_1_1223_1[1]));
    wire [1:0] far_1_1223_2;    relay_conn far_1_1223_2_a(.in(far_1_1223_1[0]), .out(far_1_1223_2[0]));    relay_conn far_1_1223_2_b(.in(far_1_1223_1[1]), .out(far_1_1223_2[1]));
    assign layer_1[203] = far_1_1223_2[0] ^ far_1_1223_2[1]; 
    wire [1:0] far_1_1224_0;    relay_conn far_1_1224_0_a(.in(layer_0[711]), .out(far_1_1224_0[0]));    relay_conn far_1_1224_0_b(.in(layer_0[835]), .out(far_1_1224_0[1]));
    wire [1:0] far_1_1224_1;    relay_conn far_1_1224_1_a(.in(far_1_1224_0[0]), .out(far_1_1224_1[0]));    relay_conn far_1_1224_1_b(.in(far_1_1224_0[1]), .out(far_1_1224_1[1]));
    wire [1:0] far_1_1224_2;    relay_conn far_1_1224_2_a(.in(far_1_1224_1[0]), .out(far_1_1224_2[0]));    relay_conn far_1_1224_2_b(.in(far_1_1224_1[1]), .out(far_1_1224_2[1]));
    assign layer_1[204] = far_1_1224_2[0]; 
    wire [1:0] far_1_1225_0;    relay_conn far_1_1225_0_a(.in(layer_0[38]), .out(far_1_1225_0[0]));    relay_conn far_1_1225_0_b(.in(layer_0[111]), .out(far_1_1225_0[1]));
    wire [1:0] far_1_1225_1;    relay_conn far_1_1225_1_a(.in(far_1_1225_0[0]), .out(far_1_1225_1[0]));    relay_conn far_1_1225_1_b(.in(far_1_1225_0[1]), .out(far_1_1225_1[1]));
    assign layer_1[205] = far_1_1225_1[1]; 
    wire [1:0] far_1_1226_0;    relay_conn far_1_1226_0_a(.in(layer_0[0]), .out(far_1_1226_0[0]));    relay_conn far_1_1226_0_b(.in(layer_0[66]), .out(far_1_1226_0[1]));
    wire [1:0] far_1_1226_1;    relay_conn far_1_1226_1_a(.in(far_1_1226_0[0]), .out(far_1_1226_1[0]));    relay_conn far_1_1226_1_b(.in(far_1_1226_0[1]), .out(far_1_1226_1[1]));
    assign layer_1[206] = ~far_1_1226_1[1] | (far_1_1226_1[0] & far_1_1226_1[1]); 
    wire [1:0] far_1_1227_0;    relay_conn far_1_1227_0_a(.in(layer_0[438]), .out(far_1_1227_0[0]));    relay_conn far_1_1227_0_b(.in(layer_0[544]), .out(far_1_1227_0[1]));
    wire [1:0] far_1_1227_1;    relay_conn far_1_1227_1_a(.in(far_1_1227_0[0]), .out(far_1_1227_1[0]));    relay_conn far_1_1227_1_b(.in(far_1_1227_0[1]), .out(far_1_1227_1[1]));
    wire [1:0] far_1_1227_2;    relay_conn far_1_1227_2_a(.in(far_1_1227_1[0]), .out(far_1_1227_2[0]));    relay_conn far_1_1227_2_b(.in(far_1_1227_1[1]), .out(far_1_1227_2[1]));
    assign layer_1[207] = ~far_1_1227_2[0] | (far_1_1227_2[0] & far_1_1227_2[1]); 
    wire [1:0] far_1_1228_0;    relay_conn far_1_1228_0_a(.in(layer_0[659]), .out(far_1_1228_0[0]));    relay_conn far_1_1228_0_b(.in(layer_0[600]), .out(far_1_1228_0[1]));
    assign layer_1[208] = ~far_1_1228_0[1] | (far_1_1228_0[0] & far_1_1228_0[1]); 
    wire [1:0] far_1_1229_0;    relay_conn far_1_1229_0_a(.in(layer_0[713]), .out(far_1_1229_0[0]));    relay_conn far_1_1229_0_b(.in(layer_0[607]), .out(far_1_1229_0[1]));
    wire [1:0] far_1_1229_1;    relay_conn far_1_1229_1_a(.in(far_1_1229_0[0]), .out(far_1_1229_1[0]));    relay_conn far_1_1229_1_b(.in(far_1_1229_0[1]), .out(far_1_1229_1[1]));
    wire [1:0] far_1_1229_2;    relay_conn far_1_1229_2_a(.in(far_1_1229_1[0]), .out(far_1_1229_2[0]));    relay_conn far_1_1229_2_b(.in(far_1_1229_1[1]), .out(far_1_1229_2[1]));
    assign layer_1[209] = ~(far_1_1229_2[0] & far_1_1229_2[1]); 
    wire [1:0] far_1_1230_0;    relay_conn far_1_1230_0_a(.in(layer_0[902]), .out(far_1_1230_0[0]));    relay_conn far_1_1230_0_b(.in(layer_0[862]), .out(far_1_1230_0[1]));
    assign layer_1[210] = ~(far_1_1230_0[0] & far_1_1230_0[1]); 
    assign layer_1[211] = ~layer_0[1006]; 
    wire [1:0] far_1_1232_0;    relay_conn far_1_1232_0_a(.in(layer_0[444]), .out(far_1_1232_0[0]));    relay_conn far_1_1232_0_b(.in(layer_0[316]), .out(far_1_1232_0[1]));
    wire [1:0] far_1_1232_1;    relay_conn far_1_1232_1_a(.in(far_1_1232_0[0]), .out(far_1_1232_1[0]));    relay_conn far_1_1232_1_b(.in(far_1_1232_0[1]), .out(far_1_1232_1[1]));
    wire [1:0] far_1_1232_2;    relay_conn far_1_1232_2_a(.in(far_1_1232_1[0]), .out(far_1_1232_2[0]));    relay_conn far_1_1232_2_b(.in(far_1_1232_1[1]), .out(far_1_1232_2[1]));
    wire [1:0] far_1_1232_3;    relay_conn far_1_1232_3_a(.in(far_1_1232_2[0]), .out(far_1_1232_3[0]));    relay_conn far_1_1232_3_b(.in(far_1_1232_2[1]), .out(far_1_1232_3[1]));
    assign layer_1[212] = far_1_1232_3[0] & far_1_1232_3[1]; 
    wire [1:0] far_1_1233_0;    relay_conn far_1_1233_0_a(.in(layer_0[229]), .out(far_1_1233_0[0]));    relay_conn far_1_1233_0_b(.in(layer_0[321]), .out(far_1_1233_0[1]));
    wire [1:0] far_1_1233_1;    relay_conn far_1_1233_1_a(.in(far_1_1233_0[0]), .out(far_1_1233_1[0]));    relay_conn far_1_1233_1_b(.in(far_1_1233_0[1]), .out(far_1_1233_1[1]));
    assign layer_1[213] = far_1_1233_1[1] & ~far_1_1233_1[0]; 
    assign layer_1[214] = ~(layer_0[1010] ^ layer_0[1012]); 
    wire [1:0] far_1_1235_0;    relay_conn far_1_1235_0_a(.in(layer_0[573]), .out(far_1_1235_0[0]));    relay_conn far_1_1235_0_b(.in(layer_0[530]), .out(far_1_1235_0[1]));
    assign layer_1[215] = far_1_1235_0[1] & ~far_1_1235_0[0]; 
    wire [1:0] far_1_1236_0;    relay_conn far_1_1236_0_a(.in(layer_0[512]), .out(far_1_1236_0[0]));    relay_conn far_1_1236_0_b(.in(layer_0[419]), .out(far_1_1236_0[1]));
    wire [1:0] far_1_1236_1;    relay_conn far_1_1236_1_a(.in(far_1_1236_0[0]), .out(far_1_1236_1[0]));    relay_conn far_1_1236_1_b(.in(far_1_1236_0[1]), .out(far_1_1236_1[1]));
    assign layer_1[216] = ~(far_1_1236_1[0] & far_1_1236_1[1]); 
    wire [1:0] far_1_1237_0;    relay_conn far_1_1237_0_a(.in(layer_0[888]), .out(far_1_1237_0[0]));    relay_conn far_1_1237_0_b(.in(layer_0[952]), .out(far_1_1237_0[1]));
    wire [1:0] far_1_1237_1;    relay_conn far_1_1237_1_a(.in(far_1_1237_0[0]), .out(far_1_1237_1[0]));    relay_conn far_1_1237_1_b(.in(far_1_1237_0[1]), .out(far_1_1237_1[1]));
    assign layer_1[217] = ~(far_1_1237_1[0] & far_1_1237_1[1]); 
    wire [1:0] far_1_1238_0;    relay_conn far_1_1238_0_a(.in(layer_0[444]), .out(far_1_1238_0[0]));    relay_conn far_1_1238_0_b(.in(layer_0[338]), .out(far_1_1238_0[1]));
    wire [1:0] far_1_1238_1;    relay_conn far_1_1238_1_a(.in(far_1_1238_0[0]), .out(far_1_1238_1[0]));    relay_conn far_1_1238_1_b(.in(far_1_1238_0[1]), .out(far_1_1238_1[1]));
    wire [1:0] far_1_1238_2;    relay_conn far_1_1238_2_a(.in(far_1_1238_1[0]), .out(far_1_1238_2[0]));    relay_conn far_1_1238_2_b(.in(far_1_1238_1[1]), .out(far_1_1238_2[1]));
    assign layer_1[218] = ~far_1_1238_2[0] | (far_1_1238_2[0] & far_1_1238_2[1]); 
    wire [1:0] far_1_1239_0;    relay_conn far_1_1239_0_a(.in(layer_0[908]), .out(far_1_1239_0[0]));    relay_conn far_1_1239_0_b(.in(layer_0[967]), .out(far_1_1239_0[1]));
    assign layer_1[219] = far_1_1239_0[0]; 
    wire [1:0] far_1_1240_0;    relay_conn far_1_1240_0_a(.in(layer_0[942]), .out(far_1_1240_0[0]));    relay_conn far_1_1240_0_b(.in(layer_0[839]), .out(far_1_1240_0[1]));
    wire [1:0] far_1_1240_1;    relay_conn far_1_1240_1_a(.in(far_1_1240_0[0]), .out(far_1_1240_1[0]));    relay_conn far_1_1240_1_b(.in(far_1_1240_0[1]), .out(far_1_1240_1[1]));
    wire [1:0] far_1_1240_2;    relay_conn far_1_1240_2_a(.in(far_1_1240_1[0]), .out(far_1_1240_2[0]));    relay_conn far_1_1240_2_b(.in(far_1_1240_1[1]), .out(far_1_1240_2[1]));
    assign layer_1[220] = far_1_1240_2[0]; 
    wire [1:0] far_1_1241_0;    relay_conn far_1_1241_0_a(.in(layer_0[834]), .out(far_1_1241_0[0]));    relay_conn far_1_1241_0_b(.in(layer_0[954]), .out(far_1_1241_0[1]));
    wire [1:0] far_1_1241_1;    relay_conn far_1_1241_1_a(.in(far_1_1241_0[0]), .out(far_1_1241_1[0]));    relay_conn far_1_1241_1_b(.in(far_1_1241_0[1]), .out(far_1_1241_1[1]));
    wire [1:0] far_1_1241_2;    relay_conn far_1_1241_2_a(.in(far_1_1241_1[0]), .out(far_1_1241_2[0]));    relay_conn far_1_1241_2_b(.in(far_1_1241_1[1]), .out(far_1_1241_2[1]));
    assign layer_1[221] = ~far_1_1241_2[0] | (far_1_1241_2[0] & far_1_1241_2[1]); 
    wire [1:0] far_1_1242_0;    relay_conn far_1_1242_0_a(.in(layer_0[344]), .out(far_1_1242_0[0]));    relay_conn far_1_1242_0_b(.in(layer_0[395]), .out(far_1_1242_0[1]));
    assign layer_1[222] = ~far_1_1242_0[1]; 
    wire [1:0] far_1_1243_0;    relay_conn far_1_1243_0_a(.in(layer_0[477]), .out(far_1_1243_0[0]));    relay_conn far_1_1243_0_b(.in(layer_0[359]), .out(far_1_1243_0[1]));
    wire [1:0] far_1_1243_1;    relay_conn far_1_1243_1_a(.in(far_1_1243_0[0]), .out(far_1_1243_1[0]));    relay_conn far_1_1243_1_b(.in(far_1_1243_0[1]), .out(far_1_1243_1[1]));
    wire [1:0] far_1_1243_2;    relay_conn far_1_1243_2_a(.in(far_1_1243_1[0]), .out(far_1_1243_2[0]));    relay_conn far_1_1243_2_b(.in(far_1_1243_1[1]), .out(far_1_1243_2[1]));
    assign layer_1[223] = ~far_1_1243_2[1]; 
    wire [1:0] far_1_1244_0;    relay_conn far_1_1244_0_a(.in(layer_0[476]), .out(far_1_1244_0[0]));    relay_conn far_1_1244_0_b(.in(layer_0[438]), .out(far_1_1244_0[1]));
    assign layer_1[224] = far_1_1244_0[1]; 
    wire [1:0] far_1_1245_0;    relay_conn far_1_1245_0_a(.in(layer_0[289]), .out(far_1_1245_0[0]));    relay_conn far_1_1245_0_b(.in(layer_0[358]), .out(far_1_1245_0[1]));
    wire [1:0] far_1_1245_1;    relay_conn far_1_1245_1_a(.in(far_1_1245_0[0]), .out(far_1_1245_1[0]));    relay_conn far_1_1245_1_b(.in(far_1_1245_0[1]), .out(far_1_1245_1[1]));
    assign layer_1[225] = ~far_1_1245_1[1]; 
    assign layer_1[226] = layer_0[402]; 
    wire [1:0] far_1_1247_0;    relay_conn far_1_1247_0_a(.in(layer_0[241]), .out(far_1_1247_0[0]));    relay_conn far_1_1247_0_b(.in(layer_0[144]), .out(far_1_1247_0[1]));
    wire [1:0] far_1_1247_1;    relay_conn far_1_1247_1_a(.in(far_1_1247_0[0]), .out(far_1_1247_1[0]));    relay_conn far_1_1247_1_b(.in(far_1_1247_0[1]), .out(far_1_1247_1[1]));
    wire [1:0] far_1_1247_2;    relay_conn far_1_1247_2_a(.in(far_1_1247_1[0]), .out(far_1_1247_2[0]));    relay_conn far_1_1247_2_b(.in(far_1_1247_1[1]), .out(far_1_1247_2[1]));
    assign layer_1[227] = ~far_1_1247_2[1] | (far_1_1247_2[0] & far_1_1247_2[1]); 
    wire [1:0] far_1_1248_0;    relay_conn far_1_1248_0_a(.in(layer_0[455]), .out(far_1_1248_0[0]));    relay_conn far_1_1248_0_b(.in(layer_0[348]), .out(far_1_1248_0[1]));
    wire [1:0] far_1_1248_1;    relay_conn far_1_1248_1_a(.in(far_1_1248_0[0]), .out(far_1_1248_1[0]));    relay_conn far_1_1248_1_b(.in(far_1_1248_0[1]), .out(far_1_1248_1[1]));
    wire [1:0] far_1_1248_2;    relay_conn far_1_1248_2_a(.in(far_1_1248_1[0]), .out(far_1_1248_2[0]));    relay_conn far_1_1248_2_b(.in(far_1_1248_1[1]), .out(far_1_1248_2[1]));
    assign layer_1[228] = ~far_1_1248_2[1]; 
    wire [1:0] far_1_1249_0;    relay_conn far_1_1249_0_a(.in(layer_0[976]), .out(far_1_1249_0[0]));    relay_conn far_1_1249_0_b(.in(layer_0[861]), .out(far_1_1249_0[1]));
    wire [1:0] far_1_1249_1;    relay_conn far_1_1249_1_a(.in(far_1_1249_0[0]), .out(far_1_1249_1[0]));    relay_conn far_1_1249_1_b(.in(far_1_1249_0[1]), .out(far_1_1249_1[1]));
    wire [1:0] far_1_1249_2;    relay_conn far_1_1249_2_a(.in(far_1_1249_1[0]), .out(far_1_1249_2[0]));    relay_conn far_1_1249_2_b(.in(far_1_1249_1[1]), .out(far_1_1249_2[1]));
    assign layer_1[229] = far_1_1249_2[0] & ~far_1_1249_2[1]; 
    wire [1:0] far_1_1250_0;    relay_conn far_1_1250_0_a(.in(layer_0[246]), .out(far_1_1250_0[0]));    relay_conn far_1_1250_0_b(.in(layer_0[283]), .out(far_1_1250_0[1]));
    assign layer_1[230] = ~(far_1_1250_0[0] ^ far_1_1250_0[1]); 
    wire [1:0] far_1_1251_0;    relay_conn far_1_1251_0_a(.in(layer_0[35]), .out(far_1_1251_0[0]));    relay_conn far_1_1251_0_b(.in(layer_0[110]), .out(far_1_1251_0[1]));
    wire [1:0] far_1_1251_1;    relay_conn far_1_1251_1_a(.in(far_1_1251_0[0]), .out(far_1_1251_1[0]));    relay_conn far_1_1251_1_b(.in(far_1_1251_0[1]), .out(far_1_1251_1[1]));
    assign layer_1[231] = ~(far_1_1251_1[0] & far_1_1251_1[1]); 
    wire [1:0] far_1_1252_0;    relay_conn far_1_1252_0_a(.in(layer_0[417]), .out(far_1_1252_0[0]));    relay_conn far_1_1252_0_b(.in(layer_0[366]), .out(far_1_1252_0[1]));
    assign layer_1[232] = far_1_1252_0[0] & far_1_1252_0[1]; 
    wire [1:0] far_1_1253_0;    relay_conn far_1_1253_0_a(.in(layer_0[702]), .out(far_1_1253_0[0]));    relay_conn far_1_1253_0_b(.in(layer_0[766]), .out(far_1_1253_0[1]));
    wire [1:0] far_1_1253_1;    relay_conn far_1_1253_1_a(.in(far_1_1253_0[0]), .out(far_1_1253_1[0]));    relay_conn far_1_1253_1_b(.in(far_1_1253_0[1]), .out(far_1_1253_1[1]));
    assign layer_1[233] = ~far_1_1253_1[1] | (far_1_1253_1[0] & far_1_1253_1[1]); 
    wire [1:0] far_1_1254_0;    relay_conn far_1_1254_0_a(.in(layer_0[314]), .out(far_1_1254_0[0]));    relay_conn far_1_1254_0_b(.in(layer_0[257]), .out(far_1_1254_0[1]));
    assign layer_1[234] = far_1_1254_0[1]; 
    assign layer_1[235] = layer_0[561]; 
    assign layer_1[236] = layer_0[855]; 
    assign layer_1[237] = layer_0[490] & ~layer_0[480]; 
    wire [1:0] far_1_1258_0;    relay_conn far_1_1258_0_a(.in(layer_0[564]), .out(far_1_1258_0[0]));    relay_conn far_1_1258_0_b(.in(layer_0[607]), .out(far_1_1258_0[1]));
    assign layer_1[238] = ~(far_1_1258_0[0] | far_1_1258_0[1]); 
    wire [1:0] far_1_1259_0;    relay_conn far_1_1259_0_a(.in(layer_0[201]), .out(far_1_1259_0[0]));    relay_conn far_1_1259_0_b(.in(layer_0[263]), .out(far_1_1259_0[1]));
    assign layer_1[239] = far_1_1259_0[0] & far_1_1259_0[1]; 
    wire [1:0] far_1_1260_0;    relay_conn far_1_1260_0_a(.in(layer_0[282]), .out(far_1_1260_0[0]));    relay_conn far_1_1260_0_b(.in(layer_0[203]), .out(far_1_1260_0[1]));
    wire [1:0] far_1_1260_1;    relay_conn far_1_1260_1_a(.in(far_1_1260_0[0]), .out(far_1_1260_1[0]));    relay_conn far_1_1260_1_b(.in(far_1_1260_0[1]), .out(far_1_1260_1[1]));
    assign layer_1[240] = ~(far_1_1260_1[0] | far_1_1260_1[1]); 
    wire [1:0] far_1_1261_0;    relay_conn far_1_1261_0_a(.in(layer_0[117]), .out(far_1_1261_0[0]));    relay_conn far_1_1261_0_b(.in(layer_0[193]), .out(far_1_1261_0[1]));
    wire [1:0] far_1_1261_1;    relay_conn far_1_1261_1_a(.in(far_1_1261_0[0]), .out(far_1_1261_1[0]));    relay_conn far_1_1261_1_b(.in(far_1_1261_0[1]), .out(far_1_1261_1[1]));
    assign layer_1[241] = far_1_1261_1[0]; 
    wire [1:0] far_1_1262_0;    relay_conn far_1_1262_0_a(.in(layer_0[47]), .out(far_1_1262_0[0]));    relay_conn far_1_1262_0_b(.in(layer_0[108]), .out(far_1_1262_0[1]));
    assign layer_1[242] = ~(far_1_1262_0[0] & far_1_1262_0[1]); 
    wire [1:0] far_1_1263_0;    relay_conn far_1_1263_0_a(.in(layer_0[158]), .out(far_1_1263_0[0]));    relay_conn far_1_1263_0_b(.in(layer_0[205]), .out(far_1_1263_0[1]));
    assign layer_1[243] = ~far_1_1263_0[1]; 
    wire [1:0] far_1_1264_0;    relay_conn far_1_1264_0_a(.in(layer_0[273]), .out(far_1_1264_0[0]));    relay_conn far_1_1264_0_b(.in(layer_0[385]), .out(far_1_1264_0[1]));
    wire [1:0] far_1_1264_1;    relay_conn far_1_1264_1_a(.in(far_1_1264_0[0]), .out(far_1_1264_1[0]));    relay_conn far_1_1264_1_b(.in(far_1_1264_0[1]), .out(far_1_1264_1[1]));
    wire [1:0] far_1_1264_2;    relay_conn far_1_1264_2_a(.in(far_1_1264_1[0]), .out(far_1_1264_2[0]));    relay_conn far_1_1264_2_b(.in(far_1_1264_1[1]), .out(far_1_1264_2[1]));
    assign layer_1[244] = far_1_1264_2[1] & ~far_1_1264_2[0]; 
    wire [1:0] far_1_1265_0;    relay_conn far_1_1265_0_a(.in(layer_0[442]), .out(far_1_1265_0[0]));    relay_conn far_1_1265_0_b(.in(layer_0[474]), .out(far_1_1265_0[1]));
    assign layer_1[245] = ~(far_1_1265_0[0] & far_1_1265_0[1]); 
    assign layer_1[246] = layer_0[490] | layer_0[505]; 
    wire [1:0] far_1_1267_0;    relay_conn far_1_1267_0_a(.in(layer_0[434]), .out(far_1_1267_0[0]));    relay_conn far_1_1267_0_b(.in(layer_0[493]), .out(far_1_1267_0[1]));
    assign layer_1[247] = ~far_1_1267_0[1] | (far_1_1267_0[0] & far_1_1267_0[1]); 
    wire [1:0] far_1_1268_0;    relay_conn far_1_1268_0_a(.in(layer_0[220]), .out(far_1_1268_0[0]));    relay_conn far_1_1268_0_b(.in(layer_0[291]), .out(far_1_1268_0[1]));
    wire [1:0] far_1_1268_1;    relay_conn far_1_1268_1_a(.in(far_1_1268_0[0]), .out(far_1_1268_1[0]));    relay_conn far_1_1268_1_b(.in(far_1_1268_0[1]), .out(far_1_1268_1[1]));
    assign layer_1[248] = far_1_1268_1[0] & ~far_1_1268_1[1]; 
    assign layer_1[249] = layer_0[323]; 
    assign layer_1[250] = ~layer_0[193]; 
    wire [1:0] far_1_1271_0;    relay_conn far_1_1271_0_a(.in(layer_0[832]), .out(far_1_1271_0[0]));    relay_conn far_1_1271_0_b(.in(layer_0[946]), .out(far_1_1271_0[1]));
    wire [1:0] far_1_1271_1;    relay_conn far_1_1271_1_a(.in(far_1_1271_0[0]), .out(far_1_1271_1[0]));    relay_conn far_1_1271_1_b(.in(far_1_1271_0[1]), .out(far_1_1271_1[1]));
    wire [1:0] far_1_1271_2;    relay_conn far_1_1271_2_a(.in(far_1_1271_1[0]), .out(far_1_1271_2[0]));    relay_conn far_1_1271_2_b(.in(far_1_1271_1[1]), .out(far_1_1271_2[1]));
    assign layer_1[251] = ~(far_1_1271_2[0] | far_1_1271_2[1]); 
    wire [1:0] far_1_1272_0;    relay_conn far_1_1272_0_a(.in(layer_0[188]), .out(far_1_1272_0[0]));    relay_conn far_1_1272_0_b(.in(layer_0[292]), .out(far_1_1272_0[1]));
    wire [1:0] far_1_1272_1;    relay_conn far_1_1272_1_a(.in(far_1_1272_0[0]), .out(far_1_1272_1[0]));    relay_conn far_1_1272_1_b(.in(far_1_1272_0[1]), .out(far_1_1272_1[1]));
    wire [1:0] far_1_1272_2;    relay_conn far_1_1272_2_a(.in(far_1_1272_1[0]), .out(far_1_1272_2[0]));    relay_conn far_1_1272_2_b(.in(far_1_1272_1[1]), .out(far_1_1272_2[1]));
    assign layer_1[252] = ~(far_1_1272_2[0] & far_1_1272_2[1]); 
    assign layer_1[253] = ~layer_0[800] | (layer_0[773] & layer_0[800]); 
    wire [1:0] far_1_1274_0;    relay_conn far_1_1274_0_a(.in(layer_0[688]), .out(far_1_1274_0[0]));    relay_conn far_1_1274_0_b(.in(layer_0[816]), .out(far_1_1274_0[1]));
    wire [1:0] far_1_1274_1;    relay_conn far_1_1274_1_a(.in(far_1_1274_0[0]), .out(far_1_1274_1[0]));    relay_conn far_1_1274_1_b(.in(far_1_1274_0[1]), .out(far_1_1274_1[1]));
    wire [1:0] far_1_1274_2;    relay_conn far_1_1274_2_a(.in(far_1_1274_1[0]), .out(far_1_1274_2[0]));    relay_conn far_1_1274_2_b(.in(far_1_1274_1[1]), .out(far_1_1274_2[1]));
    wire [1:0] far_1_1274_3;    relay_conn far_1_1274_3_a(.in(far_1_1274_2[0]), .out(far_1_1274_3[0]));    relay_conn far_1_1274_3_b(.in(far_1_1274_2[1]), .out(far_1_1274_3[1]));
    assign layer_1[254] = far_1_1274_3[0] | far_1_1274_3[1]; 
    wire [1:0] far_1_1275_0;    relay_conn far_1_1275_0_a(.in(layer_0[683]), .out(far_1_1275_0[0]));    relay_conn far_1_1275_0_b(.in(layer_0[766]), .out(far_1_1275_0[1]));
    wire [1:0] far_1_1275_1;    relay_conn far_1_1275_1_a(.in(far_1_1275_0[0]), .out(far_1_1275_1[0]));    relay_conn far_1_1275_1_b(.in(far_1_1275_0[1]), .out(far_1_1275_1[1]));
    assign layer_1[255] = far_1_1275_1[0] & far_1_1275_1[1]; 
    assign layer_1[256] = ~layer_0[65]; 
    wire [1:0] far_1_1277_0;    relay_conn far_1_1277_0_a(.in(layer_0[539]), .out(far_1_1277_0[0]));    relay_conn far_1_1277_0_b(.in(layer_0[448]), .out(far_1_1277_0[1]));
    wire [1:0] far_1_1277_1;    relay_conn far_1_1277_1_a(.in(far_1_1277_0[0]), .out(far_1_1277_1[0]));    relay_conn far_1_1277_1_b(.in(far_1_1277_0[1]), .out(far_1_1277_1[1]));
    assign layer_1[257] = far_1_1277_1[0]; 
    assign layer_1[258] = layer_0[956]; 
    assign layer_1[259] = layer_0[293]; 
    wire [1:0] far_1_1280_0;    relay_conn far_1_1280_0_a(.in(layer_0[134]), .out(far_1_1280_0[0]));    relay_conn far_1_1280_0_b(.in(layer_0[255]), .out(far_1_1280_0[1]));
    wire [1:0] far_1_1280_1;    relay_conn far_1_1280_1_a(.in(far_1_1280_0[0]), .out(far_1_1280_1[0]));    relay_conn far_1_1280_1_b(.in(far_1_1280_0[1]), .out(far_1_1280_1[1]));
    wire [1:0] far_1_1280_2;    relay_conn far_1_1280_2_a(.in(far_1_1280_1[0]), .out(far_1_1280_2[0]));    relay_conn far_1_1280_2_b(.in(far_1_1280_1[1]), .out(far_1_1280_2[1]));
    assign layer_1[260] = far_1_1280_2[0] & far_1_1280_2[1]; 
    assign layer_1[261] = ~(layer_0[244] | layer_0[265]); 
    assign layer_1[262] = ~(layer_0[789] & layer_0[773]); 
    assign layer_1[263] = ~(layer_0[814] | layer_0[793]); 
    assign layer_1[264] = ~layer_0[116]; 
    wire [1:0] far_1_1285_0;    relay_conn far_1_1285_0_a(.in(layer_0[129]), .out(far_1_1285_0[0]));    relay_conn far_1_1285_0_b(.in(layer_0[221]), .out(far_1_1285_0[1]));
    wire [1:0] far_1_1285_1;    relay_conn far_1_1285_1_a(.in(far_1_1285_0[0]), .out(far_1_1285_1[0]));    relay_conn far_1_1285_1_b(.in(far_1_1285_0[1]), .out(far_1_1285_1[1]));
    assign layer_1[265] = ~far_1_1285_1[0]; 
    wire [1:0] far_1_1286_0;    relay_conn far_1_1286_0_a(.in(layer_0[485]), .out(far_1_1286_0[0]));    relay_conn far_1_1286_0_b(.in(layer_0[595]), .out(far_1_1286_0[1]));
    wire [1:0] far_1_1286_1;    relay_conn far_1_1286_1_a(.in(far_1_1286_0[0]), .out(far_1_1286_1[0]));    relay_conn far_1_1286_1_b(.in(far_1_1286_0[1]), .out(far_1_1286_1[1]));
    wire [1:0] far_1_1286_2;    relay_conn far_1_1286_2_a(.in(far_1_1286_1[0]), .out(far_1_1286_2[0]));    relay_conn far_1_1286_2_b(.in(far_1_1286_1[1]), .out(far_1_1286_2[1]));
    assign layer_1[266] = ~far_1_1286_2[0]; 
    assign layer_1[267] = layer_0[472] & layer_0[480]; 
    wire [1:0] far_1_1288_0;    relay_conn far_1_1288_0_a(.in(layer_0[378]), .out(far_1_1288_0[0]));    relay_conn far_1_1288_0_b(.in(layer_0[346]), .out(far_1_1288_0[1]));
    assign layer_1[268] = ~far_1_1288_0[0] | (far_1_1288_0[0] & far_1_1288_0[1]); 
    wire [1:0] far_1_1289_0;    relay_conn far_1_1289_0_a(.in(layer_0[1016]), .out(far_1_1289_0[0]));    relay_conn far_1_1289_0_b(.in(layer_0[889]), .out(far_1_1289_0[1]));
    wire [1:0] far_1_1289_1;    relay_conn far_1_1289_1_a(.in(far_1_1289_0[0]), .out(far_1_1289_1[0]));    relay_conn far_1_1289_1_b(.in(far_1_1289_0[1]), .out(far_1_1289_1[1]));
    wire [1:0] far_1_1289_2;    relay_conn far_1_1289_2_a(.in(far_1_1289_1[0]), .out(far_1_1289_2[0]));    relay_conn far_1_1289_2_b(.in(far_1_1289_1[1]), .out(far_1_1289_2[1]));
    assign layer_1[269] = ~far_1_1289_2[0]; 
    wire [1:0] far_1_1290_0;    relay_conn far_1_1290_0_a(.in(layer_0[489]), .out(far_1_1290_0[0]));    relay_conn far_1_1290_0_b(.in(layer_0[454]), .out(far_1_1290_0[1]));
    assign layer_1[270] = far_1_1290_0[1] & ~far_1_1290_0[0]; 
    wire [1:0] far_1_1291_0;    relay_conn far_1_1291_0_a(.in(layer_0[779]), .out(far_1_1291_0[0]));    relay_conn far_1_1291_0_b(.in(layer_0[696]), .out(far_1_1291_0[1]));
    wire [1:0] far_1_1291_1;    relay_conn far_1_1291_1_a(.in(far_1_1291_0[0]), .out(far_1_1291_1[0]));    relay_conn far_1_1291_1_b(.in(far_1_1291_0[1]), .out(far_1_1291_1[1]));
    assign layer_1[271] = far_1_1291_1[0] & ~far_1_1291_1[1]; 
    assign layer_1[272] = layer_0[699] & ~layer_0[698]; 
    wire [1:0] far_1_1293_0;    relay_conn far_1_1293_0_a(.in(layer_0[57]), .out(far_1_1293_0[0]));    relay_conn far_1_1293_0_b(.in(layer_0[11]), .out(far_1_1293_0[1]));
    assign layer_1[273] = far_1_1293_0[1]; 
    wire [1:0] far_1_1294_0;    relay_conn far_1_1294_0_a(.in(layer_0[20]), .out(far_1_1294_0[0]));    relay_conn far_1_1294_0_b(.in(layer_0[107]), .out(far_1_1294_0[1]));
    wire [1:0] far_1_1294_1;    relay_conn far_1_1294_1_a(.in(far_1_1294_0[0]), .out(far_1_1294_1[0]));    relay_conn far_1_1294_1_b(.in(far_1_1294_0[1]), .out(far_1_1294_1[1]));
    assign layer_1[274] = far_1_1294_1[0] & far_1_1294_1[1]; 
    wire [1:0] far_1_1295_0;    relay_conn far_1_1295_0_a(.in(layer_0[528]), .out(far_1_1295_0[0]));    relay_conn far_1_1295_0_b(.in(layer_0[481]), .out(far_1_1295_0[1]));
    assign layer_1[275] = far_1_1295_0[1]; 
    wire [1:0] far_1_1296_0;    relay_conn far_1_1296_0_a(.in(layer_0[852]), .out(far_1_1296_0[0]));    relay_conn far_1_1296_0_b(.in(layer_0[915]), .out(far_1_1296_0[1]));
    assign layer_1[276] = far_1_1296_0[0]; 
    wire [1:0] far_1_1297_0;    relay_conn far_1_1297_0_a(.in(layer_0[354]), .out(far_1_1297_0[0]));    relay_conn far_1_1297_0_b(.in(layer_0[475]), .out(far_1_1297_0[1]));
    wire [1:0] far_1_1297_1;    relay_conn far_1_1297_1_a(.in(far_1_1297_0[0]), .out(far_1_1297_1[0]));    relay_conn far_1_1297_1_b(.in(far_1_1297_0[1]), .out(far_1_1297_1[1]));
    wire [1:0] far_1_1297_2;    relay_conn far_1_1297_2_a(.in(far_1_1297_1[0]), .out(far_1_1297_2[0]));    relay_conn far_1_1297_2_b(.in(far_1_1297_1[1]), .out(far_1_1297_2[1]));
    assign layer_1[277] = ~far_1_1297_2[0]; 
    wire [1:0] far_1_1298_0;    relay_conn far_1_1298_0_a(.in(layer_0[395]), .out(far_1_1298_0[0]));    relay_conn far_1_1298_0_b(.in(layer_0[352]), .out(far_1_1298_0[1]));
    assign layer_1[278] = ~(far_1_1298_0[0] & far_1_1298_0[1]); 
    wire [1:0] far_1_1299_0;    relay_conn far_1_1299_0_a(.in(layer_0[702]), .out(far_1_1299_0[0]));    relay_conn far_1_1299_0_b(.in(layer_0[773]), .out(far_1_1299_0[1]));
    wire [1:0] far_1_1299_1;    relay_conn far_1_1299_1_a(.in(far_1_1299_0[0]), .out(far_1_1299_1[0]));    relay_conn far_1_1299_1_b(.in(far_1_1299_0[1]), .out(far_1_1299_1[1]));
    assign layer_1[279] = ~(far_1_1299_1[0] & far_1_1299_1[1]); 
    assign layer_1[280] = layer_0[236] ^ layer_0[223]; 
    assign layer_1[281] = layer_0[438]; 
    wire [1:0] far_1_1302_0;    relay_conn far_1_1302_0_a(.in(layer_0[49]), .out(far_1_1302_0[0]));    relay_conn far_1_1302_0_b(.in(layer_0[177]), .out(far_1_1302_0[1]));
    wire [1:0] far_1_1302_1;    relay_conn far_1_1302_1_a(.in(far_1_1302_0[0]), .out(far_1_1302_1[0]));    relay_conn far_1_1302_1_b(.in(far_1_1302_0[1]), .out(far_1_1302_1[1]));
    wire [1:0] far_1_1302_2;    relay_conn far_1_1302_2_a(.in(far_1_1302_1[0]), .out(far_1_1302_2[0]));    relay_conn far_1_1302_2_b(.in(far_1_1302_1[1]), .out(far_1_1302_2[1]));
    wire [1:0] far_1_1302_3;    relay_conn far_1_1302_3_a(.in(far_1_1302_2[0]), .out(far_1_1302_3[0]));    relay_conn far_1_1302_3_b(.in(far_1_1302_2[1]), .out(far_1_1302_3[1]));
    assign layer_1[282] = far_1_1302_3[0] | far_1_1302_3[1]; 
    assign layer_1[283] = layer_0[302] & ~layer_0[306]; 
    wire [1:0] far_1_1304_0;    relay_conn far_1_1304_0_a(.in(layer_0[506]), .out(far_1_1304_0[0]));    relay_conn far_1_1304_0_b(.in(layer_0[557]), .out(far_1_1304_0[1]));
    assign layer_1[284] = far_1_1304_0[0] & ~far_1_1304_0[1]; 
    assign layer_1[285] = layer_0[629] & layer_0[644]; 
    wire [1:0] far_1_1306_0;    relay_conn far_1_1306_0_a(.in(layer_0[413]), .out(far_1_1306_0[0]));    relay_conn far_1_1306_0_b(.in(layer_0[347]), .out(far_1_1306_0[1]));
    wire [1:0] far_1_1306_1;    relay_conn far_1_1306_1_a(.in(far_1_1306_0[0]), .out(far_1_1306_1[0]));    relay_conn far_1_1306_1_b(.in(far_1_1306_0[1]), .out(far_1_1306_1[1]));
    assign layer_1[286] = far_1_1306_1[0]; 
    assign layer_1[287] = layer_0[261]; 
    wire [1:0] far_1_1308_0;    relay_conn far_1_1308_0_a(.in(layer_0[432]), .out(far_1_1308_0[0]));    relay_conn far_1_1308_0_b(.in(layer_0[395]), .out(far_1_1308_0[1]));
    assign layer_1[288] = far_1_1308_0[0]; 
    wire [1:0] far_1_1309_0;    relay_conn far_1_1309_0_a(.in(layer_0[497]), .out(far_1_1309_0[0]));    relay_conn far_1_1309_0_b(.in(layer_0[544]), .out(far_1_1309_0[1]));
    assign layer_1[289] = ~far_1_1309_0[0]; 
    wire [1:0] far_1_1310_0;    relay_conn far_1_1310_0_a(.in(layer_0[628]), .out(far_1_1310_0[0]));    relay_conn far_1_1310_0_b(.in(layer_0[551]), .out(far_1_1310_0[1]));
    wire [1:0] far_1_1310_1;    relay_conn far_1_1310_1_a(.in(far_1_1310_0[0]), .out(far_1_1310_1[0]));    relay_conn far_1_1310_1_b(.in(far_1_1310_0[1]), .out(far_1_1310_1[1]));
    assign layer_1[290] = ~far_1_1310_1[0] | (far_1_1310_1[0] & far_1_1310_1[1]); 
    assign layer_1[291] = ~layer_0[705]; 
    wire [1:0] far_1_1312_0;    relay_conn far_1_1312_0_a(.in(layer_0[886]), .out(far_1_1312_0[0]));    relay_conn far_1_1312_0_b(.in(layer_0[942]), .out(far_1_1312_0[1]));
    assign layer_1[292] = far_1_1312_0[0] & ~far_1_1312_0[1]; 
    wire [1:0] far_1_1313_0;    relay_conn far_1_1313_0_a(.in(layer_0[816]), .out(far_1_1313_0[0]));    relay_conn far_1_1313_0_b(.in(layer_0[705]), .out(far_1_1313_0[1]));
    wire [1:0] far_1_1313_1;    relay_conn far_1_1313_1_a(.in(far_1_1313_0[0]), .out(far_1_1313_1[0]));    relay_conn far_1_1313_1_b(.in(far_1_1313_0[1]), .out(far_1_1313_1[1]));
    wire [1:0] far_1_1313_2;    relay_conn far_1_1313_2_a(.in(far_1_1313_1[0]), .out(far_1_1313_2[0]));    relay_conn far_1_1313_2_b(.in(far_1_1313_1[1]), .out(far_1_1313_2[1]));
    assign layer_1[293] = ~far_1_1313_2[0]; 
    assign layer_1[294] = layer_0[301] & ~layer_0[326]; 
    wire [1:0] far_1_1315_0;    relay_conn far_1_1315_0_a(.in(layer_0[577]), .out(far_1_1315_0[0]));    relay_conn far_1_1315_0_b(.in(layer_0[701]), .out(far_1_1315_0[1]));
    wire [1:0] far_1_1315_1;    relay_conn far_1_1315_1_a(.in(far_1_1315_0[0]), .out(far_1_1315_1[0]));    relay_conn far_1_1315_1_b(.in(far_1_1315_0[1]), .out(far_1_1315_1[1]));
    wire [1:0] far_1_1315_2;    relay_conn far_1_1315_2_a(.in(far_1_1315_1[0]), .out(far_1_1315_2[0]));    relay_conn far_1_1315_2_b(.in(far_1_1315_1[1]), .out(far_1_1315_2[1]));
    assign layer_1[295] = ~far_1_1315_2[1] | (far_1_1315_2[0] & far_1_1315_2[1]); 
    wire [1:0] far_1_1316_0;    relay_conn far_1_1316_0_a(.in(layer_0[597]), .out(far_1_1316_0[0]));    relay_conn far_1_1316_0_b(.in(layer_0[684]), .out(far_1_1316_0[1]));
    wire [1:0] far_1_1316_1;    relay_conn far_1_1316_1_a(.in(far_1_1316_0[0]), .out(far_1_1316_1[0]));    relay_conn far_1_1316_1_b(.in(far_1_1316_0[1]), .out(far_1_1316_1[1]));
    assign layer_1[296] = far_1_1316_1[1] & ~far_1_1316_1[0]; 
    wire [1:0] far_1_1317_0;    relay_conn far_1_1317_0_a(.in(layer_0[663]), .out(far_1_1317_0[0]));    relay_conn far_1_1317_0_b(.in(layer_0[715]), .out(far_1_1317_0[1]));
    assign layer_1[297] = far_1_1317_0[0] ^ far_1_1317_0[1]; 
    assign layer_1[298] = ~(layer_0[372] & layer_0[364]); 
    wire [1:0] far_1_1319_0;    relay_conn far_1_1319_0_a(.in(layer_0[844]), .out(far_1_1319_0[0]));    relay_conn far_1_1319_0_b(.in(layer_0[964]), .out(far_1_1319_0[1]));
    wire [1:0] far_1_1319_1;    relay_conn far_1_1319_1_a(.in(far_1_1319_0[0]), .out(far_1_1319_1[0]));    relay_conn far_1_1319_1_b(.in(far_1_1319_0[1]), .out(far_1_1319_1[1]));
    wire [1:0] far_1_1319_2;    relay_conn far_1_1319_2_a(.in(far_1_1319_1[0]), .out(far_1_1319_2[0]));    relay_conn far_1_1319_2_b(.in(far_1_1319_1[1]), .out(far_1_1319_2[1]));
    assign layer_1[299] = ~(far_1_1319_2[0] ^ far_1_1319_2[1]); 
    wire [1:0] far_1_1320_0;    relay_conn far_1_1320_0_a(.in(layer_0[429]), .out(far_1_1320_0[0]));    relay_conn far_1_1320_0_b(.in(layer_0[468]), .out(far_1_1320_0[1]));
    assign layer_1[300] = ~far_1_1320_0[1] | (far_1_1320_0[0] & far_1_1320_0[1]); 
    assign layer_1[301] = ~layer_0[501]; 
    wire [1:0] far_1_1322_0;    relay_conn far_1_1322_0_a(.in(layer_0[967]), .out(far_1_1322_0[0]));    relay_conn far_1_1322_0_b(.in(layer_0[1019]), .out(far_1_1322_0[1]));
    assign layer_1[302] = far_1_1322_0[0] | far_1_1322_0[1]; 
    assign layer_1[303] = layer_0[65] ^ layer_0[62]; 
    wire [1:0] far_1_1324_0;    relay_conn far_1_1324_0_a(.in(layer_0[38]), .out(far_1_1324_0[0]));    relay_conn far_1_1324_0_b(.in(layer_0[93]), .out(far_1_1324_0[1]));
    assign layer_1[304] = ~far_1_1324_0[1]; 
    wire [1:0] far_1_1325_0;    relay_conn far_1_1325_0_a(.in(layer_0[429]), .out(far_1_1325_0[0]));    relay_conn far_1_1325_0_b(.in(layer_0[531]), .out(far_1_1325_0[1]));
    wire [1:0] far_1_1325_1;    relay_conn far_1_1325_1_a(.in(far_1_1325_0[0]), .out(far_1_1325_1[0]));    relay_conn far_1_1325_1_b(.in(far_1_1325_0[1]), .out(far_1_1325_1[1]));
    wire [1:0] far_1_1325_2;    relay_conn far_1_1325_2_a(.in(far_1_1325_1[0]), .out(far_1_1325_2[0]));    relay_conn far_1_1325_2_b(.in(far_1_1325_1[1]), .out(far_1_1325_2[1]));
    assign layer_1[305] = far_1_1325_2[1] & ~far_1_1325_2[0]; 
    wire [1:0] far_1_1326_0;    relay_conn far_1_1326_0_a(.in(layer_0[527]), .out(far_1_1326_0[0]));    relay_conn far_1_1326_0_b(.in(layer_0[429]), .out(far_1_1326_0[1]));
    wire [1:0] far_1_1326_1;    relay_conn far_1_1326_1_a(.in(far_1_1326_0[0]), .out(far_1_1326_1[0]));    relay_conn far_1_1326_1_b(.in(far_1_1326_0[1]), .out(far_1_1326_1[1]));
    wire [1:0] far_1_1326_2;    relay_conn far_1_1326_2_a(.in(far_1_1326_1[0]), .out(far_1_1326_2[0]));    relay_conn far_1_1326_2_b(.in(far_1_1326_1[1]), .out(far_1_1326_2[1]));
    assign layer_1[306] = far_1_1326_2[1]; 
    wire [1:0] far_1_1327_0;    relay_conn far_1_1327_0_a(.in(layer_0[65]), .out(far_1_1327_0[0]));    relay_conn far_1_1327_0_b(.in(layer_0[156]), .out(far_1_1327_0[1]));
    wire [1:0] far_1_1327_1;    relay_conn far_1_1327_1_a(.in(far_1_1327_0[0]), .out(far_1_1327_1[0]));    relay_conn far_1_1327_1_b(.in(far_1_1327_0[1]), .out(far_1_1327_1[1]));
    assign layer_1[307] = far_1_1327_1[0] & far_1_1327_1[1]; 
    wire [1:0] far_1_1328_0;    relay_conn far_1_1328_0_a(.in(layer_0[697]), .out(far_1_1328_0[0]));    relay_conn far_1_1328_0_b(.in(layer_0[799]), .out(far_1_1328_0[1]));
    wire [1:0] far_1_1328_1;    relay_conn far_1_1328_1_a(.in(far_1_1328_0[0]), .out(far_1_1328_1[0]));    relay_conn far_1_1328_1_b(.in(far_1_1328_0[1]), .out(far_1_1328_1[1]));
    wire [1:0] far_1_1328_2;    relay_conn far_1_1328_2_a(.in(far_1_1328_1[0]), .out(far_1_1328_2[0]));    relay_conn far_1_1328_2_b(.in(far_1_1328_1[1]), .out(far_1_1328_2[1]));
    assign layer_1[308] = ~far_1_1328_2[1]; 
    wire [1:0] far_1_1329_0;    relay_conn far_1_1329_0_a(.in(layer_0[253]), .out(far_1_1329_0[0]));    relay_conn far_1_1329_0_b(.in(layer_0[289]), .out(far_1_1329_0[1]));
    assign layer_1[309] = ~far_1_1329_0[0]; 
    assign layer_1[310] = ~(layer_0[365] & layer_0[374]); 
    wire [1:0] far_1_1331_0;    relay_conn far_1_1331_0_a(.in(layer_0[909]), .out(far_1_1331_0[0]));    relay_conn far_1_1331_0_b(.in(layer_0[833]), .out(far_1_1331_0[1]));
    wire [1:0] far_1_1331_1;    relay_conn far_1_1331_1_a(.in(far_1_1331_0[0]), .out(far_1_1331_1[0]));    relay_conn far_1_1331_1_b(.in(far_1_1331_0[1]), .out(far_1_1331_1[1]));
    assign layer_1[311] = ~far_1_1331_1[0]; 
    wire [1:0] far_1_1332_0;    relay_conn far_1_1332_0_a(.in(layer_0[810]), .out(far_1_1332_0[0]));    relay_conn far_1_1332_0_b(.in(layer_0[909]), .out(far_1_1332_0[1]));
    wire [1:0] far_1_1332_1;    relay_conn far_1_1332_1_a(.in(far_1_1332_0[0]), .out(far_1_1332_1[0]));    relay_conn far_1_1332_1_b(.in(far_1_1332_0[1]), .out(far_1_1332_1[1]));
    wire [1:0] far_1_1332_2;    relay_conn far_1_1332_2_a(.in(far_1_1332_1[0]), .out(far_1_1332_2[0]));    relay_conn far_1_1332_2_b(.in(far_1_1332_1[1]), .out(far_1_1332_2[1]));
    assign layer_1[312] = far_1_1332_2[0] & ~far_1_1332_2[1]; 
    assign layer_1[313] = ~layer_0[957]; 
    wire [1:0] far_1_1334_0;    relay_conn far_1_1334_0_a(.in(layer_0[43]), .out(far_1_1334_0[0]));    relay_conn far_1_1334_0_b(.in(layer_0[94]), .out(far_1_1334_0[1]));
    assign layer_1[314] = far_1_1334_0[0] | far_1_1334_0[1]; 
    wire [1:0] far_1_1335_0;    relay_conn far_1_1335_0_a(.in(layer_0[849]), .out(far_1_1335_0[0]));    relay_conn far_1_1335_0_b(.in(layer_0[773]), .out(far_1_1335_0[1]));
    wire [1:0] far_1_1335_1;    relay_conn far_1_1335_1_a(.in(far_1_1335_0[0]), .out(far_1_1335_1[0]));    relay_conn far_1_1335_1_b(.in(far_1_1335_0[1]), .out(far_1_1335_1[1]));
    assign layer_1[315] = far_1_1335_1[0] & far_1_1335_1[1]; 
    wire [1:0] far_1_1336_0;    relay_conn far_1_1336_0_a(.in(layer_0[2]), .out(far_1_1336_0[0]));    relay_conn far_1_1336_0_b(.in(layer_0[71]), .out(far_1_1336_0[1]));
    wire [1:0] far_1_1336_1;    relay_conn far_1_1336_1_a(.in(far_1_1336_0[0]), .out(far_1_1336_1[0]));    relay_conn far_1_1336_1_b(.in(far_1_1336_0[1]), .out(far_1_1336_1[1]));
    assign layer_1[316] = ~(far_1_1336_1[0] | far_1_1336_1[1]); 
    assign layer_1[317] = layer_0[1019] ^ layer_0[996]; 
    wire [1:0] far_1_1338_0;    relay_conn far_1_1338_0_a(.in(layer_0[441]), .out(far_1_1338_0[0]));    relay_conn far_1_1338_0_b(.in(layer_0[512]), .out(far_1_1338_0[1]));
    wire [1:0] far_1_1338_1;    relay_conn far_1_1338_1_a(.in(far_1_1338_0[0]), .out(far_1_1338_1[0]));    relay_conn far_1_1338_1_b(.in(far_1_1338_0[1]), .out(far_1_1338_1[1]));
    assign layer_1[318] = far_1_1338_1[1] & ~far_1_1338_1[0]; 
    wire [1:0] far_1_1339_0;    relay_conn far_1_1339_0_a(.in(layer_0[909]), .out(far_1_1339_0[0]));    relay_conn far_1_1339_0_b(.in(layer_0[789]), .out(far_1_1339_0[1]));
    wire [1:0] far_1_1339_1;    relay_conn far_1_1339_1_a(.in(far_1_1339_0[0]), .out(far_1_1339_1[0]));    relay_conn far_1_1339_1_b(.in(far_1_1339_0[1]), .out(far_1_1339_1[1]));
    wire [1:0] far_1_1339_2;    relay_conn far_1_1339_2_a(.in(far_1_1339_1[0]), .out(far_1_1339_2[0]));    relay_conn far_1_1339_2_b(.in(far_1_1339_1[1]), .out(far_1_1339_2[1]));
    assign layer_1[319] = ~far_1_1339_2[0]; 
    assign layer_1[320] = layer_0[686]; 
    wire [1:0] far_1_1341_0;    relay_conn far_1_1341_0_a(.in(layer_0[556]), .out(far_1_1341_0[0]));    relay_conn far_1_1341_0_b(.in(layer_0[480]), .out(far_1_1341_0[1]));
    wire [1:0] far_1_1341_1;    relay_conn far_1_1341_1_a(.in(far_1_1341_0[0]), .out(far_1_1341_1[0]));    relay_conn far_1_1341_1_b(.in(far_1_1341_0[1]), .out(far_1_1341_1[1]));
    assign layer_1[321] = ~far_1_1341_1[1] | (far_1_1341_1[0] & far_1_1341_1[1]); 
    wire [1:0] far_1_1342_0;    relay_conn far_1_1342_0_a(.in(layer_0[997]), .out(far_1_1342_0[0]));    relay_conn far_1_1342_0_b(.in(layer_0[888]), .out(far_1_1342_0[1]));
    wire [1:0] far_1_1342_1;    relay_conn far_1_1342_1_a(.in(far_1_1342_0[0]), .out(far_1_1342_1[0]));    relay_conn far_1_1342_1_b(.in(far_1_1342_0[1]), .out(far_1_1342_1[1]));
    wire [1:0] far_1_1342_2;    relay_conn far_1_1342_2_a(.in(far_1_1342_1[0]), .out(far_1_1342_2[0]));    relay_conn far_1_1342_2_b(.in(far_1_1342_1[1]), .out(far_1_1342_2[1]));
    assign layer_1[322] = far_1_1342_2[0] ^ far_1_1342_2[1]; 
    assign layer_1[323] = ~(layer_0[305] ^ layer_0[331]); 
    wire [1:0] far_1_1344_0;    relay_conn far_1_1344_0_a(.in(layer_0[21]), .out(far_1_1344_0[0]));    relay_conn far_1_1344_0_b(.in(layer_0[91]), .out(far_1_1344_0[1]));
    wire [1:0] far_1_1344_1;    relay_conn far_1_1344_1_a(.in(far_1_1344_0[0]), .out(far_1_1344_1[0]));    relay_conn far_1_1344_1_b(.in(far_1_1344_0[1]), .out(far_1_1344_1[1]));
    assign layer_1[324] = ~far_1_1344_1[0]; 
    assign layer_1[325] = ~(layer_0[93] & layer_0[73]); 
    wire [1:0] far_1_1346_0;    relay_conn far_1_1346_0_a(.in(layer_0[490]), .out(far_1_1346_0[0]));    relay_conn far_1_1346_0_b(.in(layer_0[375]), .out(far_1_1346_0[1]));
    wire [1:0] far_1_1346_1;    relay_conn far_1_1346_1_a(.in(far_1_1346_0[0]), .out(far_1_1346_1[0]));    relay_conn far_1_1346_1_b(.in(far_1_1346_0[1]), .out(far_1_1346_1[1]));
    wire [1:0] far_1_1346_2;    relay_conn far_1_1346_2_a(.in(far_1_1346_1[0]), .out(far_1_1346_2[0]));    relay_conn far_1_1346_2_b(.in(far_1_1346_1[1]), .out(far_1_1346_2[1]));
    assign layer_1[326] = far_1_1346_2[1]; 
    wire [1:0] far_1_1347_0;    relay_conn far_1_1347_0_a(.in(layer_0[484]), .out(far_1_1347_0[0]));    relay_conn far_1_1347_0_b(.in(layer_0[610]), .out(far_1_1347_0[1]));
    wire [1:0] far_1_1347_1;    relay_conn far_1_1347_1_a(.in(far_1_1347_0[0]), .out(far_1_1347_1[0]));    relay_conn far_1_1347_1_b(.in(far_1_1347_0[1]), .out(far_1_1347_1[1]));
    wire [1:0] far_1_1347_2;    relay_conn far_1_1347_2_a(.in(far_1_1347_1[0]), .out(far_1_1347_2[0]));    relay_conn far_1_1347_2_b(.in(far_1_1347_1[1]), .out(far_1_1347_2[1]));
    assign layer_1[327] = ~(far_1_1347_2[0] ^ far_1_1347_2[1]); 
    assign layer_1[328] = layer_0[487] & ~layer_0[509]; 
    wire [1:0] far_1_1349_0;    relay_conn far_1_1349_0_a(.in(layer_0[748]), .out(far_1_1349_0[0]));    relay_conn far_1_1349_0_b(.in(layer_0[696]), .out(far_1_1349_0[1]));
    assign layer_1[329] = ~(far_1_1349_0[0] | far_1_1349_0[1]); 
    wire [1:0] far_1_1350_0;    relay_conn far_1_1350_0_a(.in(layer_0[330]), .out(far_1_1350_0[0]));    relay_conn far_1_1350_0_b(.in(layer_0[204]), .out(far_1_1350_0[1]));
    wire [1:0] far_1_1350_1;    relay_conn far_1_1350_1_a(.in(far_1_1350_0[0]), .out(far_1_1350_1[0]));    relay_conn far_1_1350_1_b(.in(far_1_1350_0[1]), .out(far_1_1350_1[1]));
    wire [1:0] far_1_1350_2;    relay_conn far_1_1350_2_a(.in(far_1_1350_1[0]), .out(far_1_1350_2[0]));    relay_conn far_1_1350_2_b(.in(far_1_1350_1[1]), .out(far_1_1350_2[1]));
    assign layer_1[330] = ~(far_1_1350_2[0] & far_1_1350_2[1]); 
    wire [1:0] far_1_1351_0;    relay_conn far_1_1351_0_a(.in(layer_0[356]), .out(far_1_1351_0[0]));    relay_conn far_1_1351_0_b(.in(layer_0[263]), .out(far_1_1351_0[1]));
    wire [1:0] far_1_1351_1;    relay_conn far_1_1351_1_a(.in(far_1_1351_0[0]), .out(far_1_1351_1[0]));    relay_conn far_1_1351_1_b(.in(far_1_1351_0[1]), .out(far_1_1351_1[1]));
    assign layer_1[331] = far_1_1351_1[1] & ~far_1_1351_1[0]; 
    wire [1:0] far_1_1352_0;    relay_conn far_1_1352_0_a(.in(layer_0[394]), .out(far_1_1352_0[0]));    relay_conn far_1_1352_0_b(.in(layer_0[329]), .out(far_1_1352_0[1]));
    wire [1:0] far_1_1352_1;    relay_conn far_1_1352_1_a(.in(far_1_1352_0[0]), .out(far_1_1352_1[0]));    relay_conn far_1_1352_1_b(.in(far_1_1352_0[1]), .out(far_1_1352_1[1]));
    assign layer_1[332] = ~far_1_1352_1[1] | (far_1_1352_1[0] & far_1_1352_1[1]); 
    wire [1:0] far_1_1353_0;    relay_conn far_1_1353_0_a(.in(layer_0[706]), .out(far_1_1353_0[0]));    relay_conn far_1_1353_0_b(.in(layer_0[748]), .out(far_1_1353_0[1]));
    assign layer_1[333] = ~far_1_1353_0[1]; 
    wire [1:0] far_1_1354_0;    relay_conn far_1_1354_0_a(.in(layer_0[231]), .out(far_1_1354_0[0]));    relay_conn far_1_1354_0_b(.in(layer_0[336]), .out(far_1_1354_0[1]));
    wire [1:0] far_1_1354_1;    relay_conn far_1_1354_1_a(.in(far_1_1354_0[0]), .out(far_1_1354_1[0]));    relay_conn far_1_1354_1_b(.in(far_1_1354_0[1]), .out(far_1_1354_1[1]));
    wire [1:0] far_1_1354_2;    relay_conn far_1_1354_2_a(.in(far_1_1354_1[0]), .out(far_1_1354_2[0]));    relay_conn far_1_1354_2_b(.in(far_1_1354_1[1]), .out(far_1_1354_2[1]));
    assign layer_1[334] = ~far_1_1354_2[0]; 
    wire [1:0] far_1_1355_0;    relay_conn far_1_1355_0_a(.in(layer_0[1018]), .out(far_1_1355_0[0]));    relay_conn far_1_1355_0_b(.in(layer_0[927]), .out(far_1_1355_0[1]));
    wire [1:0] far_1_1355_1;    relay_conn far_1_1355_1_a(.in(far_1_1355_0[0]), .out(far_1_1355_1[0]));    relay_conn far_1_1355_1_b(.in(far_1_1355_0[1]), .out(far_1_1355_1[1]));
    assign layer_1[335] = far_1_1355_1[1] & ~far_1_1355_1[0]; 
    wire [1:0] far_1_1356_0;    relay_conn far_1_1356_0_a(.in(layer_0[171]), .out(far_1_1356_0[0]));    relay_conn far_1_1356_0_b(.in(layer_0[263]), .out(far_1_1356_0[1]));
    wire [1:0] far_1_1356_1;    relay_conn far_1_1356_1_a(.in(far_1_1356_0[0]), .out(far_1_1356_1[0]));    relay_conn far_1_1356_1_b(.in(far_1_1356_0[1]), .out(far_1_1356_1[1]));
    assign layer_1[336] = ~(far_1_1356_1[0] & far_1_1356_1[1]); 
    wire [1:0] far_1_1357_0;    relay_conn far_1_1357_0_a(.in(layer_0[253]), .out(far_1_1357_0[0]));    relay_conn far_1_1357_0_b(.in(layer_0[381]), .out(far_1_1357_0[1]));
    wire [1:0] far_1_1357_1;    relay_conn far_1_1357_1_a(.in(far_1_1357_0[0]), .out(far_1_1357_1[0]));    relay_conn far_1_1357_1_b(.in(far_1_1357_0[1]), .out(far_1_1357_1[1]));
    wire [1:0] far_1_1357_2;    relay_conn far_1_1357_2_a(.in(far_1_1357_1[0]), .out(far_1_1357_2[0]));    relay_conn far_1_1357_2_b(.in(far_1_1357_1[1]), .out(far_1_1357_2[1]));
    wire [1:0] far_1_1357_3;    relay_conn far_1_1357_3_a(.in(far_1_1357_2[0]), .out(far_1_1357_3[0]));    relay_conn far_1_1357_3_b(.in(far_1_1357_2[1]), .out(far_1_1357_3[1]));
    assign layer_1[337] = ~(far_1_1357_3[0] | far_1_1357_3[1]); 
    wire [1:0] far_1_1358_0;    relay_conn far_1_1358_0_a(.in(layer_0[734]), .out(far_1_1358_0[0]));    relay_conn far_1_1358_0_b(.in(layer_0[619]), .out(far_1_1358_0[1]));
    wire [1:0] far_1_1358_1;    relay_conn far_1_1358_1_a(.in(far_1_1358_0[0]), .out(far_1_1358_1[0]));    relay_conn far_1_1358_1_b(.in(far_1_1358_0[1]), .out(far_1_1358_1[1]));
    wire [1:0] far_1_1358_2;    relay_conn far_1_1358_2_a(.in(far_1_1358_1[0]), .out(far_1_1358_2[0]));    relay_conn far_1_1358_2_b(.in(far_1_1358_1[1]), .out(far_1_1358_2[1]));
    assign layer_1[338] = far_1_1358_2[1] & ~far_1_1358_2[0]; 
    wire [1:0] far_1_1359_0;    relay_conn far_1_1359_0_a(.in(layer_0[562]), .out(far_1_1359_0[0]));    relay_conn far_1_1359_0_b(.in(layer_0[512]), .out(far_1_1359_0[1]));
    assign layer_1[339] = far_1_1359_0[1] & ~far_1_1359_0[0]; 
    assign layer_1[340] = ~layer_0[914]; 
    wire [1:0] far_1_1361_0;    relay_conn far_1_1361_0_a(.in(layer_0[737]), .out(far_1_1361_0[0]));    relay_conn far_1_1361_0_b(.in(layer_0[638]), .out(far_1_1361_0[1]));
    wire [1:0] far_1_1361_1;    relay_conn far_1_1361_1_a(.in(far_1_1361_0[0]), .out(far_1_1361_1[0]));    relay_conn far_1_1361_1_b(.in(far_1_1361_0[1]), .out(far_1_1361_1[1]));
    wire [1:0] far_1_1361_2;    relay_conn far_1_1361_2_a(.in(far_1_1361_1[0]), .out(far_1_1361_2[0]));    relay_conn far_1_1361_2_b(.in(far_1_1361_1[1]), .out(far_1_1361_2[1]));
    assign layer_1[341] = ~(far_1_1361_2[0] & far_1_1361_2[1]); 
    assign layer_1[342] = layer_0[367] & ~layer_0[397]; 
    wire [1:0] far_1_1363_0;    relay_conn far_1_1363_0_a(.in(layer_0[49]), .out(far_1_1363_0[0]));    relay_conn far_1_1363_0_b(.in(layer_0[81]), .out(far_1_1363_0[1]));
    assign layer_1[343] = ~far_1_1363_0[0] | (far_1_1363_0[0] & far_1_1363_0[1]); 
    wire [1:0] far_1_1364_0;    relay_conn far_1_1364_0_a(.in(layer_0[387]), .out(far_1_1364_0[0]));    relay_conn far_1_1364_0_b(.in(layer_0[265]), .out(far_1_1364_0[1]));
    wire [1:0] far_1_1364_1;    relay_conn far_1_1364_1_a(.in(far_1_1364_0[0]), .out(far_1_1364_1[0]));    relay_conn far_1_1364_1_b(.in(far_1_1364_0[1]), .out(far_1_1364_1[1]));
    wire [1:0] far_1_1364_2;    relay_conn far_1_1364_2_a(.in(far_1_1364_1[0]), .out(far_1_1364_2[0]));    relay_conn far_1_1364_2_b(.in(far_1_1364_1[1]), .out(far_1_1364_2[1]));
    assign layer_1[344] = ~(far_1_1364_2[0] | far_1_1364_2[1]); 
    wire [1:0] far_1_1365_0;    relay_conn far_1_1365_0_a(.in(layer_0[418]), .out(far_1_1365_0[0]));    relay_conn far_1_1365_0_b(.in(layer_0[543]), .out(far_1_1365_0[1]));
    wire [1:0] far_1_1365_1;    relay_conn far_1_1365_1_a(.in(far_1_1365_0[0]), .out(far_1_1365_1[0]));    relay_conn far_1_1365_1_b(.in(far_1_1365_0[1]), .out(far_1_1365_1[1]));
    wire [1:0] far_1_1365_2;    relay_conn far_1_1365_2_a(.in(far_1_1365_1[0]), .out(far_1_1365_2[0]));    relay_conn far_1_1365_2_b(.in(far_1_1365_1[1]), .out(far_1_1365_2[1]));
    assign layer_1[345] = ~far_1_1365_2[1]; 
    wire [1:0] far_1_1366_0;    relay_conn far_1_1366_0_a(.in(layer_0[867]), .out(far_1_1366_0[0]));    relay_conn far_1_1366_0_b(.in(layer_0[909]), .out(far_1_1366_0[1]));
    assign layer_1[346] = ~far_1_1366_0[0] | (far_1_1366_0[0] & far_1_1366_0[1]); 
    wire [1:0] far_1_1367_0;    relay_conn far_1_1367_0_a(.in(layer_0[656]), .out(far_1_1367_0[0]));    relay_conn far_1_1367_0_b(.in(layer_0[543]), .out(far_1_1367_0[1]));
    wire [1:0] far_1_1367_1;    relay_conn far_1_1367_1_a(.in(far_1_1367_0[0]), .out(far_1_1367_1[0]));    relay_conn far_1_1367_1_b(.in(far_1_1367_0[1]), .out(far_1_1367_1[1]));
    wire [1:0] far_1_1367_2;    relay_conn far_1_1367_2_a(.in(far_1_1367_1[0]), .out(far_1_1367_2[0]));    relay_conn far_1_1367_2_b(.in(far_1_1367_1[1]), .out(far_1_1367_2[1]));
    assign layer_1[347] = far_1_1367_2[0] & far_1_1367_2[1]; 
    wire [1:0] far_1_1368_0;    relay_conn far_1_1368_0_a(.in(layer_0[362]), .out(far_1_1368_0[0]));    relay_conn far_1_1368_0_b(.in(layer_0[406]), .out(far_1_1368_0[1]));
    assign layer_1[348] = ~far_1_1368_0[1] | (far_1_1368_0[0] & far_1_1368_0[1]); 
    wire [1:0] far_1_1369_0;    relay_conn far_1_1369_0_a(.in(layer_0[356]), .out(far_1_1369_0[0]));    relay_conn far_1_1369_0_b(.in(layer_0[396]), .out(far_1_1369_0[1]));
    assign layer_1[349] = ~far_1_1369_0[0]; 
    wire [1:0] far_1_1370_0;    relay_conn far_1_1370_0_a(.in(layer_0[792]), .out(far_1_1370_0[0]));    relay_conn far_1_1370_0_b(.in(layer_0[879]), .out(far_1_1370_0[1]));
    wire [1:0] far_1_1370_1;    relay_conn far_1_1370_1_a(.in(far_1_1370_0[0]), .out(far_1_1370_1[0]));    relay_conn far_1_1370_1_b(.in(far_1_1370_0[1]), .out(far_1_1370_1[1]));
    assign layer_1[350] = far_1_1370_1[0] & far_1_1370_1[1]; 
    wire [1:0] far_1_1371_0;    relay_conn far_1_1371_0_a(.in(layer_0[966]), .out(far_1_1371_0[0]));    relay_conn far_1_1371_0_b(.in(layer_0[861]), .out(far_1_1371_0[1]));
    wire [1:0] far_1_1371_1;    relay_conn far_1_1371_1_a(.in(far_1_1371_0[0]), .out(far_1_1371_1[0]));    relay_conn far_1_1371_1_b(.in(far_1_1371_0[1]), .out(far_1_1371_1[1]));
    wire [1:0] far_1_1371_2;    relay_conn far_1_1371_2_a(.in(far_1_1371_1[0]), .out(far_1_1371_2[0]));    relay_conn far_1_1371_2_b(.in(far_1_1371_1[1]), .out(far_1_1371_2[1]));
    assign layer_1[351] = far_1_1371_2[0]; 
    wire [1:0] far_1_1372_0;    relay_conn far_1_1372_0_a(.in(layer_0[821]), .out(far_1_1372_0[0]));    relay_conn far_1_1372_0_b(.in(layer_0[773]), .out(far_1_1372_0[1]));
    assign layer_1[352] = ~(far_1_1372_0[0] | far_1_1372_0[1]); 
    assign layer_1[353] = ~layer_0[826] | (layer_0[855] & layer_0[826]); 
    wire [1:0] far_1_1374_0;    relay_conn far_1_1374_0_a(.in(layer_0[111]), .out(far_1_1374_0[0]));    relay_conn far_1_1374_0_b(.in(layer_0[14]), .out(far_1_1374_0[1]));
    wire [1:0] far_1_1374_1;    relay_conn far_1_1374_1_a(.in(far_1_1374_0[0]), .out(far_1_1374_1[0]));    relay_conn far_1_1374_1_b(.in(far_1_1374_0[1]), .out(far_1_1374_1[1]));
    wire [1:0] far_1_1374_2;    relay_conn far_1_1374_2_a(.in(far_1_1374_1[0]), .out(far_1_1374_2[0]));    relay_conn far_1_1374_2_b(.in(far_1_1374_1[1]), .out(far_1_1374_2[1]));
    assign layer_1[354] = ~far_1_1374_2[1]; 
    wire [1:0] far_1_1375_0;    relay_conn far_1_1375_0_a(.in(layer_0[242]), .out(far_1_1375_0[0]));    relay_conn far_1_1375_0_b(.in(layer_0[161]), .out(far_1_1375_0[1]));
    wire [1:0] far_1_1375_1;    relay_conn far_1_1375_1_a(.in(far_1_1375_0[0]), .out(far_1_1375_1[0]));    relay_conn far_1_1375_1_b(.in(far_1_1375_0[1]), .out(far_1_1375_1[1]));
    assign layer_1[355] = far_1_1375_1[0] | far_1_1375_1[1]; 
    wire [1:0] far_1_1376_0;    relay_conn far_1_1376_0_a(.in(layer_0[626]), .out(far_1_1376_0[0]));    relay_conn far_1_1376_0_b(.in(layer_0[544]), .out(far_1_1376_0[1]));
    wire [1:0] far_1_1376_1;    relay_conn far_1_1376_1_a(.in(far_1_1376_0[0]), .out(far_1_1376_1[0]));    relay_conn far_1_1376_1_b(.in(far_1_1376_0[1]), .out(far_1_1376_1[1]));
    assign layer_1[356] = ~far_1_1376_1[0]; 
    wire [1:0] far_1_1377_0;    relay_conn far_1_1377_0_a(.in(layer_0[403]), .out(far_1_1377_0[0]));    relay_conn far_1_1377_0_b(.in(layer_0[513]), .out(far_1_1377_0[1]));
    wire [1:0] far_1_1377_1;    relay_conn far_1_1377_1_a(.in(far_1_1377_0[0]), .out(far_1_1377_1[0]));    relay_conn far_1_1377_1_b(.in(far_1_1377_0[1]), .out(far_1_1377_1[1]));
    wire [1:0] far_1_1377_2;    relay_conn far_1_1377_2_a(.in(far_1_1377_1[0]), .out(far_1_1377_2[0]));    relay_conn far_1_1377_2_b(.in(far_1_1377_1[1]), .out(far_1_1377_2[1]));
    assign layer_1[357] = ~(far_1_1377_2[0] | far_1_1377_2[1]); 
    wire [1:0] far_1_1378_0;    relay_conn far_1_1378_0_a(.in(layer_0[281]), .out(far_1_1378_0[0]));    relay_conn far_1_1378_0_b(.in(layer_0[339]), .out(far_1_1378_0[1]));
    assign layer_1[358] = ~far_1_1378_0[1]; 
    assign layer_1[359] = ~layer_0[573]; 
    assign layer_1[360] = layer_0[57] | layer_0[75]; 
    assign layer_1[361] = layer_0[991] & ~layer_0[989]; 
    assign layer_1[362] = ~(layer_0[44] | layer_0[65]); 
    wire [1:0] far_1_1383_0;    relay_conn far_1_1383_0_a(.in(layer_0[964]), .out(far_1_1383_0[0]));    relay_conn far_1_1383_0_b(.in(layer_0[1004]), .out(far_1_1383_0[1]));
    assign layer_1[363] = far_1_1383_0[1] & ~far_1_1383_0[0]; 
    assign layer_1[364] = layer_0[448] | layer_0[419]; 
    wire [1:0] far_1_1385_0;    relay_conn far_1_1385_0_a(.in(layer_0[736]), .out(far_1_1385_0[0]));    relay_conn far_1_1385_0_b(.in(layer_0[799]), .out(far_1_1385_0[1]));
    assign layer_1[365] = far_1_1385_0[0] & ~far_1_1385_0[1]; 
    wire [1:0] far_1_1386_0;    relay_conn far_1_1386_0_a(.in(layer_0[65]), .out(far_1_1386_0[0]));    relay_conn far_1_1386_0_b(.in(layer_0[11]), .out(far_1_1386_0[1]));
    assign layer_1[366] = far_1_1386_0[0]; 
    wire [1:0] far_1_1387_0;    relay_conn far_1_1387_0_a(.in(layer_0[283]), .out(far_1_1387_0[0]));    relay_conn far_1_1387_0_b(.in(layer_0[337]), .out(far_1_1387_0[1]));
    assign layer_1[367] = ~(far_1_1387_0[0] & far_1_1387_0[1]); 
    wire [1:0] far_1_1388_0;    relay_conn far_1_1388_0_a(.in(layer_0[305]), .out(far_1_1388_0[0]));    relay_conn far_1_1388_0_b(.in(layer_0[243]), .out(far_1_1388_0[1]));
    assign layer_1[368] = ~(far_1_1388_0[0] | far_1_1388_0[1]); 
    assign layer_1[369] = ~layer_0[214] | (layer_0[214] & layer_0[187]); 
    wire [1:0] far_1_1390_0;    relay_conn far_1_1390_0_a(.in(layer_0[731]), .out(far_1_1390_0[0]));    relay_conn far_1_1390_0_b(.in(layer_0[855]), .out(far_1_1390_0[1]));
    wire [1:0] far_1_1390_1;    relay_conn far_1_1390_1_a(.in(far_1_1390_0[0]), .out(far_1_1390_1[0]));    relay_conn far_1_1390_1_b(.in(far_1_1390_0[1]), .out(far_1_1390_1[1]));
    wire [1:0] far_1_1390_2;    relay_conn far_1_1390_2_a(.in(far_1_1390_1[0]), .out(far_1_1390_2[0]));    relay_conn far_1_1390_2_b(.in(far_1_1390_1[1]), .out(far_1_1390_2[1]));
    assign layer_1[370] = ~(far_1_1390_2[0] ^ far_1_1390_2[1]); 
    assign layer_1[371] = layer_0[697] & layer_0[707]; 
    wire [1:0] far_1_1392_0;    relay_conn far_1_1392_0_a(.in(layer_0[507]), .out(far_1_1392_0[0]));    relay_conn far_1_1392_0_b(.in(layer_0[436]), .out(far_1_1392_0[1]));
    wire [1:0] far_1_1392_1;    relay_conn far_1_1392_1_a(.in(far_1_1392_0[0]), .out(far_1_1392_1[0]));    relay_conn far_1_1392_1_b(.in(far_1_1392_0[1]), .out(far_1_1392_1[1]));
    assign layer_1[372] = ~far_1_1392_1[0]; 
    assign layer_1[373] = layer_0[431]; 
    wire [1:0] far_1_1394_0;    relay_conn far_1_1394_0_a(.in(layer_0[43]), .out(far_1_1394_0[0]));    relay_conn far_1_1394_0_b(.in(layer_0[165]), .out(far_1_1394_0[1]));
    wire [1:0] far_1_1394_1;    relay_conn far_1_1394_1_a(.in(far_1_1394_0[0]), .out(far_1_1394_1[0]));    relay_conn far_1_1394_1_b(.in(far_1_1394_0[1]), .out(far_1_1394_1[1]));
    wire [1:0] far_1_1394_2;    relay_conn far_1_1394_2_a(.in(far_1_1394_1[0]), .out(far_1_1394_2[0]));    relay_conn far_1_1394_2_b(.in(far_1_1394_1[1]), .out(far_1_1394_2[1]));
    assign layer_1[374] = far_1_1394_2[0] & far_1_1394_2[1]; 
    wire [1:0] far_1_1395_0;    relay_conn far_1_1395_0_a(.in(layer_0[696]), .out(far_1_1395_0[0]));    relay_conn far_1_1395_0_b(.in(layer_0[798]), .out(far_1_1395_0[1]));
    wire [1:0] far_1_1395_1;    relay_conn far_1_1395_1_a(.in(far_1_1395_0[0]), .out(far_1_1395_1[0]));    relay_conn far_1_1395_1_b(.in(far_1_1395_0[1]), .out(far_1_1395_1[1]));
    wire [1:0] far_1_1395_2;    relay_conn far_1_1395_2_a(.in(far_1_1395_1[0]), .out(far_1_1395_2[0]));    relay_conn far_1_1395_2_b(.in(far_1_1395_1[1]), .out(far_1_1395_2[1]));
    assign layer_1[375] = ~far_1_1395_2[0] | (far_1_1395_2[0] & far_1_1395_2[1]); 
    wire [1:0] far_1_1396_0;    relay_conn far_1_1396_0_a(.in(layer_0[881]), .out(far_1_1396_0[0]));    relay_conn far_1_1396_0_b(.in(layer_0[1008]), .out(far_1_1396_0[1]));
    wire [1:0] far_1_1396_1;    relay_conn far_1_1396_1_a(.in(far_1_1396_0[0]), .out(far_1_1396_1[0]));    relay_conn far_1_1396_1_b(.in(far_1_1396_0[1]), .out(far_1_1396_1[1]));
    wire [1:0] far_1_1396_2;    relay_conn far_1_1396_2_a(.in(far_1_1396_1[0]), .out(far_1_1396_2[0]));    relay_conn far_1_1396_2_b(.in(far_1_1396_1[1]), .out(far_1_1396_2[1]));
    assign layer_1[376] = far_1_1396_2[1] & ~far_1_1396_2[0]; 
    wire [1:0] far_1_1397_0;    relay_conn far_1_1397_0_a(.in(layer_0[166]), .out(far_1_1397_0[0]));    relay_conn far_1_1397_0_b(.in(layer_0[66]), .out(far_1_1397_0[1]));
    wire [1:0] far_1_1397_1;    relay_conn far_1_1397_1_a(.in(far_1_1397_0[0]), .out(far_1_1397_1[0]));    relay_conn far_1_1397_1_b(.in(far_1_1397_0[1]), .out(far_1_1397_1[1]));
    wire [1:0] far_1_1397_2;    relay_conn far_1_1397_2_a(.in(far_1_1397_1[0]), .out(far_1_1397_2[0]));    relay_conn far_1_1397_2_b(.in(far_1_1397_1[1]), .out(far_1_1397_2[1]));
    assign layer_1[377] = ~far_1_1397_2[0]; 
    wire [1:0] far_1_1398_0;    relay_conn far_1_1398_0_a(.in(layer_0[143]), .out(far_1_1398_0[0]));    relay_conn far_1_1398_0_b(.in(layer_0[93]), .out(far_1_1398_0[1]));
    assign layer_1[378] = ~(far_1_1398_0[0] & far_1_1398_0[1]); 
    wire [1:0] far_1_1399_0;    relay_conn far_1_1399_0_a(.in(layer_0[651]), .out(far_1_1399_0[0]));    relay_conn far_1_1399_0_b(.in(layer_0[573]), .out(far_1_1399_0[1]));
    wire [1:0] far_1_1399_1;    relay_conn far_1_1399_1_a(.in(far_1_1399_0[0]), .out(far_1_1399_1[0]));    relay_conn far_1_1399_1_b(.in(far_1_1399_0[1]), .out(far_1_1399_1[1]));
    assign layer_1[379] = ~far_1_1399_1[1]; 
    wire [1:0] far_1_1400_0;    relay_conn far_1_1400_0_a(.in(layer_0[547]), .out(far_1_1400_0[0]));    relay_conn far_1_1400_0_b(.in(layer_0[588]), .out(far_1_1400_0[1]));
    assign layer_1[380] = far_1_1400_0[0] ^ far_1_1400_0[1]; 
    assign layer_1[381] = layer_0[32] & ~layer_0[30]; 
    wire [1:0] far_1_1402_0;    relay_conn far_1_1402_0_a(.in(layer_0[243]), .out(far_1_1402_0[0]));    relay_conn far_1_1402_0_b(.in(layer_0[283]), .out(far_1_1402_0[1]));
    assign layer_1[382] = far_1_1402_0[1] & ~far_1_1402_0[0]; 
    assign layer_1[383] = layer_0[461]; 
    wire [1:0] far_1_1404_0;    relay_conn far_1_1404_0_a(.in(layer_0[685]), .out(far_1_1404_0[0]));    relay_conn far_1_1404_0_b(.in(layer_0[559]), .out(far_1_1404_0[1]));
    wire [1:0] far_1_1404_1;    relay_conn far_1_1404_1_a(.in(far_1_1404_0[0]), .out(far_1_1404_1[0]));    relay_conn far_1_1404_1_b(.in(far_1_1404_0[1]), .out(far_1_1404_1[1]));
    wire [1:0] far_1_1404_2;    relay_conn far_1_1404_2_a(.in(far_1_1404_1[0]), .out(far_1_1404_2[0]));    relay_conn far_1_1404_2_b(.in(far_1_1404_1[1]), .out(far_1_1404_2[1]));
    assign layer_1[384] = far_1_1404_2[1] & ~far_1_1404_2[0]; 
    wire [1:0] far_1_1405_0;    relay_conn far_1_1405_0_a(.in(layer_0[162]), .out(far_1_1405_0[0]));    relay_conn far_1_1405_0_b(.in(layer_0[251]), .out(far_1_1405_0[1]));
    wire [1:0] far_1_1405_1;    relay_conn far_1_1405_1_a(.in(far_1_1405_0[0]), .out(far_1_1405_1[0]));    relay_conn far_1_1405_1_b(.in(far_1_1405_0[1]), .out(far_1_1405_1[1]));
    assign layer_1[385] = far_1_1405_1[0] & ~far_1_1405_1[1]; 
    assign layer_1[386] = ~layer_0[1014]; 
    assign layer_1[387] = ~layer_0[408] | (layer_0[408] & layer_0[438]); 
    assign layer_1[388] = layer_0[348]; 
    wire [1:0] far_1_1409_0;    relay_conn far_1_1409_0_a(.in(layer_0[313]), .out(far_1_1409_0[0]));    relay_conn far_1_1409_0_b(.in(layer_0[185]), .out(far_1_1409_0[1]));
    wire [1:0] far_1_1409_1;    relay_conn far_1_1409_1_a(.in(far_1_1409_0[0]), .out(far_1_1409_1[0]));    relay_conn far_1_1409_1_b(.in(far_1_1409_0[1]), .out(far_1_1409_1[1]));
    wire [1:0] far_1_1409_2;    relay_conn far_1_1409_2_a(.in(far_1_1409_1[0]), .out(far_1_1409_2[0]));    relay_conn far_1_1409_2_b(.in(far_1_1409_1[1]), .out(far_1_1409_2[1]));
    wire [1:0] far_1_1409_3;    relay_conn far_1_1409_3_a(.in(far_1_1409_2[0]), .out(far_1_1409_3[0]));    relay_conn far_1_1409_3_b(.in(far_1_1409_2[1]), .out(far_1_1409_3[1]));
    assign layer_1[389] = ~far_1_1409_3[1]; 
    wire [1:0] far_1_1410_0;    relay_conn far_1_1410_0_a(.in(layer_0[873]), .out(far_1_1410_0[0]));    relay_conn far_1_1410_0_b(.in(layer_0[978]), .out(far_1_1410_0[1]));
    wire [1:0] far_1_1410_1;    relay_conn far_1_1410_1_a(.in(far_1_1410_0[0]), .out(far_1_1410_1[0]));    relay_conn far_1_1410_1_b(.in(far_1_1410_0[1]), .out(far_1_1410_1[1]));
    wire [1:0] far_1_1410_2;    relay_conn far_1_1410_2_a(.in(far_1_1410_1[0]), .out(far_1_1410_2[0]));    relay_conn far_1_1410_2_b(.in(far_1_1410_1[1]), .out(far_1_1410_2[1]));
    assign layer_1[390] = far_1_1410_2[0] & far_1_1410_2[1]; 
    wire [1:0] far_1_1411_0;    relay_conn far_1_1411_0_a(.in(layer_0[489]), .out(far_1_1411_0[0]));    relay_conn far_1_1411_0_b(.in(layer_0[614]), .out(far_1_1411_0[1]));
    wire [1:0] far_1_1411_1;    relay_conn far_1_1411_1_a(.in(far_1_1411_0[0]), .out(far_1_1411_1[0]));    relay_conn far_1_1411_1_b(.in(far_1_1411_0[1]), .out(far_1_1411_1[1]));
    wire [1:0] far_1_1411_2;    relay_conn far_1_1411_2_a(.in(far_1_1411_1[0]), .out(far_1_1411_2[0]));    relay_conn far_1_1411_2_b(.in(far_1_1411_1[1]), .out(far_1_1411_2[1]));
    assign layer_1[391] = far_1_1411_2[0] & ~far_1_1411_2[1]; 
    wire [1:0] far_1_1412_0;    relay_conn far_1_1412_0_a(.in(layer_0[380]), .out(far_1_1412_0[0]));    relay_conn far_1_1412_0_b(.in(layer_0[322]), .out(far_1_1412_0[1]));
    assign layer_1[392] = far_1_1412_0[0] & ~far_1_1412_0[1]; 
    wire [1:0] far_1_1413_0;    relay_conn far_1_1413_0_a(.in(layer_0[148]), .out(far_1_1413_0[0]));    relay_conn far_1_1413_0_b(.in(layer_0[71]), .out(far_1_1413_0[1]));
    wire [1:0] far_1_1413_1;    relay_conn far_1_1413_1_a(.in(far_1_1413_0[0]), .out(far_1_1413_1[0]));    relay_conn far_1_1413_1_b(.in(far_1_1413_0[1]), .out(far_1_1413_1[1]));
    assign layer_1[393] = ~far_1_1413_1[0] | (far_1_1413_1[0] & far_1_1413_1[1]); 
    wire [1:0] far_1_1414_0;    relay_conn far_1_1414_0_a(.in(layer_0[192]), .out(far_1_1414_0[0]));    relay_conn far_1_1414_0_b(.in(layer_0[285]), .out(far_1_1414_0[1]));
    wire [1:0] far_1_1414_1;    relay_conn far_1_1414_1_a(.in(far_1_1414_0[0]), .out(far_1_1414_1[0]));    relay_conn far_1_1414_1_b(.in(far_1_1414_0[1]), .out(far_1_1414_1[1]));
    assign layer_1[394] = ~far_1_1414_1[0] | (far_1_1414_1[0] & far_1_1414_1[1]); 
    wire [1:0] far_1_1415_0;    relay_conn far_1_1415_0_a(.in(layer_0[313]), .out(far_1_1415_0[0]));    relay_conn far_1_1415_0_b(.in(layer_0[210]), .out(far_1_1415_0[1]));
    wire [1:0] far_1_1415_1;    relay_conn far_1_1415_1_a(.in(far_1_1415_0[0]), .out(far_1_1415_1[0]));    relay_conn far_1_1415_1_b(.in(far_1_1415_0[1]), .out(far_1_1415_1[1]));
    wire [1:0] far_1_1415_2;    relay_conn far_1_1415_2_a(.in(far_1_1415_1[0]), .out(far_1_1415_2[0]));    relay_conn far_1_1415_2_b(.in(far_1_1415_1[1]), .out(far_1_1415_2[1]));
    assign layer_1[395] = ~(far_1_1415_2[0] ^ far_1_1415_2[1]); 
    wire [1:0] far_1_1416_0;    relay_conn far_1_1416_0_a(.in(layer_0[272]), .out(far_1_1416_0[0]));    relay_conn far_1_1416_0_b(.in(layer_0[237]), .out(far_1_1416_0[1]));
    assign layer_1[396] = far_1_1416_0[0] | far_1_1416_0[1]; 
    assign layer_1[397] = layer_0[389] & ~layer_0[367]; 
    wire [1:0] far_1_1418_0;    relay_conn far_1_1418_0_a(.in(layer_0[1009]), .out(far_1_1418_0[0]));    relay_conn far_1_1418_0_b(.in(layer_0[896]), .out(far_1_1418_0[1]));
    wire [1:0] far_1_1418_1;    relay_conn far_1_1418_1_a(.in(far_1_1418_0[0]), .out(far_1_1418_1[0]));    relay_conn far_1_1418_1_b(.in(far_1_1418_0[1]), .out(far_1_1418_1[1]));
    wire [1:0] far_1_1418_2;    relay_conn far_1_1418_2_a(.in(far_1_1418_1[0]), .out(far_1_1418_2[0]));    relay_conn far_1_1418_2_b(.in(far_1_1418_1[1]), .out(far_1_1418_2[1]));
    assign layer_1[398] = far_1_1418_2[0] | far_1_1418_2[1]; 
    wire [1:0] far_1_1419_0;    relay_conn far_1_1419_0_a(.in(layer_0[564]), .out(far_1_1419_0[0]));    relay_conn far_1_1419_0_b(.in(layer_0[446]), .out(far_1_1419_0[1]));
    wire [1:0] far_1_1419_1;    relay_conn far_1_1419_1_a(.in(far_1_1419_0[0]), .out(far_1_1419_1[0]));    relay_conn far_1_1419_1_b(.in(far_1_1419_0[1]), .out(far_1_1419_1[1]));
    wire [1:0] far_1_1419_2;    relay_conn far_1_1419_2_a(.in(far_1_1419_1[0]), .out(far_1_1419_2[0]));    relay_conn far_1_1419_2_b(.in(far_1_1419_1[1]), .out(far_1_1419_2[1]));
    assign layer_1[399] = ~far_1_1419_2[0]; 
    wire [1:0] far_1_1420_0;    relay_conn far_1_1420_0_a(.in(layer_0[1017]), .out(far_1_1420_0[0]));    relay_conn far_1_1420_0_b(.in(layer_0[891]), .out(far_1_1420_0[1]));
    wire [1:0] far_1_1420_1;    relay_conn far_1_1420_1_a(.in(far_1_1420_0[0]), .out(far_1_1420_1[0]));    relay_conn far_1_1420_1_b(.in(far_1_1420_0[1]), .out(far_1_1420_1[1]));
    wire [1:0] far_1_1420_2;    relay_conn far_1_1420_2_a(.in(far_1_1420_1[0]), .out(far_1_1420_2[0]));    relay_conn far_1_1420_2_b(.in(far_1_1420_1[1]), .out(far_1_1420_2[1]));
    assign layer_1[400] = far_1_1420_2[0] & ~far_1_1420_2[1]; 
    wire [1:0] far_1_1421_0;    relay_conn far_1_1421_0_a(.in(layer_0[836]), .out(far_1_1421_0[0]));    relay_conn far_1_1421_0_b(.in(layer_0[786]), .out(far_1_1421_0[1]));
    assign layer_1[401] = far_1_1421_0[0] & ~far_1_1421_0[1]; 
    wire [1:0] far_1_1422_0;    relay_conn far_1_1422_0_a(.in(layer_0[983]), .out(far_1_1422_0[0]));    relay_conn far_1_1422_0_b(.in(layer_0[937]), .out(far_1_1422_0[1]));
    assign layer_1[402] = far_1_1422_0[1] & ~far_1_1422_0[0]; 
    wire [1:0] far_1_1423_0;    relay_conn far_1_1423_0_a(.in(layer_0[810]), .out(far_1_1423_0[0]));    relay_conn far_1_1423_0_b(.in(layer_0[856]), .out(far_1_1423_0[1]));
    assign layer_1[403] = far_1_1423_0[1] & ~far_1_1423_0[0]; 
    wire [1:0] far_1_1424_0;    relay_conn far_1_1424_0_a(.in(layer_0[785]), .out(far_1_1424_0[0]));    relay_conn far_1_1424_0_b(.in(layer_0[896]), .out(far_1_1424_0[1]));
    wire [1:0] far_1_1424_1;    relay_conn far_1_1424_1_a(.in(far_1_1424_0[0]), .out(far_1_1424_1[0]));    relay_conn far_1_1424_1_b(.in(far_1_1424_0[1]), .out(far_1_1424_1[1]));
    wire [1:0] far_1_1424_2;    relay_conn far_1_1424_2_a(.in(far_1_1424_1[0]), .out(far_1_1424_2[0]));    relay_conn far_1_1424_2_b(.in(far_1_1424_1[1]), .out(far_1_1424_2[1]));
    assign layer_1[404] = ~far_1_1424_2[0] | (far_1_1424_2[0] & far_1_1424_2[1]); 
    wire [1:0] far_1_1425_0;    relay_conn far_1_1425_0_a(.in(layer_0[676]), .out(far_1_1425_0[0]));    relay_conn far_1_1425_0_b(.in(layer_0[734]), .out(far_1_1425_0[1]));
    assign layer_1[405] = ~far_1_1425_0[0] | (far_1_1425_0[0] & far_1_1425_0[1]); 
    assign layer_1[406] = layer_0[334]; 
    assign layer_1[407] = ~(layer_0[923] | layer_0[899]); 
    wire [1:0] far_1_1428_0;    relay_conn far_1_1428_0_a(.in(layer_0[30]), .out(far_1_1428_0[0]));    relay_conn far_1_1428_0_b(.in(layer_0[147]), .out(far_1_1428_0[1]));
    wire [1:0] far_1_1428_1;    relay_conn far_1_1428_1_a(.in(far_1_1428_0[0]), .out(far_1_1428_1[0]));    relay_conn far_1_1428_1_b(.in(far_1_1428_0[1]), .out(far_1_1428_1[1]));
    wire [1:0] far_1_1428_2;    relay_conn far_1_1428_2_a(.in(far_1_1428_1[0]), .out(far_1_1428_2[0]));    relay_conn far_1_1428_2_b(.in(far_1_1428_1[1]), .out(far_1_1428_2[1]));
    assign layer_1[408] = ~far_1_1428_2[1] | (far_1_1428_2[0] & far_1_1428_2[1]); 
    wire [1:0] far_1_1429_0;    relay_conn far_1_1429_0_a(.in(layer_0[67]), .out(far_1_1429_0[0]));    relay_conn far_1_1429_0_b(.in(layer_0[19]), .out(far_1_1429_0[1]));
    assign layer_1[409] = ~far_1_1429_0[0]; 
    wire [1:0] far_1_1430_0;    relay_conn far_1_1430_0_a(.in(layer_0[256]), .out(far_1_1430_0[0]));    relay_conn far_1_1430_0_b(.in(layer_0[337]), .out(far_1_1430_0[1]));
    wire [1:0] far_1_1430_1;    relay_conn far_1_1430_1_a(.in(far_1_1430_0[0]), .out(far_1_1430_1[0]));    relay_conn far_1_1430_1_b(.in(far_1_1430_0[1]), .out(far_1_1430_1[1]));
    assign layer_1[410] = far_1_1430_1[0] | far_1_1430_1[1]; 
    assign layer_1[411] = ~(layer_0[644] | layer_0[628]); 
    wire [1:0] far_1_1432_0;    relay_conn far_1_1432_0_a(.in(layer_0[961]), .out(far_1_1432_0[0]));    relay_conn far_1_1432_0_b(.in(layer_0[845]), .out(far_1_1432_0[1]));
    wire [1:0] far_1_1432_1;    relay_conn far_1_1432_1_a(.in(far_1_1432_0[0]), .out(far_1_1432_1[0]));    relay_conn far_1_1432_1_b(.in(far_1_1432_0[1]), .out(far_1_1432_1[1]));
    wire [1:0] far_1_1432_2;    relay_conn far_1_1432_2_a(.in(far_1_1432_1[0]), .out(far_1_1432_2[0]));    relay_conn far_1_1432_2_b(.in(far_1_1432_1[1]), .out(far_1_1432_2[1]));
    assign layer_1[412] = ~(far_1_1432_2[0] & far_1_1432_2[1]); 
    assign layer_1[413] = layer_0[933] ^ layer_0[954]; 
    wire [1:0] far_1_1434_0;    relay_conn far_1_1434_0_a(.in(layer_0[672]), .out(far_1_1434_0[0]));    relay_conn far_1_1434_0_b(.in(layer_0[590]), .out(far_1_1434_0[1]));
    wire [1:0] far_1_1434_1;    relay_conn far_1_1434_1_a(.in(far_1_1434_0[0]), .out(far_1_1434_1[0]));    relay_conn far_1_1434_1_b(.in(far_1_1434_0[1]), .out(far_1_1434_1[1]));
    assign layer_1[414] = ~(far_1_1434_1[0] | far_1_1434_1[1]); 
    wire [1:0] far_1_1435_0;    relay_conn far_1_1435_0_a(.in(layer_0[853]), .out(far_1_1435_0[0]));    relay_conn far_1_1435_0_b(.in(layer_0[773]), .out(far_1_1435_0[1]));
    wire [1:0] far_1_1435_1;    relay_conn far_1_1435_1_a(.in(far_1_1435_0[0]), .out(far_1_1435_1[0]));    relay_conn far_1_1435_1_b(.in(far_1_1435_0[1]), .out(far_1_1435_1[1]));
    assign layer_1[415] = far_1_1435_1[0] & far_1_1435_1[1]; 
    assign layer_1[416] = ~layer_0[475] | (layer_0[475] & layer_0[451]); 
    wire [1:0] far_1_1437_0;    relay_conn far_1_1437_0_a(.in(layer_0[706]), .out(far_1_1437_0[0]));    relay_conn far_1_1437_0_b(.in(layer_0[741]), .out(far_1_1437_0[1]));
    assign layer_1[417] = far_1_1437_0[0]; 
    wire [1:0] far_1_1438_0;    relay_conn far_1_1438_0_a(.in(layer_0[699]), .out(far_1_1438_0[0]));    relay_conn far_1_1438_0_b(.in(layer_0[748]), .out(far_1_1438_0[1]));
    assign layer_1[418] = ~far_1_1438_0[1] | (far_1_1438_0[0] & far_1_1438_0[1]); 
    wire [1:0] far_1_1439_0;    relay_conn far_1_1439_0_a(.in(layer_0[816]), .out(far_1_1439_0[0]));    relay_conn far_1_1439_0_b(.in(layer_0[914]), .out(far_1_1439_0[1]));
    wire [1:0] far_1_1439_1;    relay_conn far_1_1439_1_a(.in(far_1_1439_0[0]), .out(far_1_1439_1[0]));    relay_conn far_1_1439_1_b(.in(far_1_1439_0[1]), .out(far_1_1439_1[1]));
    wire [1:0] far_1_1439_2;    relay_conn far_1_1439_2_a(.in(far_1_1439_1[0]), .out(far_1_1439_2[0]));    relay_conn far_1_1439_2_b(.in(far_1_1439_1[1]), .out(far_1_1439_2[1]));
    assign layer_1[419] = far_1_1439_2[1]; 
    assign layer_1[420] = layer_0[412] & ~layer_0[396]; 
    assign layer_1[421] = ~layer_0[590] | (layer_0[590] & layer_0[592]); 
    assign layer_1[422] = layer_0[401]; 
    wire [1:0] far_1_1443_0;    relay_conn far_1_1443_0_a(.in(layer_0[395]), .out(far_1_1443_0[0]));    relay_conn far_1_1443_0_b(.in(layer_0[330]), .out(far_1_1443_0[1]));
    wire [1:0] far_1_1443_1;    relay_conn far_1_1443_1_a(.in(far_1_1443_0[0]), .out(far_1_1443_1[0]));    relay_conn far_1_1443_1_b(.in(far_1_1443_0[1]), .out(far_1_1443_1[1]));
    assign layer_1[423] = far_1_1443_1[1] & ~far_1_1443_1[0]; 
    wire [1:0] far_1_1444_0;    relay_conn far_1_1444_0_a(.in(layer_0[752]), .out(far_1_1444_0[0]));    relay_conn far_1_1444_0_b(.in(layer_0[708]), .out(far_1_1444_0[1]));
    assign layer_1[424] = far_1_1444_0[0] & far_1_1444_0[1]; 
    wire [1:0] far_1_1445_0;    relay_conn far_1_1445_0_a(.in(layer_0[607]), .out(far_1_1445_0[0]));    relay_conn far_1_1445_0_b(.in(layer_0[656]), .out(far_1_1445_0[1]));
    assign layer_1[425] = ~(far_1_1445_0[0] | far_1_1445_0[1]); 
    wire [1:0] far_1_1446_0;    relay_conn far_1_1446_0_a(.in(layer_0[886]), .out(far_1_1446_0[0]));    relay_conn far_1_1446_0_b(.in(layer_0[768]), .out(far_1_1446_0[1]));
    wire [1:0] far_1_1446_1;    relay_conn far_1_1446_1_a(.in(far_1_1446_0[0]), .out(far_1_1446_1[0]));    relay_conn far_1_1446_1_b(.in(far_1_1446_0[1]), .out(far_1_1446_1[1]));
    wire [1:0] far_1_1446_2;    relay_conn far_1_1446_2_a(.in(far_1_1446_1[0]), .out(far_1_1446_2[0]));    relay_conn far_1_1446_2_b(.in(far_1_1446_1[1]), .out(far_1_1446_2[1]));
    assign layer_1[426] = far_1_1446_2[1] & ~far_1_1446_2[0]; 
    assign layer_1[427] = layer_0[697]; 
    wire [1:0] far_1_1448_0;    relay_conn far_1_1448_0_a(.in(layer_0[395]), .out(far_1_1448_0[0]));    relay_conn far_1_1448_0_b(.in(layer_0[475]), .out(far_1_1448_0[1]));
    wire [1:0] far_1_1448_1;    relay_conn far_1_1448_1_a(.in(far_1_1448_0[0]), .out(far_1_1448_1[0]));    relay_conn far_1_1448_1_b(.in(far_1_1448_0[1]), .out(far_1_1448_1[1]));
    assign layer_1[428] = far_1_1448_1[0]; 
    wire [1:0] far_1_1449_0;    relay_conn far_1_1449_0_a(.in(layer_0[204]), .out(far_1_1449_0[0]));    relay_conn far_1_1449_0_b(.in(layer_0[124]), .out(far_1_1449_0[1]));
    wire [1:0] far_1_1449_1;    relay_conn far_1_1449_1_a(.in(far_1_1449_0[0]), .out(far_1_1449_1[0]));    relay_conn far_1_1449_1_b(.in(far_1_1449_0[1]), .out(far_1_1449_1[1]));
    assign layer_1[429] = ~far_1_1449_1[1]; 
    wire [1:0] far_1_1450_0;    relay_conn far_1_1450_0_a(.in(layer_0[974]), .out(far_1_1450_0[0]));    relay_conn far_1_1450_0_b(.in(layer_0[852]), .out(far_1_1450_0[1]));
    wire [1:0] far_1_1450_1;    relay_conn far_1_1450_1_a(.in(far_1_1450_0[0]), .out(far_1_1450_1[0]));    relay_conn far_1_1450_1_b(.in(far_1_1450_0[1]), .out(far_1_1450_1[1]));
    wire [1:0] far_1_1450_2;    relay_conn far_1_1450_2_a(.in(far_1_1450_1[0]), .out(far_1_1450_2[0]));    relay_conn far_1_1450_2_b(.in(far_1_1450_1[1]), .out(far_1_1450_2[1]));
    assign layer_1[430] = ~(far_1_1450_2[0] | far_1_1450_2[1]); 
    assign layer_1[431] = layer_0[237]; 
    wire [1:0] far_1_1452_0;    relay_conn far_1_1452_0_a(.in(layer_0[422]), .out(far_1_1452_0[0]));    relay_conn far_1_1452_0_b(.in(layer_0[372]), .out(far_1_1452_0[1]));
    assign layer_1[432] = ~far_1_1452_0[1] | (far_1_1452_0[0] & far_1_1452_0[1]); 
    wire [1:0] far_1_1453_0;    relay_conn far_1_1453_0_a(.in(layer_0[237]), .out(far_1_1453_0[0]));    relay_conn far_1_1453_0_b(.in(layer_0[347]), .out(far_1_1453_0[1]));
    wire [1:0] far_1_1453_1;    relay_conn far_1_1453_1_a(.in(far_1_1453_0[0]), .out(far_1_1453_1[0]));    relay_conn far_1_1453_1_b(.in(far_1_1453_0[1]), .out(far_1_1453_1[1]));
    wire [1:0] far_1_1453_2;    relay_conn far_1_1453_2_a(.in(far_1_1453_1[0]), .out(far_1_1453_2[0]));    relay_conn far_1_1453_2_b(.in(far_1_1453_1[1]), .out(far_1_1453_2[1]));
    assign layer_1[433] = ~(far_1_1453_2[0] | far_1_1453_2[1]); 
    assign layer_1[434] = ~(layer_0[367] ^ layer_0[346]); 
    assign layer_1[435] = ~layer_0[395]; 
    wire [1:0] far_1_1456_0;    relay_conn far_1_1456_0_a(.in(layer_0[379]), .out(far_1_1456_0[0]));    relay_conn far_1_1456_0_b(.in(layer_0[256]), .out(far_1_1456_0[1]));
    wire [1:0] far_1_1456_1;    relay_conn far_1_1456_1_a(.in(far_1_1456_0[0]), .out(far_1_1456_1[0]));    relay_conn far_1_1456_1_b(.in(far_1_1456_0[1]), .out(far_1_1456_1[1]));
    wire [1:0] far_1_1456_2;    relay_conn far_1_1456_2_a(.in(far_1_1456_1[0]), .out(far_1_1456_2[0]));    relay_conn far_1_1456_2_b(.in(far_1_1456_1[1]), .out(far_1_1456_2[1]));
    assign layer_1[436] = ~far_1_1456_2[1] | (far_1_1456_2[0] & far_1_1456_2[1]); 
    wire [1:0] far_1_1457_0;    relay_conn far_1_1457_0_a(.in(layer_0[338]), .out(far_1_1457_0[0]));    relay_conn far_1_1457_0_b(.in(layer_0[391]), .out(far_1_1457_0[1]));
    assign layer_1[437] = far_1_1457_0[0] | far_1_1457_0[1]; 
    wire [1:0] far_1_1458_0;    relay_conn far_1_1458_0_a(.in(layer_0[506]), .out(far_1_1458_0[0]));    relay_conn far_1_1458_0_b(.in(layer_0[444]), .out(far_1_1458_0[1]));
    assign layer_1[438] = ~(far_1_1458_0[0] & far_1_1458_0[1]); 
    wire [1:0] far_1_1459_0;    relay_conn far_1_1459_0_a(.in(layer_0[807]), .out(far_1_1459_0[0]));    relay_conn far_1_1459_0_b(.in(layer_0[931]), .out(far_1_1459_0[1]));
    wire [1:0] far_1_1459_1;    relay_conn far_1_1459_1_a(.in(far_1_1459_0[0]), .out(far_1_1459_1[0]));    relay_conn far_1_1459_1_b(.in(far_1_1459_0[1]), .out(far_1_1459_1[1]));
    wire [1:0] far_1_1459_2;    relay_conn far_1_1459_2_a(.in(far_1_1459_1[0]), .out(far_1_1459_2[0]));    relay_conn far_1_1459_2_b(.in(far_1_1459_1[1]), .out(far_1_1459_2[1]));
    assign layer_1[439] = far_1_1459_2[0]; 
    wire [1:0] far_1_1460_0;    relay_conn far_1_1460_0_a(.in(layer_0[339]), .out(far_1_1460_0[0]));    relay_conn far_1_1460_0_b(.in(layer_0[454]), .out(far_1_1460_0[1]));
    wire [1:0] far_1_1460_1;    relay_conn far_1_1460_1_a(.in(far_1_1460_0[0]), .out(far_1_1460_1[0]));    relay_conn far_1_1460_1_b(.in(far_1_1460_0[1]), .out(far_1_1460_1[1]));
    wire [1:0] far_1_1460_2;    relay_conn far_1_1460_2_a(.in(far_1_1460_1[0]), .out(far_1_1460_2[0]));    relay_conn far_1_1460_2_b(.in(far_1_1460_1[1]), .out(far_1_1460_2[1]));
    assign layer_1[440] = ~far_1_1460_2[0] | (far_1_1460_2[0] & far_1_1460_2[1]); 
    wire [1:0] far_1_1461_0;    relay_conn far_1_1461_0_a(.in(layer_0[988]), .out(far_1_1461_0[0]));    relay_conn far_1_1461_0_b(.in(layer_0[916]), .out(far_1_1461_0[1]));
    wire [1:0] far_1_1461_1;    relay_conn far_1_1461_1_a(.in(far_1_1461_0[0]), .out(far_1_1461_1[0]));    relay_conn far_1_1461_1_b(.in(far_1_1461_0[1]), .out(far_1_1461_1[1]));
    assign layer_1[441] = far_1_1461_1[1] & ~far_1_1461_1[0]; 
    wire [1:0] far_1_1462_0;    relay_conn far_1_1462_0_a(.in(layer_0[865]), .out(far_1_1462_0[0]));    relay_conn far_1_1462_0_b(.in(layer_0[827]), .out(far_1_1462_0[1]));
    assign layer_1[442] = far_1_1462_0[0] & ~far_1_1462_0[1]; 
    wire [1:0] far_1_1463_0;    relay_conn far_1_1463_0_a(.in(layer_0[214]), .out(far_1_1463_0[0]));    relay_conn far_1_1463_0_b(.in(layer_0[121]), .out(far_1_1463_0[1]));
    wire [1:0] far_1_1463_1;    relay_conn far_1_1463_1_a(.in(far_1_1463_0[0]), .out(far_1_1463_1[0]));    relay_conn far_1_1463_1_b(.in(far_1_1463_0[1]), .out(far_1_1463_1[1]));
    assign layer_1[443] = far_1_1463_1[0]; 
    assign layer_1[444] = ~(layer_0[647] | layer_0[621]); 
    wire [1:0] far_1_1465_0;    relay_conn far_1_1465_0_a(.in(layer_0[871]), .out(far_1_1465_0[0]));    relay_conn far_1_1465_0_b(.in(layer_0[985]), .out(far_1_1465_0[1]));
    wire [1:0] far_1_1465_1;    relay_conn far_1_1465_1_a(.in(far_1_1465_0[0]), .out(far_1_1465_1[0]));    relay_conn far_1_1465_1_b(.in(far_1_1465_0[1]), .out(far_1_1465_1[1]));
    wire [1:0] far_1_1465_2;    relay_conn far_1_1465_2_a(.in(far_1_1465_1[0]), .out(far_1_1465_2[0]));    relay_conn far_1_1465_2_b(.in(far_1_1465_1[1]), .out(far_1_1465_2[1]));
    assign layer_1[445] = ~far_1_1465_2[0] | (far_1_1465_2[0] & far_1_1465_2[1]); 
    wire [1:0] far_1_1466_0;    relay_conn far_1_1466_0_a(.in(layer_0[841]), .out(far_1_1466_0[0]));    relay_conn far_1_1466_0_b(.in(layer_0[888]), .out(far_1_1466_0[1]));
    assign layer_1[446] = far_1_1466_0[0] & far_1_1466_0[1]; 
    wire [1:0] far_1_1467_0;    relay_conn far_1_1467_0_a(.in(layer_0[543]), .out(far_1_1467_0[0]));    relay_conn far_1_1467_0_b(.in(layer_0[430]), .out(far_1_1467_0[1]));
    wire [1:0] far_1_1467_1;    relay_conn far_1_1467_1_a(.in(far_1_1467_0[0]), .out(far_1_1467_1[0]));    relay_conn far_1_1467_1_b(.in(far_1_1467_0[1]), .out(far_1_1467_1[1]));
    wire [1:0] far_1_1467_2;    relay_conn far_1_1467_2_a(.in(far_1_1467_1[0]), .out(far_1_1467_2[0]));    relay_conn far_1_1467_2_b(.in(far_1_1467_1[1]), .out(far_1_1467_2[1]));
    assign layer_1[447] = ~(far_1_1467_2[0] ^ far_1_1467_2[1]); 
    assign layer_1[448] = layer_0[954] & layer_0[964]; 
    wire [1:0] far_1_1469_0;    relay_conn far_1_1469_0_a(.in(layer_0[768]), .out(far_1_1469_0[0]));    relay_conn far_1_1469_0_b(.in(layer_0[707]), .out(far_1_1469_0[1]));
    assign layer_1[449] = ~(far_1_1469_0[0] ^ far_1_1469_0[1]); 
    assign layer_1[450] = ~(layer_0[257] ^ layer_0[240]); 
    wire [1:0] far_1_1471_0;    relay_conn far_1_1471_0_a(.in(layer_0[277]), .out(far_1_1471_0[0]));    relay_conn far_1_1471_0_b(.in(layer_0[208]), .out(far_1_1471_0[1]));
    wire [1:0] far_1_1471_1;    relay_conn far_1_1471_1_a(.in(far_1_1471_0[0]), .out(far_1_1471_1[0]));    relay_conn far_1_1471_1_b(.in(far_1_1471_0[1]), .out(far_1_1471_1[1]));
    assign layer_1[451] = ~far_1_1471_1[1]; 
    wire [1:0] far_1_1472_0;    relay_conn far_1_1472_0_a(.in(layer_0[926]), .out(far_1_1472_0[0]));    relay_conn far_1_1472_0_b(.in(layer_0[984]), .out(far_1_1472_0[1]));
    assign layer_1[452] = far_1_1472_0[1] & ~far_1_1472_0[0]; 
    wire [1:0] far_1_1473_0;    relay_conn far_1_1473_0_a(.in(layer_0[676]), .out(far_1_1473_0[0]));    relay_conn far_1_1473_0_b(.in(layer_0[590]), .out(far_1_1473_0[1]));
    wire [1:0] far_1_1473_1;    relay_conn far_1_1473_1_a(.in(far_1_1473_0[0]), .out(far_1_1473_1[0]));    relay_conn far_1_1473_1_b(.in(far_1_1473_0[1]), .out(far_1_1473_1[1]));
    assign layer_1[453] = far_1_1473_1[1]; 
    wire [1:0] far_1_1474_0;    relay_conn far_1_1474_0_a(.in(layer_0[954]), .out(far_1_1474_0[0]));    relay_conn far_1_1474_0_b(.in(layer_0[841]), .out(far_1_1474_0[1]));
    wire [1:0] far_1_1474_1;    relay_conn far_1_1474_1_a(.in(far_1_1474_0[0]), .out(far_1_1474_1[0]));    relay_conn far_1_1474_1_b(.in(far_1_1474_0[1]), .out(far_1_1474_1[1]));
    wire [1:0] far_1_1474_2;    relay_conn far_1_1474_2_a(.in(far_1_1474_1[0]), .out(far_1_1474_2[0]));    relay_conn far_1_1474_2_b(.in(far_1_1474_1[1]), .out(far_1_1474_2[1]));
    assign layer_1[454] = far_1_1474_2[0]; 
    wire [1:0] far_1_1475_0;    relay_conn far_1_1475_0_a(.in(layer_0[936]), .out(far_1_1475_0[0]));    relay_conn far_1_1475_0_b(.in(layer_0[880]), .out(far_1_1475_0[1]));
    assign layer_1[455] = far_1_1475_0[0]; 
    wire [1:0] far_1_1476_0;    relay_conn far_1_1476_0_a(.in(layer_0[621]), .out(far_1_1476_0[0]));    relay_conn far_1_1476_0_b(.in(layer_0[497]), .out(far_1_1476_0[1]));
    wire [1:0] far_1_1476_1;    relay_conn far_1_1476_1_a(.in(far_1_1476_0[0]), .out(far_1_1476_1[0]));    relay_conn far_1_1476_1_b(.in(far_1_1476_0[1]), .out(far_1_1476_1[1]));
    wire [1:0] far_1_1476_2;    relay_conn far_1_1476_2_a(.in(far_1_1476_1[0]), .out(far_1_1476_2[0]));    relay_conn far_1_1476_2_b(.in(far_1_1476_1[1]), .out(far_1_1476_2[1]));
    assign layer_1[456] = far_1_1476_2[0] ^ far_1_1476_2[1]; 
    assign layer_1[457] = ~layer_0[839] | (layer_0[839] & layer_0[823]); 
    wire [1:0] far_1_1478_0;    relay_conn far_1_1478_0_a(.in(layer_0[91]), .out(far_1_1478_0[0]));    relay_conn far_1_1478_0_b(.in(layer_0[45]), .out(far_1_1478_0[1]));
    assign layer_1[458] = ~far_1_1478_0[0] | (far_1_1478_0[0] & far_1_1478_0[1]); 
    wire [1:0] far_1_1479_0;    relay_conn far_1_1479_0_a(.in(layer_0[85]), .out(far_1_1479_0[0]));    relay_conn far_1_1479_0_b(.in(layer_0[15]), .out(far_1_1479_0[1]));
    wire [1:0] far_1_1479_1;    relay_conn far_1_1479_1_a(.in(far_1_1479_0[0]), .out(far_1_1479_1[0]));    relay_conn far_1_1479_1_b(.in(far_1_1479_0[1]), .out(far_1_1479_1[1]));
    assign layer_1[459] = ~far_1_1479_1[1] | (far_1_1479_1[0] & far_1_1479_1[1]); 
    wire [1:0] far_1_1480_0;    relay_conn far_1_1480_0_a(.in(layer_0[216]), .out(far_1_1480_0[0]));    relay_conn far_1_1480_0_b(.in(layer_0[321]), .out(far_1_1480_0[1]));
    wire [1:0] far_1_1480_1;    relay_conn far_1_1480_1_a(.in(far_1_1480_0[0]), .out(far_1_1480_1[0]));    relay_conn far_1_1480_1_b(.in(far_1_1480_0[1]), .out(far_1_1480_1[1]));
    wire [1:0] far_1_1480_2;    relay_conn far_1_1480_2_a(.in(far_1_1480_1[0]), .out(far_1_1480_2[0]));    relay_conn far_1_1480_2_b(.in(far_1_1480_1[1]), .out(far_1_1480_2[1]));
    assign layer_1[460] = far_1_1480_2[0] & ~far_1_1480_2[1]; 
    assign layer_1[461] = layer_0[339] & layer_0[308]; 
    wire [1:0] far_1_1482_0;    relay_conn far_1_1482_0_a(.in(layer_0[897]), .out(far_1_1482_0[0]));    relay_conn far_1_1482_0_b(.in(layer_0[855]), .out(far_1_1482_0[1]));
    assign layer_1[462] = far_1_1482_0[1] & ~far_1_1482_0[0]; 
    wire [1:0] far_1_1483_0;    relay_conn far_1_1483_0_a(.in(layer_0[834]), .out(far_1_1483_0[0]));    relay_conn far_1_1483_0_b(.in(layer_0[954]), .out(far_1_1483_0[1]));
    wire [1:0] far_1_1483_1;    relay_conn far_1_1483_1_a(.in(far_1_1483_0[0]), .out(far_1_1483_1[0]));    relay_conn far_1_1483_1_b(.in(far_1_1483_0[1]), .out(far_1_1483_1[1]));
    wire [1:0] far_1_1483_2;    relay_conn far_1_1483_2_a(.in(far_1_1483_1[0]), .out(far_1_1483_2[0]));    relay_conn far_1_1483_2_b(.in(far_1_1483_1[1]), .out(far_1_1483_2[1]));
    assign layer_1[463] = far_1_1483_2[0] | far_1_1483_2[1]; 
    wire [1:0] far_1_1484_0;    relay_conn far_1_1484_0_a(.in(layer_0[1019]), .out(far_1_1484_0[0]));    relay_conn far_1_1484_0_b(.in(layer_0[897]), .out(far_1_1484_0[1]));
    wire [1:0] far_1_1484_1;    relay_conn far_1_1484_1_a(.in(far_1_1484_0[0]), .out(far_1_1484_1[0]));    relay_conn far_1_1484_1_b(.in(far_1_1484_0[1]), .out(far_1_1484_1[1]));
    wire [1:0] far_1_1484_2;    relay_conn far_1_1484_2_a(.in(far_1_1484_1[0]), .out(far_1_1484_2[0]));    relay_conn far_1_1484_2_b(.in(far_1_1484_1[1]), .out(far_1_1484_2[1]));
    assign layer_1[464] = ~far_1_1484_2[1] | (far_1_1484_2[0] & far_1_1484_2[1]); 
    wire [1:0] far_1_1485_0;    relay_conn far_1_1485_0_a(.in(layer_0[187]), .out(far_1_1485_0[0]));    relay_conn far_1_1485_0_b(.in(layer_0[315]), .out(far_1_1485_0[1]));
    wire [1:0] far_1_1485_1;    relay_conn far_1_1485_1_a(.in(far_1_1485_0[0]), .out(far_1_1485_1[0]));    relay_conn far_1_1485_1_b(.in(far_1_1485_0[1]), .out(far_1_1485_1[1]));
    wire [1:0] far_1_1485_2;    relay_conn far_1_1485_2_a(.in(far_1_1485_1[0]), .out(far_1_1485_2[0]));    relay_conn far_1_1485_2_b(.in(far_1_1485_1[1]), .out(far_1_1485_2[1]));
    wire [1:0] far_1_1485_3;    relay_conn far_1_1485_3_a(.in(far_1_1485_2[0]), .out(far_1_1485_3[0]));    relay_conn far_1_1485_3_b(.in(far_1_1485_2[1]), .out(far_1_1485_3[1]));
    assign layer_1[465] = far_1_1485_3[0] & ~far_1_1485_3[1]; 
    wire [1:0] far_1_1486_0;    relay_conn far_1_1486_0_a(.in(layer_0[921]), .out(far_1_1486_0[0]));    relay_conn far_1_1486_0_b(.in(layer_0[858]), .out(far_1_1486_0[1]));
    assign layer_1[466] = ~far_1_1486_0[1]; 
    assign layer_1[467] = layer_0[81]; 
    wire [1:0] far_1_1488_0;    relay_conn far_1_1488_0_a(.in(layer_0[67]), .out(far_1_1488_0[0]));    relay_conn far_1_1488_0_b(.in(layer_0[161]), .out(far_1_1488_0[1]));
    wire [1:0] far_1_1488_1;    relay_conn far_1_1488_1_a(.in(far_1_1488_0[0]), .out(far_1_1488_1[0]));    relay_conn far_1_1488_1_b(.in(far_1_1488_0[1]), .out(far_1_1488_1[1]));
    assign layer_1[468] = far_1_1488_1[0] & far_1_1488_1[1]; 
    wire [1:0] far_1_1489_0;    relay_conn far_1_1489_0_a(.in(layer_0[65]), .out(far_1_1489_0[0]));    relay_conn far_1_1489_0_b(.in(layer_0[114]), .out(far_1_1489_0[1]));
    assign layer_1[469] = far_1_1489_0[0] & far_1_1489_0[1]; 
    wire [1:0] far_1_1490_0;    relay_conn far_1_1490_0_a(.in(layer_0[852]), .out(far_1_1490_0[0]));    relay_conn far_1_1490_0_b(.in(layer_0[899]), .out(far_1_1490_0[1]));
    assign layer_1[470] = far_1_1490_0[0] | far_1_1490_0[1]; 
    wire [1:0] far_1_1491_0;    relay_conn far_1_1491_0_a(.in(layer_0[246]), .out(far_1_1491_0[0]));    relay_conn far_1_1491_0_b(.in(layer_0[131]), .out(far_1_1491_0[1]));
    wire [1:0] far_1_1491_1;    relay_conn far_1_1491_1_a(.in(far_1_1491_0[0]), .out(far_1_1491_1[0]));    relay_conn far_1_1491_1_b(.in(far_1_1491_0[1]), .out(far_1_1491_1[1]));
    wire [1:0] far_1_1491_2;    relay_conn far_1_1491_2_a(.in(far_1_1491_1[0]), .out(far_1_1491_2[0]));    relay_conn far_1_1491_2_b(.in(far_1_1491_1[1]), .out(far_1_1491_2[1]));
    assign layer_1[471] = far_1_1491_2[1]; 
    assign layer_1[472] = ~layer_0[580]; 
    wire [1:0] far_1_1493_0;    relay_conn far_1_1493_0_a(.in(layer_0[964]), .out(far_1_1493_0[0]));    relay_conn far_1_1493_0_b(.in(layer_0[927]), .out(far_1_1493_0[1]));
    assign layer_1[473] = ~(far_1_1493_0[0] | far_1_1493_0[1]); 
    wire [1:0] far_1_1494_0;    relay_conn far_1_1494_0_a(.in(layer_0[57]), .out(far_1_1494_0[0]));    relay_conn far_1_1494_0_b(.in(layer_0[116]), .out(far_1_1494_0[1]));
    assign layer_1[474] = ~far_1_1494_0[0] | (far_1_1494_0[0] & far_1_1494_0[1]); 
    wire [1:0] far_1_1495_0;    relay_conn far_1_1495_0_a(.in(layer_0[347]), .out(far_1_1495_0[0]));    relay_conn far_1_1495_0_b(.in(layer_0[301]), .out(far_1_1495_0[1]));
    assign layer_1[475] = far_1_1495_0[0] & ~far_1_1495_0[1]; 
    assign layer_1[476] = ~(layer_0[356] & layer_0[367]); 
    assign layer_1[477] = ~(layer_0[246] | layer_0[242]); 
    wire [1:0] far_1_1498_0;    relay_conn far_1_1498_0_a(.in(layer_0[400]), .out(far_1_1498_0[0]));    relay_conn far_1_1498_0_b(.in(layer_0[284]), .out(far_1_1498_0[1]));
    wire [1:0] far_1_1498_1;    relay_conn far_1_1498_1_a(.in(far_1_1498_0[0]), .out(far_1_1498_1[0]));    relay_conn far_1_1498_1_b(.in(far_1_1498_0[1]), .out(far_1_1498_1[1]));
    wire [1:0] far_1_1498_2;    relay_conn far_1_1498_2_a(.in(far_1_1498_1[0]), .out(far_1_1498_2[0]));    relay_conn far_1_1498_2_b(.in(far_1_1498_1[1]), .out(far_1_1498_2[1]));
    assign layer_1[478] = far_1_1498_2[0]; 
    wire [1:0] far_1_1499_0;    relay_conn far_1_1499_0_a(.in(layer_0[251]), .out(far_1_1499_0[0]));    relay_conn far_1_1499_0_b(.in(layer_0[336]), .out(far_1_1499_0[1]));
    wire [1:0] far_1_1499_1;    relay_conn far_1_1499_1_a(.in(far_1_1499_0[0]), .out(far_1_1499_1[0]));    relay_conn far_1_1499_1_b(.in(far_1_1499_0[1]), .out(far_1_1499_1[1]));
    assign layer_1[479] = far_1_1499_1[0] & ~far_1_1499_1[1]; 
    wire [1:0] far_1_1500_0;    relay_conn far_1_1500_0_a(.in(layer_0[579]), .out(far_1_1500_0[0]));    relay_conn far_1_1500_0_b(.in(layer_0[505]), .out(far_1_1500_0[1]));
    wire [1:0] far_1_1500_1;    relay_conn far_1_1500_1_a(.in(far_1_1500_0[0]), .out(far_1_1500_1[0]));    relay_conn far_1_1500_1_b(.in(far_1_1500_0[1]), .out(far_1_1500_1[1]));
    assign layer_1[480] = ~far_1_1500_1[1] | (far_1_1500_1[0] & far_1_1500_1[1]); 
    wire [1:0] far_1_1501_0;    relay_conn far_1_1501_0_a(.in(layer_0[122]), .out(far_1_1501_0[0]));    relay_conn far_1_1501_0_b(.in(layer_0[65]), .out(far_1_1501_0[1]));
    assign layer_1[481] = far_1_1501_0[0] & far_1_1501_0[1]; 
    wire [1:0] far_1_1502_0;    relay_conn far_1_1502_0_a(.in(layer_0[478]), .out(far_1_1502_0[0]));    relay_conn far_1_1502_0_b(.in(layer_0[572]), .out(far_1_1502_0[1]));
    wire [1:0] far_1_1502_1;    relay_conn far_1_1502_1_a(.in(far_1_1502_0[0]), .out(far_1_1502_1[0]));    relay_conn far_1_1502_1_b(.in(far_1_1502_0[1]), .out(far_1_1502_1[1]));
    assign layer_1[482] = far_1_1502_1[0] & ~far_1_1502_1[1]; 
    assign layer_1[483] = ~(layer_0[400] | layer_0[403]); 
    wire [1:0] far_1_1504_0;    relay_conn far_1_1504_0_a(.in(layer_0[997]), .out(far_1_1504_0[0]));    relay_conn far_1_1504_0_b(.in(layer_0[915]), .out(far_1_1504_0[1]));
    wire [1:0] far_1_1504_1;    relay_conn far_1_1504_1_a(.in(far_1_1504_0[0]), .out(far_1_1504_1[0]));    relay_conn far_1_1504_1_b(.in(far_1_1504_0[1]), .out(far_1_1504_1[1]));
    assign layer_1[484] = ~(far_1_1504_1[0] | far_1_1504_1[1]); 
    wire [1:0] far_1_1505_0;    relay_conn far_1_1505_0_a(.in(layer_0[441]), .out(far_1_1505_0[0]));    relay_conn far_1_1505_0_b(.in(layer_0[482]), .out(far_1_1505_0[1]));
    assign layer_1[485] = far_1_1505_0[1] & ~far_1_1505_0[0]; 
    wire [1:0] far_1_1506_0;    relay_conn far_1_1506_0_a(.in(layer_0[85]), .out(far_1_1506_0[0]));    relay_conn far_1_1506_0_b(.in(layer_0[8]), .out(far_1_1506_0[1]));
    wire [1:0] far_1_1506_1;    relay_conn far_1_1506_1_a(.in(far_1_1506_0[0]), .out(far_1_1506_1[0]));    relay_conn far_1_1506_1_b(.in(far_1_1506_0[1]), .out(far_1_1506_1[1]));
    assign layer_1[486] = far_1_1506_1[0] ^ far_1_1506_1[1]; 
    wire [1:0] far_1_1507_0;    relay_conn far_1_1507_0_a(.in(layer_0[915]), .out(far_1_1507_0[0]));    relay_conn far_1_1507_0_b(.in(layer_0[829]), .out(far_1_1507_0[1]));
    wire [1:0] far_1_1507_1;    relay_conn far_1_1507_1_a(.in(far_1_1507_0[0]), .out(far_1_1507_1[0]));    relay_conn far_1_1507_1_b(.in(far_1_1507_0[1]), .out(far_1_1507_1[1]));
    assign layer_1[487] = ~(far_1_1507_1[0] ^ far_1_1507_1[1]); 
    assign layer_1[488] = layer_0[187]; 
    wire [1:0] far_1_1509_0;    relay_conn far_1_1509_0_a(.in(layer_0[444]), .out(far_1_1509_0[0]));    relay_conn far_1_1509_0_b(.in(layer_0[396]), .out(far_1_1509_0[1]));
    assign layer_1[489] = ~(far_1_1509_0[0] | far_1_1509_0[1]); 
    assign layer_1[490] = layer_0[658] & ~layer_0[638]; 
    assign layer_1[491] = ~(layer_0[827] | layer_0[847]); 
    wire [1:0] far_1_1512_0;    relay_conn far_1_1512_0_a(.in(layer_0[314]), .out(far_1_1512_0[0]));    relay_conn far_1_1512_0_b(.in(layer_0[395]), .out(far_1_1512_0[1]));
    wire [1:0] far_1_1512_1;    relay_conn far_1_1512_1_a(.in(far_1_1512_0[0]), .out(far_1_1512_1[0]));    relay_conn far_1_1512_1_b(.in(far_1_1512_0[1]), .out(far_1_1512_1[1]));
    assign layer_1[492] = far_1_1512_1[0] & ~far_1_1512_1[1]; 
    wire [1:0] far_1_1513_0;    relay_conn far_1_1513_0_a(.in(layer_0[484]), .out(far_1_1513_0[0]));    relay_conn far_1_1513_0_b(.in(layer_0[412]), .out(far_1_1513_0[1]));
    wire [1:0] far_1_1513_1;    relay_conn far_1_1513_1_a(.in(far_1_1513_0[0]), .out(far_1_1513_1[0]));    relay_conn far_1_1513_1_b(.in(far_1_1513_0[1]), .out(far_1_1513_1[1]));
    assign layer_1[493] = ~(far_1_1513_1[0] & far_1_1513_1[1]); 
    wire [1:0] far_1_1514_0;    relay_conn far_1_1514_0_a(.in(layer_0[676]), .out(far_1_1514_0[0]));    relay_conn far_1_1514_0_b(.in(layer_0[583]), .out(far_1_1514_0[1]));
    wire [1:0] far_1_1514_1;    relay_conn far_1_1514_1_a(.in(far_1_1514_0[0]), .out(far_1_1514_1[0]));    relay_conn far_1_1514_1_b(.in(far_1_1514_0[1]), .out(far_1_1514_1[1]));
    assign layer_1[494] = far_1_1514_1[0] & far_1_1514_1[1]; 
    wire [1:0] far_1_1515_0;    relay_conn far_1_1515_0_a(.in(layer_0[187]), .out(far_1_1515_0[0]));    relay_conn far_1_1515_0_b(.in(layer_0[267]), .out(far_1_1515_0[1]));
    wire [1:0] far_1_1515_1;    relay_conn far_1_1515_1_a(.in(far_1_1515_0[0]), .out(far_1_1515_1[0]));    relay_conn far_1_1515_1_b(.in(far_1_1515_0[1]), .out(far_1_1515_1[1]));
    assign layer_1[495] = far_1_1515_1[0] ^ far_1_1515_1[1]; 
    wire [1:0] far_1_1516_0;    relay_conn far_1_1516_0_a(.in(layer_0[523]), .out(far_1_1516_0[0]));    relay_conn far_1_1516_0_b(.in(layer_0[420]), .out(far_1_1516_0[1]));
    wire [1:0] far_1_1516_1;    relay_conn far_1_1516_1_a(.in(far_1_1516_0[0]), .out(far_1_1516_1[0]));    relay_conn far_1_1516_1_b(.in(far_1_1516_0[1]), .out(far_1_1516_1[1]));
    wire [1:0] far_1_1516_2;    relay_conn far_1_1516_2_a(.in(far_1_1516_1[0]), .out(far_1_1516_2[0]));    relay_conn far_1_1516_2_b(.in(far_1_1516_1[1]), .out(far_1_1516_2[1]));
    assign layer_1[496] = ~far_1_1516_2[0] | (far_1_1516_2[0] & far_1_1516_2[1]); 
    assign layer_1[497] = ~(layer_0[395] & layer_0[419]); 
    wire [1:0] far_1_1518_0;    relay_conn far_1_1518_0_a(.in(layer_0[471]), .out(far_1_1518_0[0]));    relay_conn far_1_1518_0_b(.in(layer_0[354]), .out(far_1_1518_0[1]));
    wire [1:0] far_1_1518_1;    relay_conn far_1_1518_1_a(.in(far_1_1518_0[0]), .out(far_1_1518_1[0]));    relay_conn far_1_1518_1_b(.in(far_1_1518_0[1]), .out(far_1_1518_1[1]));
    wire [1:0] far_1_1518_2;    relay_conn far_1_1518_2_a(.in(far_1_1518_1[0]), .out(far_1_1518_2[0]));    relay_conn far_1_1518_2_b(.in(far_1_1518_1[1]), .out(far_1_1518_2[1]));
    assign layer_1[498] = ~far_1_1518_2[1]; 
    assign layer_1[499] = layer_0[74] | layer_0[94]; 
    wire [1:0] far_1_1520_0;    relay_conn far_1_1520_0_a(.in(layer_0[438]), .out(far_1_1520_0[0]));    relay_conn far_1_1520_0_b(.in(layer_0[543]), .out(far_1_1520_0[1]));
    wire [1:0] far_1_1520_1;    relay_conn far_1_1520_1_a(.in(far_1_1520_0[0]), .out(far_1_1520_1[0]));    relay_conn far_1_1520_1_b(.in(far_1_1520_0[1]), .out(far_1_1520_1[1]));
    wire [1:0] far_1_1520_2;    relay_conn far_1_1520_2_a(.in(far_1_1520_1[0]), .out(far_1_1520_2[0]));    relay_conn far_1_1520_2_b(.in(far_1_1520_1[1]), .out(far_1_1520_2[1]));
    assign layer_1[500] = ~far_1_1520_2[0]; 
    wire [1:0] far_1_1521_0;    relay_conn far_1_1521_0_a(.in(layer_0[681]), .out(far_1_1521_0[0]));    relay_conn far_1_1521_0_b(.in(layer_0[777]), .out(far_1_1521_0[1]));
    wire [1:0] far_1_1521_1;    relay_conn far_1_1521_1_a(.in(far_1_1521_0[0]), .out(far_1_1521_1[0]));    relay_conn far_1_1521_1_b(.in(far_1_1521_0[1]), .out(far_1_1521_1[1]));
    wire [1:0] far_1_1521_2;    relay_conn far_1_1521_2_a(.in(far_1_1521_1[0]), .out(far_1_1521_2[0]));    relay_conn far_1_1521_2_b(.in(far_1_1521_1[1]), .out(far_1_1521_2[1]));
    assign layer_1[501] = far_1_1521_2[0] & ~far_1_1521_2[1]; 
    assign layer_1[502] = ~(layer_0[512] & layer_0[508]); 
    wire [1:0] far_1_1523_0;    relay_conn far_1_1523_0_a(.in(layer_0[277]), .out(far_1_1523_0[0]));    relay_conn far_1_1523_0_b(.in(layer_0[150]), .out(far_1_1523_0[1]));
    wire [1:0] far_1_1523_1;    relay_conn far_1_1523_1_a(.in(far_1_1523_0[0]), .out(far_1_1523_1[0]));    relay_conn far_1_1523_1_b(.in(far_1_1523_0[1]), .out(far_1_1523_1[1]));
    wire [1:0] far_1_1523_2;    relay_conn far_1_1523_2_a(.in(far_1_1523_1[0]), .out(far_1_1523_2[0]));    relay_conn far_1_1523_2_b(.in(far_1_1523_1[1]), .out(far_1_1523_2[1]));
    assign layer_1[503] = ~(far_1_1523_2[0] & far_1_1523_2[1]); 
    wire [1:0] far_1_1524_0;    relay_conn far_1_1524_0_a(.in(layer_0[964]), .out(far_1_1524_0[0]));    relay_conn far_1_1524_0_b(.in(layer_0[859]), .out(far_1_1524_0[1]));
    wire [1:0] far_1_1524_1;    relay_conn far_1_1524_1_a(.in(far_1_1524_0[0]), .out(far_1_1524_1[0]));    relay_conn far_1_1524_1_b(.in(far_1_1524_0[1]), .out(far_1_1524_1[1]));
    wire [1:0] far_1_1524_2;    relay_conn far_1_1524_2_a(.in(far_1_1524_1[0]), .out(far_1_1524_2[0]));    relay_conn far_1_1524_2_b(.in(far_1_1524_1[1]), .out(far_1_1524_2[1]));
    assign layer_1[504] = ~far_1_1524_2[1]; 
    wire [1:0] far_1_1525_0;    relay_conn far_1_1525_0_a(.in(layer_0[381]), .out(far_1_1525_0[0]));    relay_conn far_1_1525_0_b(.in(layer_0[431]), .out(far_1_1525_0[1]));
    assign layer_1[505] = ~(far_1_1525_0[0] | far_1_1525_0[1]); 
    assign layer_1[506] = layer_0[444] & ~layer_0[467]; 
    assign layer_1[507] = layer_0[123] & layer_0[95]; 
    assign layer_1[508] = ~(layer_0[413] & layer_0[391]); 
    wire [1:0] far_1_1529_0;    relay_conn far_1_1529_0_a(.in(layer_0[535]), .out(far_1_1529_0[0]));    relay_conn far_1_1529_0_b(.in(layer_0[412]), .out(far_1_1529_0[1]));
    wire [1:0] far_1_1529_1;    relay_conn far_1_1529_1_a(.in(far_1_1529_0[0]), .out(far_1_1529_1[0]));    relay_conn far_1_1529_1_b(.in(far_1_1529_0[1]), .out(far_1_1529_1[1]));
    wire [1:0] far_1_1529_2;    relay_conn far_1_1529_2_a(.in(far_1_1529_1[0]), .out(far_1_1529_2[0]));    relay_conn far_1_1529_2_b(.in(far_1_1529_1[1]), .out(far_1_1529_2[1]));
    assign layer_1[509] = far_1_1529_2[1] & ~far_1_1529_2[0]; 
    wire [1:0] far_1_1530_0;    relay_conn far_1_1530_0_a(.in(layer_0[379]), .out(far_1_1530_0[0]));    relay_conn far_1_1530_0_b(.in(layer_0[254]), .out(far_1_1530_0[1]));
    wire [1:0] far_1_1530_1;    relay_conn far_1_1530_1_a(.in(far_1_1530_0[0]), .out(far_1_1530_1[0]));    relay_conn far_1_1530_1_b(.in(far_1_1530_0[1]), .out(far_1_1530_1[1]));
    wire [1:0] far_1_1530_2;    relay_conn far_1_1530_2_a(.in(far_1_1530_1[0]), .out(far_1_1530_2[0]));    relay_conn far_1_1530_2_b(.in(far_1_1530_1[1]), .out(far_1_1530_2[1]));
    assign layer_1[510] = ~(far_1_1530_2[0] & far_1_1530_2[1]); 
    wire [1:0] far_1_1531_0;    relay_conn far_1_1531_0_a(.in(layer_0[305]), .out(far_1_1531_0[0]));    relay_conn far_1_1531_0_b(.in(layer_0[224]), .out(far_1_1531_0[1]));
    wire [1:0] far_1_1531_1;    relay_conn far_1_1531_1_a(.in(far_1_1531_0[0]), .out(far_1_1531_1[0]));    relay_conn far_1_1531_1_b(.in(far_1_1531_0[1]), .out(far_1_1531_1[1]));
    assign layer_1[511] = far_1_1531_1[1] & ~far_1_1531_1[0]; 
    wire [1:0] far_1_1532_0;    relay_conn far_1_1532_0_a(.in(layer_0[1]), .out(far_1_1532_0[0]));    relay_conn far_1_1532_0_b(.in(layer_0[94]), .out(far_1_1532_0[1]));
    wire [1:0] far_1_1532_1;    relay_conn far_1_1532_1_a(.in(far_1_1532_0[0]), .out(far_1_1532_1[0]));    relay_conn far_1_1532_1_b(.in(far_1_1532_0[1]), .out(far_1_1532_1[1]));
    assign layer_1[512] = far_1_1532_1[1]; 
    wire [1:0] far_1_1533_0;    relay_conn far_1_1533_0_a(.in(layer_0[378]), .out(far_1_1533_0[0]));    relay_conn far_1_1533_0_b(.in(layer_0[253]), .out(far_1_1533_0[1]));
    wire [1:0] far_1_1533_1;    relay_conn far_1_1533_1_a(.in(far_1_1533_0[0]), .out(far_1_1533_1[0]));    relay_conn far_1_1533_1_b(.in(far_1_1533_0[1]), .out(far_1_1533_1[1]));
    wire [1:0] far_1_1533_2;    relay_conn far_1_1533_2_a(.in(far_1_1533_1[0]), .out(far_1_1533_2[0]));    relay_conn far_1_1533_2_b(.in(far_1_1533_1[1]), .out(far_1_1533_2[1]));
    assign layer_1[513] = ~(far_1_1533_2[0] | far_1_1533_2[1]); 
    wire [1:0] far_1_1534_0;    relay_conn far_1_1534_0_a(.in(layer_0[828]), .out(far_1_1534_0[0]));    relay_conn far_1_1534_0_b(.in(layer_0[896]), .out(far_1_1534_0[1]));
    wire [1:0] far_1_1534_1;    relay_conn far_1_1534_1_a(.in(far_1_1534_0[0]), .out(far_1_1534_1[0]));    relay_conn far_1_1534_1_b(.in(far_1_1534_0[1]), .out(far_1_1534_1[1]));
    assign layer_1[514] = ~far_1_1534_1[0]; 
    assign layer_1[515] = ~(layer_0[304] ^ layer_0[309]); 
    wire [1:0] far_1_1536_0;    relay_conn far_1_1536_0_a(.in(layer_0[438]), .out(far_1_1536_0[0]));    relay_conn far_1_1536_0_b(.in(layer_0[330]), .out(far_1_1536_0[1]));
    wire [1:0] far_1_1536_1;    relay_conn far_1_1536_1_a(.in(far_1_1536_0[0]), .out(far_1_1536_1[0]));    relay_conn far_1_1536_1_b(.in(far_1_1536_0[1]), .out(far_1_1536_1[1]));
    wire [1:0] far_1_1536_2;    relay_conn far_1_1536_2_a(.in(far_1_1536_1[0]), .out(far_1_1536_2[0]));    relay_conn far_1_1536_2_b(.in(far_1_1536_1[1]), .out(far_1_1536_2[1]));
    assign layer_1[516] = far_1_1536_2[0] & far_1_1536_2[1]; 
    wire [1:0] far_1_1537_0;    relay_conn far_1_1537_0_a(.in(layer_0[627]), .out(far_1_1537_0[0]));    relay_conn far_1_1537_0_b(.in(layer_0[501]), .out(far_1_1537_0[1]));
    wire [1:0] far_1_1537_1;    relay_conn far_1_1537_1_a(.in(far_1_1537_0[0]), .out(far_1_1537_1[0]));    relay_conn far_1_1537_1_b(.in(far_1_1537_0[1]), .out(far_1_1537_1[1]));
    wire [1:0] far_1_1537_2;    relay_conn far_1_1537_2_a(.in(far_1_1537_1[0]), .out(far_1_1537_2[0]));    relay_conn far_1_1537_2_b(.in(far_1_1537_1[1]), .out(far_1_1537_2[1]));
    assign layer_1[517] = ~far_1_1537_2[1]; 
    wire [1:0] far_1_1538_0;    relay_conn far_1_1538_0_a(.in(layer_0[513]), .out(far_1_1538_0[0]));    relay_conn far_1_1538_0_b(.in(layer_0[555]), .out(far_1_1538_0[1]));
    assign layer_1[518] = far_1_1538_0[0] & ~far_1_1538_0[1]; 
    wire [1:0] far_1_1539_0;    relay_conn far_1_1539_0_a(.in(layer_0[762]), .out(far_1_1539_0[0]));    relay_conn far_1_1539_0_b(.in(layer_0[870]), .out(far_1_1539_0[1]));
    wire [1:0] far_1_1539_1;    relay_conn far_1_1539_1_a(.in(far_1_1539_0[0]), .out(far_1_1539_1[0]));    relay_conn far_1_1539_1_b(.in(far_1_1539_0[1]), .out(far_1_1539_1[1]));
    wire [1:0] far_1_1539_2;    relay_conn far_1_1539_2_a(.in(far_1_1539_1[0]), .out(far_1_1539_2[0]));    relay_conn far_1_1539_2_b(.in(far_1_1539_1[1]), .out(far_1_1539_2[1]));
    assign layer_1[519] = far_1_1539_2[0]; 
    wire [1:0] far_1_1540_0;    relay_conn far_1_1540_0_a(.in(layer_0[272]), .out(far_1_1540_0[0]));    relay_conn far_1_1540_0_b(.in(layer_0[392]), .out(far_1_1540_0[1]));
    wire [1:0] far_1_1540_1;    relay_conn far_1_1540_1_a(.in(far_1_1540_0[0]), .out(far_1_1540_1[0]));    relay_conn far_1_1540_1_b(.in(far_1_1540_0[1]), .out(far_1_1540_1[1]));
    wire [1:0] far_1_1540_2;    relay_conn far_1_1540_2_a(.in(far_1_1540_1[0]), .out(far_1_1540_2[0]));    relay_conn far_1_1540_2_b(.in(far_1_1540_1[1]), .out(far_1_1540_2[1]));
    assign layer_1[520] = far_1_1540_2[0] & far_1_1540_2[1]; 
    assign layer_1[521] = ~layer_0[841] | (layer_0[860] & layer_0[841]); 
    assign layer_1[522] = layer_0[16] & ~layer_0[42]; 
    wire [1:0] far_1_1543_0;    relay_conn far_1_1543_0_a(.in(layer_0[358]), .out(far_1_1543_0[0]));    relay_conn far_1_1543_0_b(.in(layer_0[253]), .out(far_1_1543_0[1]));
    wire [1:0] far_1_1543_1;    relay_conn far_1_1543_1_a(.in(far_1_1543_0[0]), .out(far_1_1543_1[0]));    relay_conn far_1_1543_1_b(.in(far_1_1543_0[1]), .out(far_1_1543_1[1]));
    wire [1:0] far_1_1543_2;    relay_conn far_1_1543_2_a(.in(far_1_1543_1[0]), .out(far_1_1543_2[0]));    relay_conn far_1_1543_2_b(.in(far_1_1543_1[1]), .out(far_1_1543_2[1]));
    assign layer_1[523] = ~far_1_1543_2[0] | (far_1_1543_2[0] & far_1_1543_2[1]); 
    wire [1:0] far_1_1544_0;    relay_conn far_1_1544_0_a(.in(layer_0[798]), .out(far_1_1544_0[0]));    relay_conn far_1_1544_0_b(.in(layer_0[838]), .out(far_1_1544_0[1]));
    assign layer_1[524] = far_1_1544_0[0] | far_1_1544_0[1]; 
    assign layer_1[525] = ~layer_0[879] | (layer_0[879] & layer_0[853]); 
    wire [1:0] far_1_1546_0;    relay_conn far_1_1546_0_a(.in(layer_0[384]), .out(far_1_1546_0[0]));    relay_conn far_1_1546_0_b(.in(layer_0[476]), .out(far_1_1546_0[1]));
    wire [1:0] far_1_1546_1;    relay_conn far_1_1546_1_a(.in(far_1_1546_0[0]), .out(far_1_1546_1[0]));    relay_conn far_1_1546_1_b(.in(far_1_1546_0[1]), .out(far_1_1546_1[1]));
    assign layer_1[526] = ~far_1_1546_1[0] | (far_1_1546_1[0] & far_1_1546_1[1]); 
    wire [1:0] far_1_1547_0;    relay_conn far_1_1547_0_a(.in(layer_0[200]), .out(far_1_1547_0[0]));    relay_conn far_1_1547_0_b(.in(layer_0[115]), .out(far_1_1547_0[1]));
    wire [1:0] far_1_1547_1;    relay_conn far_1_1547_1_a(.in(far_1_1547_0[0]), .out(far_1_1547_1[0]));    relay_conn far_1_1547_1_b(.in(far_1_1547_0[1]), .out(far_1_1547_1[1]));
    assign layer_1[527] = ~far_1_1547_1[1]; 
    wire [1:0] far_1_1548_0;    relay_conn far_1_1548_0_a(.in(layer_0[834]), .out(far_1_1548_0[0]));    relay_conn far_1_1548_0_b(.in(layer_0[750]), .out(far_1_1548_0[1]));
    wire [1:0] far_1_1548_1;    relay_conn far_1_1548_1_a(.in(far_1_1548_0[0]), .out(far_1_1548_1[0]));    relay_conn far_1_1548_1_b(.in(far_1_1548_0[1]), .out(far_1_1548_1[1]));
    assign layer_1[528] = ~(far_1_1548_1[0] ^ far_1_1548_1[1]); 
    assign layer_1[529] = layer_0[847] & layer_0[826]; 
    wire [1:0] far_1_1550_0;    relay_conn far_1_1550_0_a(.in(layer_0[906]), .out(far_1_1550_0[0]));    relay_conn far_1_1550_0_b(.in(layer_0[866]), .out(far_1_1550_0[1]));
    assign layer_1[530] = ~far_1_1550_0[1]; 
    wire [1:0] far_1_1551_0;    relay_conn far_1_1551_0_a(.in(layer_0[187]), .out(far_1_1551_0[0]));    relay_conn far_1_1551_0_b(.in(layer_0[70]), .out(far_1_1551_0[1]));
    wire [1:0] far_1_1551_1;    relay_conn far_1_1551_1_a(.in(far_1_1551_0[0]), .out(far_1_1551_1[0]));    relay_conn far_1_1551_1_b(.in(far_1_1551_0[1]), .out(far_1_1551_1[1]));
    wire [1:0] far_1_1551_2;    relay_conn far_1_1551_2_a(.in(far_1_1551_1[0]), .out(far_1_1551_2[0]));    relay_conn far_1_1551_2_b(.in(far_1_1551_1[1]), .out(far_1_1551_2[1]));
    assign layer_1[531] = far_1_1551_2[0] | far_1_1551_2[1]; 
    wire [1:0] far_1_1552_0;    relay_conn far_1_1552_0_a(.in(layer_0[54]), .out(far_1_1552_0[0]));    relay_conn far_1_1552_0_b(.in(layer_0[108]), .out(far_1_1552_0[1]));
    assign layer_1[532] = ~(far_1_1552_0[0] | far_1_1552_0[1]); 
    assign layer_1[533] = layer_0[293] & ~layer_0[291]; 
    assign layer_1[534] = layer_0[858] & layer_0[886]; 
    wire [1:0] far_1_1555_0;    relay_conn far_1_1555_0_a(.in(layer_0[511]), .out(far_1_1555_0[0]));    relay_conn far_1_1555_0_b(.in(layer_0[559]), .out(far_1_1555_0[1]));
    assign layer_1[535] = far_1_1555_0[0] & ~far_1_1555_0[1]; 
    wire [1:0] far_1_1556_0;    relay_conn far_1_1556_0_a(.in(layer_0[331]), .out(far_1_1556_0[0]));    relay_conn far_1_1556_0_b(.in(layer_0[208]), .out(far_1_1556_0[1]));
    wire [1:0] far_1_1556_1;    relay_conn far_1_1556_1_a(.in(far_1_1556_0[0]), .out(far_1_1556_1[0]));    relay_conn far_1_1556_1_b(.in(far_1_1556_0[1]), .out(far_1_1556_1[1]));
    wire [1:0] far_1_1556_2;    relay_conn far_1_1556_2_a(.in(far_1_1556_1[0]), .out(far_1_1556_2[0]));    relay_conn far_1_1556_2_b(.in(far_1_1556_1[1]), .out(far_1_1556_2[1]));
    assign layer_1[536] = ~far_1_1556_2[0]; 
    wire [1:0] far_1_1557_0;    relay_conn far_1_1557_0_a(.in(layer_0[89]), .out(far_1_1557_0[0]));    relay_conn far_1_1557_0_b(.in(layer_0[156]), .out(far_1_1557_0[1]));
    wire [1:0] far_1_1557_1;    relay_conn far_1_1557_1_a(.in(far_1_1557_0[0]), .out(far_1_1557_1[0]));    relay_conn far_1_1557_1_b(.in(far_1_1557_0[1]), .out(far_1_1557_1[1]));
    assign layer_1[537] = ~far_1_1557_1[0] | (far_1_1557_1[0] & far_1_1557_1[1]); 
    assign layer_1[538] = ~layer_0[415]; 
    wire [1:0] far_1_1559_0;    relay_conn far_1_1559_0_a(.in(layer_0[839]), .out(far_1_1559_0[0]));    relay_conn far_1_1559_0_b(.in(layer_0[734]), .out(far_1_1559_0[1]));
    wire [1:0] far_1_1559_1;    relay_conn far_1_1559_1_a(.in(far_1_1559_0[0]), .out(far_1_1559_1[0]));    relay_conn far_1_1559_1_b(.in(far_1_1559_0[1]), .out(far_1_1559_1[1]));
    wire [1:0] far_1_1559_2;    relay_conn far_1_1559_2_a(.in(far_1_1559_1[0]), .out(far_1_1559_2[0]));    relay_conn far_1_1559_2_b(.in(far_1_1559_1[1]), .out(far_1_1559_2[1]));
    assign layer_1[539] = ~(far_1_1559_2[0] | far_1_1559_2[1]); 
    assign layer_1[540] = ~(layer_0[255] ^ layer_0[265]); 
    wire [1:0] far_1_1561_0;    relay_conn far_1_1561_0_a(.in(layer_0[828]), .out(far_1_1561_0[0]));    relay_conn far_1_1561_0_b(.in(layer_0[954]), .out(far_1_1561_0[1]));
    wire [1:0] far_1_1561_1;    relay_conn far_1_1561_1_a(.in(far_1_1561_0[0]), .out(far_1_1561_1[0]));    relay_conn far_1_1561_1_b(.in(far_1_1561_0[1]), .out(far_1_1561_1[1]));
    wire [1:0] far_1_1561_2;    relay_conn far_1_1561_2_a(.in(far_1_1561_1[0]), .out(far_1_1561_2[0]));    relay_conn far_1_1561_2_b(.in(far_1_1561_1[1]), .out(far_1_1561_2[1]));
    assign layer_1[541] = ~far_1_1561_2[0] | (far_1_1561_2[0] & far_1_1561_2[1]); 
    wire [1:0] far_1_1562_0;    relay_conn far_1_1562_0_a(.in(layer_0[996]), .out(far_1_1562_0[0]));    relay_conn far_1_1562_0_b(.in(layer_0[896]), .out(far_1_1562_0[1]));
    wire [1:0] far_1_1562_1;    relay_conn far_1_1562_1_a(.in(far_1_1562_0[0]), .out(far_1_1562_1[0]));    relay_conn far_1_1562_1_b(.in(far_1_1562_0[1]), .out(far_1_1562_1[1]));
    wire [1:0] far_1_1562_2;    relay_conn far_1_1562_2_a(.in(far_1_1562_1[0]), .out(far_1_1562_2[0]));    relay_conn far_1_1562_2_b(.in(far_1_1562_1[1]), .out(far_1_1562_2[1]));
    assign layer_1[542] = ~(far_1_1562_2[0] & far_1_1562_2[1]); 
    wire [1:0] far_1_1563_0;    relay_conn far_1_1563_0_a(.in(layer_0[484]), .out(far_1_1563_0[0]));    relay_conn far_1_1563_0_b(.in(layer_0[380]), .out(far_1_1563_0[1]));
    wire [1:0] far_1_1563_1;    relay_conn far_1_1563_1_a(.in(far_1_1563_0[0]), .out(far_1_1563_1[0]));    relay_conn far_1_1563_1_b(.in(far_1_1563_0[1]), .out(far_1_1563_1[1]));
    wire [1:0] far_1_1563_2;    relay_conn far_1_1563_2_a(.in(far_1_1563_1[0]), .out(far_1_1563_2[0]));    relay_conn far_1_1563_2_b(.in(far_1_1563_1[1]), .out(far_1_1563_2[1]));
    assign layer_1[543] = far_1_1563_2[1] & ~far_1_1563_2[0]; 
    wire [1:0] far_1_1564_0;    relay_conn far_1_1564_0_a(.in(layer_0[626]), .out(far_1_1564_0[0]));    relay_conn far_1_1564_0_b(.in(layer_0[580]), .out(far_1_1564_0[1]));
    assign layer_1[544] = far_1_1564_0[0] | far_1_1564_0[1]; 
    wire [1:0] far_1_1565_0;    relay_conn far_1_1565_0_a(.in(layer_0[861]), .out(far_1_1565_0[0]));    relay_conn far_1_1565_0_b(.in(layer_0[821]), .out(far_1_1565_0[1]));
    assign layer_1[545] = far_1_1565_0[0] & ~far_1_1565_0[1]; 
    wire [1:0] far_1_1566_0;    relay_conn far_1_1566_0_a(.in(layer_0[546]), .out(far_1_1566_0[0]));    relay_conn far_1_1566_0_b(.in(layer_0[446]), .out(far_1_1566_0[1]));
    wire [1:0] far_1_1566_1;    relay_conn far_1_1566_1_a(.in(far_1_1566_0[0]), .out(far_1_1566_1[0]));    relay_conn far_1_1566_1_b(.in(far_1_1566_0[1]), .out(far_1_1566_1[1]));
    wire [1:0] far_1_1566_2;    relay_conn far_1_1566_2_a(.in(far_1_1566_1[0]), .out(far_1_1566_2[0]));    relay_conn far_1_1566_2_b(.in(far_1_1566_1[1]), .out(far_1_1566_2[1]));
    assign layer_1[546] = far_1_1566_2[1] & ~far_1_1566_2[0]; 
    assign layer_1[547] = layer_0[37] & ~layer_0[30]; 
    wire [1:0] far_1_1568_0;    relay_conn far_1_1568_0_a(.in(layer_0[734]), .out(far_1_1568_0[0]));    relay_conn far_1_1568_0_b(.in(layer_0[834]), .out(far_1_1568_0[1]));
    wire [1:0] far_1_1568_1;    relay_conn far_1_1568_1_a(.in(far_1_1568_0[0]), .out(far_1_1568_1[0]));    relay_conn far_1_1568_1_b(.in(far_1_1568_0[1]), .out(far_1_1568_1[1]));
    wire [1:0] far_1_1568_2;    relay_conn far_1_1568_2_a(.in(far_1_1568_1[0]), .out(far_1_1568_2[0]));    relay_conn far_1_1568_2_b(.in(far_1_1568_1[1]), .out(far_1_1568_2[1]));
    assign layer_1[548] = ~far_1_1568_2[0]; 
    assign layer_1[549] = ~(layer_0[27] | layer_0[51]); 
    wire [1:0] far_1_1570_0;    relay_conn far_1_1570_0_a(.in(layer_0[819]), .out(far_1_1570_0[0]));    relay_conn far_1_1570_0_b(.in(layer_0[896]), .out(far_1_1570_0[1]));
    wire [1:0] far_1_1570_1;    relay_conn far_1_1570_1_a(.in(far_1_1570_0[0]), .out(far_1_1570_1[0]));    relay_conn far_1_1570_1_b(.in(far_1_1570_0[1]), .out(far_1_1570_1[1]));
    assign layer_1[550] = far_1_1570_1[1] & ~far_1_1570_1[0]; 
    assign layer_1[551] = ~(layer_0[355] & layer_0[337]); 
    wire [1:0] far_1_1572_0;    relay_conn far_1_1572_0_a(.in(layer_0[908]), .out(far_1_1572_0[0]));    relay_conn far_1_1572_0_b(.in(layer_0[849]), .out(far_1_1572_0[1]));
    assign layer_1[552] = ~(far_1_1572_0[0] | far_1_1572_0[1]); 
    wire [1:0] far_1_1573_0;    relay_conn far_1_1573_0_a(.in(layer_0[866]), .out(far_1_1573_0[0]));    relay_conn far_1_1573_0_b(.in(layer_0[992]), .out(far_1_1573_0[1]));
    wire [1:0] far_1_1573_1;    relay_conn far_1_1573_1_a(.in(far_1_1573_0[0]), .out(far_1_1573_1[0]));    relay_conn far_1_1573_1_b(.in(far_1_1573_0[1]), .out(far_1_1573_1[1]));
    wire [1:0] far_1_1573_2;    relay_conn far_1_1573_2_a(.in(far_1_1573_1[0]), .out(far_1_1573_2[0]));    relay_conn far_1_1573_2_b(.in(far_1_1573_1[1]), .out(far_1_1573_2[1]));
    assign layer_1[553] = ~far_1_1573_2[1]; 
    wire [1:0] far_1_1574_0;    relay_conn far_1_1574_0_a(.in(layer_0[579]), .out(far_1_1574_0[0]));    relay_conn far_1_1574_0_b(.in(layer_0[704]), .out(far_1_1574_0[1]));
    wire [1:0] far_1_1574_1;    relay_conn far_1_1574_1_a(.in(far_1_1574_0[0]), .out(far_1_1574_1[0]));    relay_conn far_1_1574_1_b(.in(far_1_1574_0[1]), .out(far_1_1574_1[1]));
    wire [1:0] far_1_1574_2;    relay_conn far_1_1574_2_a(.in(far_1_1574_1[0]), .out(far_1_1574_2[0]));    relay_conn far_1_1574_2_b(.in(far_1_1574_1[1]), .out(far_1_1574_2[1]));
    assign layer_1[554] = ~(far_1_1574_2[0] | far_1_1574_2[1]); 
    assign layer_1[555] = layer_0[591]; 
    wire [1:0] far_1_1576_0;    relay_conn far_1_1576_0_a(.in(layer_0[992]), .out(far_1_1576_0[0]));    relay_conn far_1_1576_0_b(.in(layer_0[916]), .out(far_1_1576_0[1]));
    wire [1:0] far_1_1576_1;    relay_conn far_1_1576_1_a(.in(far_1_1576_0[0]), .out(far_1_1576_1[0]));    relay_conn far_1_1576_1_b(.in(far_1_1576_0[1]), .out(far_1_1576_1[1]));
    assign layer_1[556] = ~(far_1_1576_1[0] | far_1_1576_1[1]); 
    wire [1:0] far_1_1577_0;    relay_conn far_1_1577_0_a(.in(layer_0[530]), .out(far_1_1577_0[0]));    relay_conn far_1_1577_0_b(.in(layer_0[600]), .out(far_1_1577_0[1]));
    wire [1:0] far_1_1577_1;    relay_conn far_1_1577_1_a(.in(far_1_1577_0[0]), .out(far_1_1577_1[0]));    relay_conn far_1_1577_1_b(.in(far_1_1577_0[1]), .out(far_1_1577_1[1]));
    assign layer_1[557] = far_1_1577_1[0]; 
    wire [1:0] far_1_1578_0;    relay_conn far_1_1578_0_a(.in(layer_0[272]), .out(far_1_1578_0[0]));    relay_conn far_1_1578_0_b(.in(layer_0[208]), .out(far_1_1578_0[1]));
    wire [1:0] far_1_1578_1;    relay_conn far_1_1578_1_a(.in(far_1_1578_0[0]), .out(far_1_1578_1[0]));    relay_conn far_1_1578_1_b(.in(far_1_1578_0[1]), .out(far_1_1578_1[1]));
    assign layer_1[558] = ~(far_1_1578_1[0] | far_1_1578_1[1]); 
    assign layer_1[559] = ~(layer_0[626] | layer_0[640]); 
    wire [1:0] far_1_1580_0;    relay_conn far_1_1580_0_a(.in(layer_0[644]), .out(far_1_1580_0[0]));    relay_conn far_1_1580_0_b(.in(layer_0[606]), .out(far_1_1580_0[1]));
    assign layer_1[560] = ~(far_1_1580_0[0] & far_1_1580_0[1]); 
    wire [1:0] far_1_1581_0;    relay_conn far_1_1581_0_a(.in(layer_0[65]), .out(far_1_1581_0[0]));    relay_conn far_1_1581_0_b(.in(layer_0[147]), .out(far_1_1581_0[1]));
    wire [1:0] far_1_1581_1;    relay_conn far_1_1581_1_a(.in(far_1_1581_0[0]), .out(far_1_1581_1[0]));    relay_conn far_1_1581_1_b(.in(far_1_1581_0[1]), .out(far_1_1581_1[1]));
    assign layer_1[561] = ~(far_1_1581_1[0] | far_1_1581_1[1]); 
    wire [1:0] far_1_1582_0;    relay_conn far_1_1582_0_a(.in(layer_0[731]), .out(far_1_1582_0[0]));    relay_conn far_1_1582_0_b(.in(layer_0[807]), .out(far_1_1582_0[1]));
    wire [1:0] far_1_1582_1;    relay_conn far_1_1582_1_a(.in(far_1_1582_0[0]), .out(far_1_1582_1[0]));    relay_conn far_1_1582_1_b(.in(far_1_1582_0[1]), .out(far_1_1582_1[1]));
    assign layer_1[562] = ~far_1_1582_1[0] | (far_1_1582_1[0] & far_1_1582_1[1]); 
    assign layer_1[563] = ~(layer_0[967] & layer_0[966]); 
    assign layer_1[564] = layer_0[442] & ~layer_0[420]; 
    wire [1:0] far_1_1585_0;    relay_conn far_1_1585_0_a(.in(layer_0[21]), .out(far_1_1585_0[0]));    relay_conn far_1_1585_0_b(.in(layer_0[84]), .out(far_1_1585_0[1]));
    assign layer_1[565] = ~(far_1_1585_0[0] ^ far_1_1585_0[1]); 
    wire [1:0] far_1_1586_0;    relay_conn far_1_1586_0_a(.in(layer_0[14]), .out(far_1_1586_0[0]));    relay_conn far_1_1586_0_b(.in(layer_0[126]), .out(far_1_1586_0[1]));
    wire [1:0] far_1_1586_1;    relay_conn far_1_1586_1_a(.in(far_1_1586_0[0]), .out(far_1_1586_1[0]));    relay_conn far_1_1586_1_b(.in(far_1_1586_0[1]), .out(far_1_1586_1[1]));
    wire [1:0] far_1_1586_2;    relay_conn far_1_1586_2_a(.in(far_1_1586_1[0]), .out(far_1_1586_2[0]));    relay_conn far_1_1586_2_b(.in(far_1_1586_1[1]), .out(far_1_1586_2[1]));
    assign layer_1[566] = ~far_1_1586_2[1]; 
    wire [1:0] far_1_1587_0;    relay_conn far_1_1587_0_a(.in(layer_0[699]), .out(far_1_1587_0[0]));    relay_conn far_1_1587_0_b(.in(layer_0[644]), .out(far_1_1587_0[1]));
    assign layer_1[567] = ~(far_1_1587_0[0] ^ far_1_1587_0[1]); 
    wire [1:0] far_1_1588_0;    relay_conn far_1_1588_0_a(.in(layer_0[998]), .out(far_1_1588_0[0]));    relay_conn far_1_1588_0_b(.in(layer_0[914]), .out(far_1_1588_0[1]));
    wire [1:0] far_1_1588_1;    relay_conn far_1_1588_1_a(.in(far_1_1588_0[0]), .out(far_1_1588_1[0]));    relay_conn far_1_1588_1_b(.in(far_1_1588_0[1]), .out(far_1_1588_1[1]));
    assign layer_1[568] = far_1_1588_1[0]; 
    wire [1:0] far_1_1589_0;    relay_conn far_1_1589_0_a(.in(layer_0[336]), .out(far_1_1589_0[0]));    relay_conn far_1_1589_0_b(.in(layer_0[461]), .out(far_1_1589_0[1]));
    wire [1:0] far_1_1589_1;    relay_conn far_1_1589_1_a(.in(far_1_1589_0[0]), .out(far_1_1589_1[0]));    relay_conn far_1_1589_1_b(.in(far_1_1589_0[1]), .out(far_1_1589_1[1]));
    wire [1:0] far_1_1589_2;    relay_conn far_1_1589_2_a(.in(far_1_1589_1[0]), .out(far_1_1589_2[0]));    relay_conn far_1_1589_2_b(.in(far_1_1589_1[1]), .out(far_1_1589_2[1]));
    assign layer_1[569] = ~(far_1_1589_2[0] | far_1_1589_2[1]); 
    wire [1:0] far_1_1590_0;    relay_conn far_1_1590_0_a(.in(layer_0[638]), .out(far_1_1590_0[0]));    relay_conn far_1_1590_0_b(.in(layer_0[528]), .out(far_1_1590_0[1]));
    wire [1:0] far_1_1590_1;    relay_conn far_1_1590_1_a(.in(far_1_1590_0[0]), .out(far_1_1590_1[0]));    relay_conn far_1_1590_1_b(.in(far_1_1590_0[1]), .out(far_1_1590_1[1]));
    wire [1:0] far_1_1590_2;    relay_conn far_1_1590_2_a(.in(far_1_1590_1[0]), .out(far_1_1590_2[0]));    relay_conn far_1_1590_2_b(.in(far_1_1590_1[1]), .out(far_1_1590_2[1]));
    assign layer_1[570] = far_1_1590_2[1] & ~far_1_1590_2[0]; 
    wire [1:0] far_1_1591_0;    relay_conn far_1_1591_0_a(.in(layer_0[874]), .out(far_1_1591_0[0]));    relay_conn far_1_1591_0_b(.in(layer_0[789]), .out(far_1_1591_0[1]));
    wire [1:0] far_1_1591_1;    relay_conn far_1_1591_1_a(.in(far_1_1591_0[0]), .out(far_1_1591_1[0]));    relay_conn far_1_1591_1_b(.in(far_1_1591_0[1]), .out(far_1_1591_1[1]));
    assign layer_1[571] = far_1_1591_1[0] & far_1_1591_1[1]; 
    wire [1:0] far_1_1592_0;    relay_conn far_1_1592_0_a(.in(layer_0[914]), .out(far_1_1592_0[0]));    relay_conn far_1_1592_0_b(.in(layer_0[1012]), .out(far_1_1592_0[1]));
    wire [1:0] far_1_1592_1;    relay_conn far_1_1592_1_a(.in(far_1_1592_0[0]), .out(far_1_1592_1[0]));    relay_conn far_1_1592_1_b(.in(far_1_1592_0[1]), .out(far_1_1592_1[1]));
    wire [1:0] far_1_1592_2;    relay_conn far_1_1592_2_a(.in(far_1_1592_1[0]), .out(far_1_1592_2[0]));    relay_conn far_1_1592_2_b(.in(far_1_1592_1[1]), .out(far_1_1592_2[1]));
    assign layer_1[572] = ~(far_1_1592_2[0] & far_1_1592_2[1]); 
    wire [1:0] far_1_1593_0;    relay_conn far_1_1593_0_a(.in(layer_0[83]), .out(far_1_1593_0[0]));    relay_conn far_1_1593_0_b(.in(layer_0[194]), .out(far_1_1593_0[1]));
    wire [1:0] far_1_1593_1;    relay_conn far_1_1593_1_a(.in(far_1_1593_0[0]), .out(far_1_1593_1[0]));    relay_conn far_1_1593_1_b(.in(far_1_1593_0[1]), .out(far_1_1593_1[1]));
    wire [1:0] far_1_1593_2;    relay_conn far_1_1593_2_a(.in(far_1_1593_1[0]), .out(far_1_1593_2[0]));    relay_conn far_1_1593_2_b(.in(far_1_1593_1[1]), .out(far_1_1593_2[1]));
    assign layer_1[573] = ~(far_1_1593_2[0] | far_1_1593_2[1]); 
    wire [1:0] far_1_1594_0;    relay_conn far_1_1594_0_a(.in(layer_0[849]), .out(far_1_1594_0[0]));    relay_conn far_1_1594_0_b(.in(layer_0[752]), .out(far_1_1594_0[1]));
    wire [1:0] far_1_1594_1;    relay_conn far_1_1594_1_a(.in(far_1_1594_0[0]), .out(far_1_1594_1[0]));    relay_conn far_1_1594_1_b(.in(far_1_1594_0[1]), .out(far_1_1594_1[1]));
    wire [1:0] far_1_1594_2;    relay_conn far_1_1594_2_a(.in(far_1_1594_1[0]), .out(far_1_1594_2[0]));    relay_conn far_1_1594_2_b(.in(far_1_1594_1[1]), .out(far_1_1594_2[1]));
    assign layer_1[574] = ~(far_1_1594_2[0] & far_1_1594_2[1]); 
    assign layer_1[575] = ~(layer_0[625] | layer_0[601]); 
    wire [1:0] far_1_1596_0;    relay_conn far_1_1596_0_a(.in(layer_0[137]), .out(far_1_1596_0[0]));    relay_conn far_1_1596_0_b(.in(layer_0[193]), .out(far_1_1596_0[1]));
    assign layer_1[576] = far_1_1596_0[0]; 
    assign layer_1[577] = ~layer_0[1000] | (layer_0[1000] & layer_0[984]); 
    wire [1:0] far_1_1598_0;    relay_conn far_1_1598_0_a(.in(layer_0[252]), .out(far_1_1598_0[0]));    relay_conn far_1_1598_0_b(.in(layer_0[356]), .out(far_1_1598_0[1]));
    wire [1:0] far_1_1598_1;    relay_conn far_1_1598_1_a(.in(far_1_1598_0[0]), .out(far_1_1598_1[0]));    relay_conn far_1_1598_1_b(.in(far_1_1598_0[1]), .out(far_1_1598_1[1]));
    wire [1:0] far_1_1598_2;    relay_conn far_1_1598_2_a(.in(far_1_1598_1[0]), .out(far_1_1598_2[0]));    relay_conn far_1_1598_2_b(.in(far_1_1598_1[1]), .out(far_1_1598_2[1]));
    assign layer_1[578] = far_1_1598_2[0] & ~far_1_1598_2[1]; 
    wire [1:0] far_1_1599_0;    relay_conn far_1_1599_0_a(.in(layer_0[640]), .out(far_1_1599_0[0]));    relay_conn far_1_1599_0_b(.in(layer_0[731]), .out(far_1_1599_0[1]));
    wire [1:0] far_1_1599_1;    relay_conn far_1_1599_1_a(.in(far_1_1599_0[0]), .out(far_1_1599_1[0]));    relay_conn far_1_1599_1_b(.in(far_1_1599_0[1]), .out(far_1_1599_1[1]));
    assign layer_1[579] = ~(far_1_1599_1[0] | far_1_1599_1[1]); 
    wire [1:0] far_1_1600_0;    relay_conn far_1_1600_0_a(.in(layer_0[322]), .out(far_1_1600_0[0]));    relay_conn far_1_1600_0_b(.in(layer_0[272]), .out(far_1_1600_0[1]));
    assign layer_1[580] = far_1_1600_0[1]; 
    wire [1:0] far_1_1601_0;    relay_conn far_1_1601_0_a(.in(layer_0[299]), .out(far_1_1601_0[0]));    relay_conn far_1_1601_0_b(.in(layer_0[184]), .out(far_1_1601_0[1]));
    wire [1:0] far_1_1601_1;    relay_conn far_1_1601_1_a(.in(far_1_1601_0[0]), .out(far_1_1601_1[0]));    relay_conn far_1_1601_1_b(.in(far_1_1601_0[1]), .out(far_1_1601_1[1]));
    wire [1:0] far_1_1601_2;    relay_conn far_1_1601_2_a(.in(far_1_1601_1[0]), .out(far_1_1601_2[0]));    relay_conn far_1_1601_2_b(.in(far_1_1601_1[1]), .out(far_1_1601_2[1]));
    assign layer_1[581] = far_1_1601_2[1] & ~far_1_1601_2[0]; 
    wire [1:0] far_1_1602_0;    relay_conn far_1_1602_0_a(.in(layer_0[551]), .out(far_1_1602_0[0]));    relay_conn far_1_1602_0_b(.in(layer_0[679]), .out(far_1_1602_0[1]));
    wire [1:0] far_1_1602_1;    relay_conn far_1_1602_1_a(.in(far_1_1602_0[0]), .out(far_1_1602_1[0]));    relay_conn far_1_1602_1_b(.in(far_1_1602_0[1]), .out(far_1_1602_1[1]));
    wire [1:0] far_1_1602_2;    relay_conn far_1_1602_2_a(.in(far_1_1602_1[0]), .out(far_1_1602_2[0]));    relay_conn far_1_1602_2_b(.in(far_1_1602_1[1]), .out(far_1_1602_2[1]));
    wire [1:0] far_1_1602_3;    relay_conn far_1_1602_3_a(.in(far_1_1602_2[0]), .out(far_1_1602_3[0]));    relay_conn far_1_1602_3_b(.in(far_1_1602_2[1]), .out(far_1_1602_3[1]));
    assign layer_1[582] = far_1_1602_3[0] | far_1_1602_3[1]; 
    wire [1:0] far_1_1603_0;    relay_conn far_1_1603_0_a(.in(layer_0[886]), .out(far_1_1603_0[0]));    relay_conn far_1_1603_0_b(.in(layer_0[938]), .out(far_1_1603_0[1]));
    assign layer_1[583] = ~far_1_1603_0[0]; 
    wire [1:0] far_1_1604_0;    relay_conn far_1_1604_0_a(.in(layer_0[629]), .out(far_1_1604_0[0]));    relay_conn far_1_1604_0_b(.in(layer_0[596]), .out(far_1_1604_0[1]));
    assign layer_1[584] = ~far_1_1604_0[1] | (far_1_1604_0[0] & far_1_1604_0[1]); 
    wire [1:0] far_1_1605_0;    relay_conn far_1_1605_0_a(.in(layer_0[32]), .out(far_1_1605_0[0]));    relay_conn far_1_1605_0_b(.in(layer_0[99]), .out(far_1_1605_0[1]));
    wire [1:0] far_1_1605_1;    relay_conn far_1_1605_1_a(.in(far_1_1605_0[0]), .out(far_1_1605_1[0]));    relay_conn far_1_1605_1_b(.in(far_1_1605_0[1]), .out(far_1_1605_1[1]));
    assign layer_1[585] = far_1_1605_1[0] & ~far_1_1605_1[1]; 
    wire [1:0] far_1_1606_0;    relay_conn far_1_1606_0_a(.in(layer_0[408]), .out(far_1_1606_0[0]));    relay_conn far_1_1606_0_b(.in(layer_0[480]), .out(far_1_1606_0[1]));
    wire [1:0] far_1_1606_1;    relay_conn far_1_1606_1_a(.in(far_1_1606_0[0]), .out(far_1_1606_1[0]));    relay_conn far_1_1606_1_b(.in(far_1_1606_0[1]), .out(far_1_1606_1[1]));
    assign layer_1[586] = far_1_1606_1[0] & ~far_1_1606_1[1]; 
    wire [1:0] far_1_1607_0;    relay_conn far_1_1607_0_a(.in(layer_0[770]), .out(far_1_1607_0[0]));    relay_conn far_1_1607_0_b(.in(layer_0[659]), .out(far_1_1607_0[1]));
    wire [1:0] far_1_1607_1;    relay_conn far_1_1607_1_a(.in(far_1_1607_0[0]), .out(far_1_1607_1[0]));    relay_conn far_1_1607_1_b(.in(far_1_1607_0[1]), .out(far_1_1607_1[1]));
    wire [1:0] far_1_1607_2;    relay_conn far_1_1607_2_a(.in(far_1_1607_1[0]), .out(far_1_1607_2[0]));    relay_conn far_1_1607_2_b(.in(far_1_1607_1[1]), .out(far_1_1607_2[1]));
    assign layer_1[587] = far_1_1607_2[0] ^ far_1_1607_2[1]; 
    wire [1:0] far_1_1608_0;    relay_conn far_1_1608_0_a(.in(layer_0[334]), .out(far_1_1608_0[0]));    relay_conn far_1_1608_0_b(.in(layer_0[443]), .out(far_1_1608_0[1]));
    wire [1:0] far_1_1608_1;    relay_conn far_1_1608_1_a(.in(far_1_1608_0[0]), .out(far_1_1608_1[0]));    relay_conn far_1_1608_1_b(.in(far_1_1608_0[1]), .out(far_1_1608_1[1]));
    wire [1:0] far_1_1608_2;    relay_conn far_1_1608_2_a(.in(far_1_1608_1[0]), .out(far_1_1608_2[0]));    relay_conn far_1_1608_2_b(.in(far_1_1608_1[1]), .out(far_1_1608_2[1]));
    assign layer_1[588] = far_1_1608_2[0] & ~far_1_1608_2[1]; 
    wire [1:0] far_1_1609_0;    relay_conn far_1_1609_0_a(.in(layer_0[721]), .out(far_1_1609_0[0]));    relay_conn far_1_1609_0_b(.in(layer_0[833]), .out(far_1_1609_0[1]));
    wire [1:0] far_1_1609_1;    relay_conn far_1_1609_1_a(.in(far_1_1609_0[0]), .out(far_1_1609_1[0]));    relay_conn far_1_1609_1_b(.in(far_1_1609_0[1]), .out(far_1_1609_1[1]));
    wire [1:0] far_1_1609_2;    relay_conn far_1_1609_2_a(.in(far_1_1609_1[0]), .out(far_1_1609_2[0]));    relay_conn far_1_1609_2_b(.in(far_1_1609_1[1]), .out(far_1_1609_2[1]));
    assign layer_1[589] = far_1_1609_2[0] ^ far_1_1609_2[1]; 
    wire [1:0] far_1_1610_0;    relay_conn far_1_1610_0_a(.in(layer_0[683]), .out(far_1_1610_0[0]));    relay_conn far_1_1610_0_b(.in(layer_0[562]), .out(far_1_1610_0[1]));
    wire [1:0] far_1_1610_1;    relay_conn far_1_1610_1_a(.in(far_1_1610_0[0]), .out(far_1_1610_1[0]));    relay_conn far_1_1610_1_b(.in(far_1_1610_0[1]), .out(far_1_1610_1[1]));
    wire [1:0] far_1_1610_2;    relay_conn far_1_1610_2_a(.in(far_1_1610_1[0]), .out(far_1_1610_2[0]));    relay_conn far_1_1610_2_b(.in(far_1_1610_1[1]), .out(far_1_1610_2[1]));
    assign layer_1[590] = ~far_1_1610_2[1]; 
    wire [1:0] far_1_1611_0;    relay_conn far_1_1611_0_a(.in(layer_0[432]), .out(far_1_1611_0[0]));    relay_conn far_1_1611_0_b(.in(layer_0[485]), .out(far_1_1611_0[1]));
    assign layer_1[591] = far_1_1611_0[0] & far_1_1611_0[1]; 
    wire [1:0] far_1_1612_0;    relay_conn far_1_1612_0_a(.in(layer_0[480]), .out(far_1_1612_0[0]));    relay_conn far_1_1612_0_b(.in(layer_0[397]), .out(far_1_1612_0[1]));
    wire [1:0] far_1_1612_1;    relay_conn far_1_1612_1_a(.in(far_1_1612_0[0]), .out(far_1_1612_1[0]));    relay_conn far_1_1612_1_b(.in(far_1_1612_0[1]), .out(far_1_1612_1[1]));
    assign layer_1[592] = ~(far_1_1612_1[0] | far_1_1612_1[1]); 
    assign layer_1[593] = ~(layer_0[723] & layer_0[752]); 
    wire [1:0] far_1_1614_0;    relay_conn far_1_1614_0_a(.in(layer_0[1]), .out(far_1_1614_0[0]));    relay_conn far_1_1614_0_b(.in(layer_0[37]), .out(far_1_1614_0[1]));
    assign layer_1[594] = far_1_1614_0[0] ^ far_1_1614_0[1]; 
    wire [1:0] far_1_1615_0;    relay_conn far_1_1615_0_a(.in(layer_0[780]), .out(far_1_1615_0[0]));    relay_conn far_1_1615_0_b(.in(layer_0[834]), .out(far_1_1615_0[1]));
    assign layer_1[595] = far_1_1615_0[0]; 
    assign layer_1[596] = layer_0[202] | layer_0[204]; 
    assign layer_1[597] = ~(layer_0[773] & layer_0[790]); 
    wire [1:0] far_1_1618_0;    relay_conn far_1_1618_0_a(.in(layer_0[761]), .out(far_1_1618_0[0]));    relay_conn far_1_1618_0_b(.in(layer_0[708]), .out(far_1_1618_0[1]));
    assign layer_1[598] = ~far_1_1618_0[1] | (far_1_1618_0[0] & far_1_1618_0[1]); 
    wire [1:0] far_1_1619_0;    relay_conn far_1_1619_0_a(.in(layer_0[272]), .out(far_1_1619_0[0]));    relay_conn far_1_1619_0_b(.in(layer_0[329]), .out(far_1_1619_0[1]));
    assign layer_1[599] = far_1_1619_0[0] | far_1_1619_0[1]; 
    assign layer_1[600] = layer_0[346] & layer_0[361]; 
    wire [1:0] far_1_1621_0;    relay_conn far_1_1621_0_a(.in(layer_0[125]), .out(far_1_1621_0[0]));    relay_conn far_1_1621_0_b(.in(layer_0[205]), .out(far_1_1621_0[1]));
    wire [1:0] far_1_1621_1;    relay_conn far_1_1621_1_a(.in(far_1_1621_0[0]), .out(far_1_1621_1[0]));    relay_conn far_1_1621_1_b(.in(far_1_1621_0[1]), .out(far_1_1621_1[1]));
    assign layer_1[601] = ~(far_1_1621_1[0] & far_1_1621_1[1]); 
    wire [1:0] far_1_1622_0;    relay_conn far_1_1622_0_a(.in(layer_0[505]), .out(far_1_1622_0[0]));    relay_conn far_1_1622_0_b(.in(layer_0[389]), .out(far_1_1622_0[1]));
    wire [1:0] far_1_1622_1;    relay_conn far_1_1622_1_a(.in(far_1_1622_0[0]), .out(far_1_1622_1[0]));    relay_conn far_1_1622_1_b(.in(far_1_1622_0[1]), .out(far_1_1622_1[1]));
    wire [1:0] far_1_1622_2;    relay_conn far_1_1622_2_a(.in(far_1_1622_1[0]), .out(far_1_1622_2[0]));    relay_conn far_1_1622_2_b(.in(far_1_1622_1[1]), .out(far_1_1622_2[1]));
    assign layer_1[602] = far_1_1622_2[1] & ~far_1_1622_2[0]; 
    wire [1:0] far_1_1623_0;    relay_conn far_1_1623_0_a(.in(layer_0[511]), .out(far_1_1623_0[0]));    relay_conn far_1_1623_0_b(.in(layer_0[406]), .out(far_1_1623_0[1]));
    wire [1:0] far_1_1623_1;    relay_conn far_1_1623_1_a(.in(far_1_1623_0[0]), .out(far_1_1623_1[0]));    relay_conn far_1_1623_1_b(.in(far_1_1623_0[1]), .out(far_1_1623_1[1]));
    wire [1:0] far_1_1623_2;    relay_conn far_1_1623_2_a(.in(far_1_1623_1[0]), .out(far_1_1623_2[0]));    relay_conn far_1_1623_2_b(.in(far_1_1623_1[1]), .out(far_1_1623_2[1]));
    assign layer_1[603] = far_1_1623_2[0] | far_1_1623_2[1]; 
    assign layer_1[604] = layer_0[330] & ~layer_0[351]; 
    wire [1:0] far_1_1625_0;    relay_conn far_1_1625_0_a(.in(layer_0[489]), .out(far_1_1625_0[0]));    relay_conn far_1_1625_0_b(.in(layer_0[450]), .out(far_1_1625_0[1]));
    assign layer_1[605] = ~(far_1_1625_0[0] | far_1_1625_0[1]); 
    wire [1:0] far_1_1626_0;    relay_conn far_1_1626_0_a(.in(layer_0[614]), .out(far_1_1626_0[0]));    relay_conn far_1_1626_0_b(.in(layer_0[569]), .out(far_1_1626_0[1]));
    assign layer_1[606] = ~(far_1_1626_0[0] & far_1_1626_0[1]); 
    assign layer_1[607] = ~layer_0[374] | (layer_0[374] & layer_0[395]); 
    wire [1:0] far_1_1628_0;    relay_conn far_1_1628_0_a(.in(layer_0[452]), .out(far_1_1628_0[0]));    relay_conn far_1_1628_0_b(.in(layer_0[547]), .out(far_1_1628_0[1]));
    wire [1:0] far_1_1628_1;    relay_conn far_1_1628_1_a(.in(far_1_1628_0[0]), .out(far_1_1628_1[0]));    relay_conn far_1_1628_1_b(.in(far_1_1628_0[1]), .out(far_1_1628_1[1]));
    assign layer_1[608] = ~far_1_1628_1[0]; 
    wire [1:0] far_1_1629_0;    relay_conn far_1_1629_0_a(.in(layer_0[174]), .out(far_1_1629_0[0]));    relay_conn far_1_1629_0_b(.in(layer_0[119]), .out(far_1_1629_0[1]));
    assign layer_1[609] = ~far_1_1629_0[1] | (far_1_1629_0[0] & far_1_1629_0[1]); 
    assign layer_1[610] = ~(layer_0[315] | layer_0[343]); 
    wire [1:0] far_1_1631_0;    relay_conn far_1_1631_0_a(.in(layer_0[841]), .out(far_1_1631_0[0]));    relay_conn far_1_1631_0_b(.in(layer_0[793]), .out(far_1_1631_0[1]));
    assign layer_1[611] = ~far_1_1631_0[0]; 
    wire [1:0] far_1_1632_0;    relay_conn far_1_1632_0_a(.in(layer_0[512]), .out(far_1_1632_0[0]));    relay_conn far_1_1632_0_b(.in(layer_0[441]), .out(far_1_1632_0[1]));
    wire [1:0] far_1_1632_1;    relay_conn far_1_1632_1_a(.in(far_1_1632_0[0]), .out(far_1_1632_1[0]));    relay_conn far_1_1632_1_b(.in(far_1_1632_0[1]), .out(far_1_1632_1[1]));
    assign layer_1[612] = ~far_1_1632_1[0]; 
    wire [1:0] far_1_1633_0;    relay_conn far_1_1633_0_a(.in(layer_0[847]), .out(far_1_1633_0[0]));    relay_conn far_1_1633_0_b(.in(layer_0[926]), .out(far_1_1633_0[1]));
    wire [1:0] far_1_1633_1;    relay_conn far_1_1633_1_a(.in(far_1_1633_0[0]), .out(far_1_1633_1[0]));    relay_conn far_1_1633_1_b(.in(far_1_1633_0[1]), .out(far_1_1633_1[1]));
    assign layer_1[613] = ~far_1_1633_1[1] | (far_1_1633_1[0] & far_1_1633_1[1]); 
    wire [1:0] far_1_1634_0;    relay_conn far_1_1634_0_a(.in(layer_0[1010]), .out(far_1_1634_0[0]));    relay_conn far_1_1634_0_b(.in(layer_0[893]), .out(far_1_1634_0[1]));
    wire [1:0] far_1_1634_1;    relay_conn far_1_1634_1_a(.in(far_1_1634_0[0]), .out(far_1_1634_1[0]));    relay_conn far_1_1634_1_b(.in(far_1_1634_0[1]), .out(far_1_1634_1[1]));
    wire [1:0] far_1_1634_2;    relay_conn far_1_1634_2_a(.in(far_1_1634_1[0]), .out(far_1_1634_2[0]));    relay_conn far_1_1634_2_b(.in(far_1_1634_1[1]), .out(far_1_1634_2[1]));
    assign layer_1[614] = far_1_1634_2[1] & ~far_1_1634_2[0]; 
    wire [1:0] far_1_1635_0;    relay_conn far_1_1635_0_a(.in(layer_0[198]), .out(far_1_1635_0[0]));    relay_conn far_1_1635_0_b(.in(layer_0[282]), .out(far_1_1635_0[1]));
    wire [1:0] far_1_1635_1;    relay_conn far_1_1635_1_a(.in(far_1_1635_0[0]), .out(far_1_1635_1[0]));    relay_conn far_1_1635_1_b(.in(far_1_1635_0[1]), .out(far_1_1635_1[1]));
    assign layer_1[615] = ~(far_1_1635_1[0] & far_1_1635_1[1]); 
    wire [1:0] far_1_1636_0;    relay_conn far_1_1636_0_a(.in(layer_0[699]), .out(far_1_1636_0[0]));    relay_conn far_1_1636_0_b(.in(layer_0[768]), .out(far_1_1636_0[1]));
    wire [1:0] far_1_1636_1;    relay_conn far_1_1636_1_a(.in(far_1_1636_0[0]), .out(far_1_1636_1[0]));    relay_conn far_1_1636_1_b(.in(far_1_1636_0[1]), .out(far_1_1636_1[1]));
    assign layer_1[616] = ~far_1_1636_1[0]; 
    assign layer_1[617] = ~layer_0[923] | (layer_0[945] & layer_0[923]); 
    wire [1:0] far_1_1638_0;    relay_conn far_1_1638_0_a(.in(layer_0[367]), .out(far_1_1638_0[0]));    relay_conn far_1_1638_0_b(.in(layer_0[444]), .out(far_1_1638_0[1]));
    wire [1:0] far_1_1638_1;    relay_conn far_1_1638_1_a(.in(far_1_1638_0[0]), .out(far_1_1638_1[0]));    relay_conn far_1_1638_1_b(.in(far_1_1638_0[1]), .out(far_1_1638_1[1]));
    assign layer_1[618] = ~far_1_1638_1[1] | (far_1_1638_1[0] & far_1_1638_1[1]); 
    assign layer_1[619] = layer_0[66] | layer_0[71]; 
    wire [1:0] far_1_1640_0;    relay_conn far_1_1640_0_a(.in(layer_0[562]), .out(far_1_1640_0[0]));    relay_conn far_1_1640_0_b(.in(layer_0[446]), .out(far_1_1640_0[1]));
    wire [1:0] far_1_1640_1;    relay_conn far_1_1640_1_a(.in(far_1_1640_0[0]), .out(far_1_1640_1[0]));    relay_conn far_1_1640_1_b(.in(far_1_1640_0[1]), .out(far_1_1640_1[1]));
    wire [1:0] far_1_1640_2;    relay_conn far_1_1640_2_a(.in(far_1_1640_1[0]), .out(far_1_1640_2[0]));    relay_conn far_1_1640_2_b(.in(far_1_1640_1[1]), .out(far_1_1640_2[1]));
    assign layer_1[620] = ~far_1_1640_2[0] | (far_1_1640_2[0] & far_1_1640_2[1]); 
    assign layer_1[621] = layer_0[57] & ~layer_0[85]; 
    wire [1:0] far_1_1642_0;    relay_conn far_1_1642_0_a(.in(layer_0[493]), .out(far_1_1642_0[0]));    relay_conn far_1_1642_0_b(.in(layer_0[397]), .out(far_1_1642_0[1]));
    wire [1:0] far_1_1642_1;    relay_conn far_1_1642_1_a(.in(far_1_1642_0[0]), .out(far_1_1642_1[0]));    relay_conn far_1_1642_1_b(.in(far_1_1642_0[1]), .out(far_1_1642_1[1]));
    wire [1:0] far_1_1642_2;    relay_conn far_1_1642_2_a(.in(far_1_1642_1[0]), .out(far_1_1642_2[0]));    relay_conn far_1_1642_2_b(.in(far_1_1642_1[1]), .out(far_1_1642_2[1]));
    assign layer_1[622] = far_1_1642_2[0]; 
    assign layer_1[623] = layer_0[629]; 
    wire [1:0] far_1_1644_0;    relay_conn far_1_1644_0_a(.in(layer_0[356]), .out(far_1_1644_0[0]));    relay_conn far_1_1644_0_b(.in(layer_0[245]), .out(far_1_1644_0[1]));
    wire [1:0] far_1_1644_1;    relay_conn far_1_1644_1_a(.in(far_1_1644_0[0]), .out(far_1_1644_1[0]));    relay_conn far_1_1644_1_b(.in(far_1_1644_0[1]), .out(far_1_1644_1[1]));
    wire [1:0] far_1_1644_2;    relay_conn far_1_1644_2_a(.in(far_1_1644_1[0]), .out(far_1_1644_2[0]));    relay_conn far_1_1644_2_b(.in(far_1_1644_1[1]), .out(far_1_1644_2[1]));
    assign layer_1[624] = far_1_1644_2[1]; 
    wire [1:0] far_1_1645_0;    relay_conn far_1_1645_0_a(.in(layer_0[475]), .out(far_1_1645_0[0]));    relay_conn far_1_1645_0_b(.in(layer_0[438]), .out(far_1_1645_0[1]));
    assign layer_1[625] = far_1_1645_0[0] ^ far_1_1645_0[1]; 
    assign layer_1[626] = ~layer_0[640] | (layer_0[669] & layer_0[640]); 
    wire [1:0] far_1_1647_0;    relay_conn far_1_1647_0_a(.in(layer_0[973]), .out(far_1_1647_0[0]));    relay_conn far_1_1647_0_b(.in(layer_0[936]), .out(far_1_1647_0[1]));
    assign layer_1[627] = ~far_1_1647_0[0] | (far_1_1647_0[0] & far_1_1647_0[1]); 
    wire [1:0] far_1_1648_0;    relay_conn far_1_1648_0_a(.in(layer_0[881]), .out(far_1_1648_0[0]));    relay_conn far_1_1648_0_b(.in(layer_0[841]), .out(far_1_1648_0[1]));
    assign layer_1[628] = far_1_1648_0[0] & far_1_1648_0[1]; 
    wire [1:0] far_1_1649_0;    relay_conn far_1_1649_0_a(.in(layer_0[461]), .out(far_1_1649_0[0]));    relay_conn far_1_1649_0_b(.in(layer_0[361]), .out(far_1_1649_0[1]));
    wire [1:0] far_1_1649_1;    relay_conn far_1_1649_1_a(.in(far_1_1649_0[0]), .out(far_1_1649_1[0]));    relay_conn far_1_1649_1_b(.in(far_1_1649_0[1]), .out(far_1_1649_1[1]));
    wire [1:0] far_1_1649_2;    relay_conn far_1_1649_2_a(.in(far_1_1649_1[0]), .out(far_1_1649_2[0]));    relay_conn far_1_1649_2_b(.in(far_1_1649_1[1]), .out(far_1_1649_2[1]));
    assign layer_1[629] = ~far_1_1649_2[0]; 
    assign layer_1[630] = ~layer_0[438] | (layer_0[438] & layer_0[468]); 
    wire [1:0] far_1_1651_0;    relay_conn far_1_1651_0_a(.in(layer_0[387]), .out(far_1_1651_0[0]));    relay_conn far_1_1651_0_b(.in(layer_0[316]), .out(far_1_1651_0[1]));
    wire [1:0] far_1_1651_1;    relay_conn far_1_1651_1_a(.in(far_1_1651_0[0]), .out(far_1_1651_1[0]));    relay_conn far_1_1651_1_b(.in(far_1_1651_0[1]), .out(far_1_1651_1[1]));
    assign layer_1[631] = ~far_1_1651_1[0] | (far_1_1651_1[0] & far_1_1651_1[1]); 
    assign layer_1[632] = ~layer_0[604]; 
    wire [1:0] far_1_1653_0;    relay_conn far_1_1653_0_a(.in(layer_0[220]), .out(far_1_1653_0[0]));    relay_conn far_1_1653_0_b(.in(layer_0[115]), .out(far_1_1653_0[1]));
    wire [1:0] far_1_1653_1;    relay_conn far_1_1653_1_a(.in(far_1_1653_0[0]), .out(far_1_1653_1[0]));    relay_conn far_1_1653_1_b(.in(far_1_1653_0[1]), .out(far_1_1653_1[1]));
    wire [1:0] far_1_1653_2;    relay_conn far_1_1653_2_a(.in(far_1_1653_1[0]), .out(far_1_1653_2[0]));    relay_conn far_1_1653_2_b(.in(far_1_1653_1[1]), .out(far_1_1653_2[1]));
    assign layer_1[633] = far_1_1653_2[1]; 
    wire [1:0] far_1_1654_0;    relay_conn far_1_1654_0_a(.in(layer_0[173]), .out(far_1_1654_0[0]));    relay_conn far_1_1654_0_b(.in(layer_0[85]), .out(far_1_1654_0[1]));
    wire [1:0] far_1_1654_1;    relay_conn far_1_1654_1_a(.in(far_1_1654_0[0]), .out(far_1_1654_1[0]));    relay_conn far_1_1654_1_b(.in(far_1_1654_0[1]), .out(far_1_1654_1[1]));
    assign layer_1[634] = far_1_1654_1[0] & ~far_1_1654_1[1]; 
    assign layer_1[635] = layer_0[843] | layer_0[861]; 
    wire [1:0] far_1_1656_0;    relay_conn far_1_1656_0_a(.in(layer_0[686]), .out(far_1_1656_0[0]));    relay_conn far_1_1656_0_b(.in(layer_0[599]), .out(far_1_1656_0[1]));
    wire [1:0] far_1_1656_1;    relay_conn far_1_1656_1_a(.in(far_1_1656_0[0]), .out(far_1_1656_1[0]));    relay_conn far_1_1656_1_b(.in(far_1_1656_0[1]), .out(far_1_1656_1[1]));
    assign layer_1[636] = far_1_1656_1[0]; 
    assign layer_1[637] = layer_0[1019] & layer_0[988]; 
    wire [1:0] far_1_1658_0;    relay_conn far_1_1658_0_a(.in(layer_0[468]), .out(far_1_1658_0[0]));    relay_conn far_1_1658_0_b(.in(layer_0[432]), .out(far_1_1658_0[1]));
    assign layer_1[638] = far_1_1658_0[0] ^ far_1_1658_0[1]; 
    wire [1:0] far_1_1659_0;    relay_conn far_1_1659_0_a(.in(layer_0[799]), .out(far_1_1659_0[0]));    relay_conn far_1_1659_0_b(.in(layer_0[699]), .out(far_1_1659_0[1]));
    wire [1:0] far_1_1659_1;    relay_conn far_1_1659_1_a(.in(far_1_1659_0[0]), .out(far_1_1659_1[0]));    relay_conn far_1_1659_1_b(.in(far_1_1659_0[1]), .out(far_1_1659_1[1]));
    wire [1:0] far_1_1659_2;    relay_conn far_1_1659_2_a(.in(far_1_1659_1[0]), .out(far_1_1659_2[0]));    relay_conn far_1_1659_2_b(.in(far_1_1659_1[1]), .out(far_1_1659_2[1]));
    assign layer_1[639] = far_1_1659_2[1] & ~far_1_1659_2[0]; 
    wire [1:0] far_1_1660_0;    relay_conn far_1_1660_0_a(.in(layer_0[237]), .out(far_1_1660_0[0]));    relay_conn far_1_1660_0_b(.in(layer_0[287]), .out(far_1_1660_0[1]));
    assign layer_1[640] = ~far_1_1660_0[1]; 
    wire [1:0] far_1_1661_0;    relay_conn far_1_1661_0_a(.in(layer_0[876]), .out(far_1_1661_0[0]));    relay_conn far_1_1661_0_b(.in(layer_0[999]), .out(far_1_1661_0[1]));
    wire [1:0] far_1_1661_1;    relay_conn far_1_1661_1_a(.in(far_1_1661_0[0]), .out(far_1_1661_1[0]));    relay_conn far_1_1661_1_b(.in(far_1_1661_0[1]), .out(far_1_1661_1[1]));
    wire [1:0] far_1_1661_2;    relay_conn far_1_1661_2_a(.in(far_1_1661_1[0]), .out(far_1_1661_2[0]));    relay_conn far_1_1661_2_b(.in(far_1_1661_1[1]), .out(far_1_1661_2[1]));
    assign layer_1[641] = far_1_1661_2[1] & ~far_1_1661_2[0]; 
    wire [1:0] far_1_1662_0;    relay_conn far_1_1662_0_a(.in(layer_0[621]), .out(far_1_1662_0[0]));    relay_conn far_1_1662_0_b(.in(layer_0[579]), .out(far_1_1662_0[1]));
    assign layer_1[642] = ~far_1_1662_0[1] | (far_1_1662_0[0] & far_1_1662_0[1]); 
    assign layer_1[643] = layer_0[656]; 
    wire [1:0] far_1_1664_0;    relay_conn far_1_1664_0_a(.in(layer_0[285]), .out(far_1_1664_0[0]));    relay_conn far_1_1664_0_b(.in(layer_0[194]), .out(far_1_1664_0[1]));
    wire [1:0] far_1_1664_1;    relay_conn far_1_1664_1_a(.in(far_1_1664_0[0]), .out(far_1_1664_1[0]));    relay_conn far_1_1664_1_b(.in(far_1_1664_0[1]), .out(far_1_1664_1[1]));
    assign layer_1[644] = ~(far_1_1664_1[0] & far_1_1664_1[1]); 
    wire [1:0] far_1_1665_0;    relay_conn far_1_1665_0_a(.in(layer_0[178]), .out(far_1_1665_0[0]));    relay_conn far_1_1665_0_b(.in(layer_0[117]), .out(far_1_1665_0[1]));
    assign layer_1[645] = far_1_1665_0[1] & ~far_1_1665_0[0]; 
    wire [1:0] far_1_1666_0;    relay_conn far_1_1666_0_a(.in(layer_0[690]), .out(far_1_1666_0[0]));    relay_conn far_1_1666_0_b(.in(layer_0[741]), .out(far_1_1666_0[1]));
    assign layer_1[646] = far_1_1666_0[1] & ~far_1_1666_0[0]; 
    wire [1:0] far_1_1667_0;    relay_conn far_1_1667_0_a(.in(layer_0[756]), .out(far_1_1667_0[0]));    relay_conn far_1_1667_0_b(.in(layer_0[821]), .out(far_1_1667_0[1]));
    wire [1:0] far_1_1667_1;    relay_conn far_1_1667_1_a(.in(far_1_1667_0[0]), .out(far_1_1667_1[0]));    relay_conn far_1_1667_1_b(.in(far_1_1667_0[1]), .out(far_1_1667_1[1]));
    assign layer_1[647] = ~(far_1_1667_1[0] & far_1_1667_1[1]); 
    assign layer_1[648] = ~layer_0[728] | (layer_0[728] & layer_0[698]); 
    wire [1:0] far_1_1669_0;    relay_conn far_1_1669_0_a(.in(layer_0[672]), .out(far_1_1669_0[0]));    relay_conn far_1_1669_0_b(.in(layer_0[793]), .out(far_1_1669_0[1]));
    wire [1:0] far_1_1669_1;    relay_conn far_1_1669_1_a(.in(far_1_1669_0[0]), .out(far_1_1669_1[0]));    relay_conn far_1_1669_1_b(.in(far_1_1669_0[1]), .out(far_1_1669_1[1]));
    wire [1:0] far_1_1669_2;    relay_conn far_1_1669_2_a(.in(far_1_1669_1[0]), .out(far_1_1669_2[0]));    relay_conn far_1_1669_2_b(.in(far_1_1669_1[1]), .out(far_1_1669_2[1]));
    assign layer_1[649] = far_1_1669_2[1] & ~far_1_1669_2[0]; 
    wire [1:0] far_1_1670_0;    relay_conn far_1_1670_0_a(.in(layer_0[107]), .out(far_1_1670_0[0]));    relay_conn far_1_1670_0_b(.in(layer_0[204]), .out(far_1_1670_0[1]));
    wire [1:0] far_1_1670_1;    relay_conn far_1_1670_1_a(.in(far_1_1670_0[0]), .out(far_1_1670_1[0]));    relay_conn far_1_1670_1_b(.in(far_1_1670_0[1]), .out(far_1_1670_1[1]));
    wire [1:0] far_1_1670_2;    relay_conn far_1_1670_2_a(.in(far_1_1670_1[0]), .out(far_1_1670_2[0]));    relay_conn far_1_1670_2_b(.in(far_1_1670_1[1]), .out(far_1_1670_2[1]));
    assign layer_1[650] = ~far_1_1670_2[0]; 
    assign layer_1[651] = ~(layer_0[973] & layer_0[995]); 
    wire [1:0] far_1_1672_0;    relay_conn far_1_1672_0_a(.in(layer_0[400]), .out(far_1_1672_0[0]));    relay_conn far_1_1672_0_b(.in(layer_0[514]), .out(far_1_1672_0[1]));
    wire [1:0] far_1_1672_1;    relay_conn far_1_1672_1_a(.in(far_1_1672_0[0]), .out(far_1_1672_1[0]));    relay_conn far_1_1672_1_b(.in(far_1_1672_0[1]), .out(far_1_1672_1[1]));
    wire [1:0] far_1_1672_2;    relay_conn far_1_1672_2_a(.in(far_1_1672_1[0]), .out(far_1_1672_2[0]));    relay_conn far_1_1672_2_b(.in(far_1_1672_1[1]), .out(far_1_1672_2[1]));
    assign layer_1[652] = far_1_1672_2[0] | far_1_1672_2[1]; 
    wire [1:0] far_1_1673_0;    relay_conn far_1_1673_0_a(.in(layer_0[699]), .out(far_1_1673_0[0]));    relay_conn far_1_1673_0_b(.in(layer_0[815]), .out(far_1_1673_0[1]));
    wire [1:0] far_1_1673_1;    relay_conn far_1_1673_1_a(.in(far_1_1673_0[0]), .out(far_1_1673_1[0]));    relay_conn far_1_1673_1_b(.in(far_1_1673_0[1]), .out(far_1_1673_1[1]));
    wire [1:0] far_1_1673_2;    relay_conn far_1_1673_2_a(.in(far_1_1673_1[0]), .out(far_1_1673_2[0]));    relay_conn far_1_1673_2_b(.in(far_1_1673_1[1]), .out(far_1_1673_2[1]));
    assign layer_1[653] = far_1_1673_2[0] & ~far_1_1673_2[1]; 
    wire [1:0] far_1_1674_0;    relay_conn far_1_1674_0_a(.in(layer_0[911]), .out(far_1_1674_0[0]));    relay_conn far_1_1674_0_b(.in(layer_0[846]), .out(far_1_1674_0[1]));
    wire [1:0] far_1_1674_1;    relay_conn far_1_1674_1_a(.in(far_1_1674_0[0]), .out(far_1_1674_1[0]));    relay_conn far_1_1674_1_b(.in(far_1_1674_0[1]), .out(far_1_1674_1[1]));
    assign layer_1[654] = ~(far_1_1674_1[0] | far_1_1674_1[1]); 
    wire [1:0] far_1_1675_0;    relay_conn far_1_1675_0_a(.in(layer_0[754]), .out(far_1_1675_0[0]));    relay_conn far_1_1675_0_b(.in(layer_0[656]), .out(far_1_1675_0[1]));
    wire [1:0] far_1_1675_1;    relay_conn far_1_1675_1_a(.in(far_1_1675_0[0]), .out(far_1_1675_1[0]));    relay_conn far_1_1675_1_b(.in(far_1_1675_0[1]), .out(far_1_1675_1[1]));
    wire [1:0] far_1_1675_2;    relay_conn far_1_1675_2_a(.in(far_1_1675_1[0]), .out(far_1_1675_2[0]));    relay_conn far_1_1675_2_b(.in(far_1_1675_1[1]), .out(far_1_1675_2[1]));
    assign layer_1[655] = ~far_1_1675_2[1]; 
    wire [1:0] far_1_1676_0;    relay_conn far_1_1676_0_a(.in(layer_0[734]), .out(far_1_1676_0[0]));    relay_conn far_1_1676_0_b(.in(layer_0[795]), .out(far_1_1676_0[1]));
    assign layer_1[656] = ~far_1_1676_0[0]; 
    assign layer_1[657] = ~layer_0[455] | (layer_0[478] & layer_0[455]); 
    wire [1:0] far_1_1678_0;    relay_conn far_1_1678_0_a(.in(layer_0[361]), .out(far_1_1678_0[0]));    relay_conn far_1_1678_0_b(.in(layer_0[441]), .out(far_1_1678_0[1]));
    wire [1:0] far_1_1678_1;    relay_conn far_1_1678_1_a(.in(far_1_1678_0[0]), .out(far_1_1678_1[0]));    relay_conn far_1_1678_1_b(.in(far_1_1678_0[1]), .out(far_1_1678_1[1]));
    assign layer_1[658] = far_1_1678_1[0] ^ far_1_1678_1[1]; 
    wire [1:0] far_1_1679_0;    relay_conn far_1_1679_0_a(.in(layer_0[75]), .out(far_1_1679_0[0]));    relay_conn far_1_1679_0_b(.in(layer_0[131]), .out(far_1_1679_0[1]));
    assign layer_1[659] = far_1_1679_0[0] | far_1_1679_0[1]; 
    wire [1:0] far_1_1680_0;    relay_conn far_1_1680_0_a(.in(layer_0[91]), .out(far_1_1680_0[0]));    relay_conn far_1_1680_0_b(.in(layer_0[188]), .out(far_1_1680_0[1]));
    wire [1:0] far_1_1680_1;    relay_conn far_1_1680_1_a(.in(far_1_1680_0[0]), .out(far_1_1680_1[0]));    relay_conn far_1_1680_1_b(.in(far_1_1680_0[1]), .out(far_1_1680_1[1]));
    wire [1:0] far_1_1680_2;    relay_conn far_1_1680_2_a(.in(far_1_1680_1[0]), .out(far_1_1680_2[0]));    relay_conn far_1_1680_2_b(.in(far_1_1680_1[1]), .out(far_1_1680_2[1]));
    assign layer_1[660] = ~(far_1_1680_2[0] | far_1_1680_2[1]); 
    wire [1:0] far_1_1681_0;    relay_conn far_1_1681_0_a(.in(layer_0[883]), .out(far_1_1681_0[0]));    relay_conn far_1_1681_0_b(.in(layer_0[947]), .out(far_1_1681_0[1]));
    wire [1:0] far_1_1681_1;    relay_conn far_1_1681_1_a(.in(far_1_1681_0[0]), .out(far_1_1681_1[0]));    relay_conn far_1_1681_1_b(.in(far_1_1681_0[1]), .out(far_1_1681_1[1]));
    assign layer_1[661] = far_1_1681_1[0]; 
    wire [1:0] far_1_1682_0;    relay_conn far_1_1682_0_a(.in(layer_0[185]), .out(far_1_1682_0[0]));    relay_conn far_1_1682_0_b(.in(layer_0[107]), .out(far_1_1682_0[1]));
    wire [1:0] far_1_1682_1;    relay_conn far_1_1682_1_a(.in(far_1_1682_0[0]), .out(far_1_1682_1[0]));    relay_conn far_1_1682_1_b(.in(far_1_1682_0[1]), .out(far_1_1682_1[1]));
    assign layer_1[662] = far_1_1682_1[1] & ~far_1_1682_1[0]; 
    assign layer_1[663] = ~layer_0[942] | (layer_0[942] & layer_0[938]); 
    assign layer_1[664] = ~layer_0[73]; 
    wire [1:0] far_1_1685_0;    relay_conn far_1_1685_0_a(.in(layer_0[404]), .out(far_1_1685_0[0]));    relay_conn far_1_1685_0_b(.in(layer_0[505]), .out(far_1_1685_0[1]));
    wire [1:0] far_1_1685_1;    relay_conn far_1_1685_1_a(.in(far_1_1685_0[0]), .out(far_1_1685_1[0]));    relay_conn far_1_1685_1_b(.in(far_1_1685_0[1]), .out(far_1_1685_1[1]));
    wire [1:0] far_1_1685_2;    relay_conn far_1_1685_2_a(.in(far_1_1685_1[0]), .out(far_1_1685_2[0]));    relay_conn far_1_1685_2_b(.in(far_1_1685_1[1]), .out(far_1_1685_2[1]));
    assign layer_1[665] = ~(far_1_1685_2[0] | far_1_1685_2[1]); 
    wire [1:0] far_1_1686_0;    relay_conn far_1_1686_0_a(.in(layer_0[412]), .out(far_1_1686_0[0]));    relay_conn far_1_1686_0_b(.in(layer_0[468]), .out(far_1_1686_0[1]));
    assign layer_1[666] = far_1_1686_0[1]; 
    assign layer_1[667] = layer_0[366]; 
    wire [1:0] far_1_1688_0;    relay_conn far_1_1688_0_a(.in(layer_0[280]), .out(far_1_1688_0[0]));    relay_conn far_1_1688_0_b(.in(layer_0[356]), .out(far_1_1688_0[1]));
    wire [1:0] far_1_1688_1;    relay_conn far_1_1688_1_a(.in(far_1_1688_0[0]), .out(far_1_1688_1[0]));    relay_conn far_1_1688_1_b(.in(far_1_1688_0[1]), .out(far_1_1688_1[1]));
    assign layer_1[668] = far_1_1688_1[0] | far_1_1688_1[1]; 
    wire [1:0] far_1_1689_0;    relay_conn far_1_1689_0_a(.in(layer_0[656]), .out(far_1_1689_0[0]));    relay_conn far_1_1689_0_b(.in(layer_0[588]), .out(far_1_1689_0[1]));
    wire [1:0] far_1_1689_1;    relay_conn far_1_1689_1_a(.in(far_1_1689_0[0]), .out(far_1_1689_1[0]));    relay_conn far_1_1689_1_b(.in(far_1_1689_0[1]), .out(far_1_1689_1[1]));
    assign layer_1[669] = ~far_1_1689_1[1]; 
    assign layer_1[670] = ~layer_0[397] | (layer_0[415] & layer_0[397]); 
    wire [1:0] far_1_1691_0;    relay_conn far_1_1691_0_a(.in(layer_0[525]), .out(far_1_1691_0[0]));    relay_conn far_1_1691_0_b(.in(layer_0[562]), .out(far_1_1691_0[1]));
    assign layer_1[671] = ~far_1_1691_0[0] | (far_1_1691_0[0] & far_1_1691_0[1]); 
    wire [1:0] far_1_1692_0;    relay_conn far_1_1692_0_a(.in(layer_0[125]), .out(far_1_1692_0[0]));    relay_conn far_1_1692_0_b(.in(layer_0[242]), .out(far_1_1692_0[1]));
    wire [1:0] far_1_1692_1;    relay_conn far_1_1692_1_a(.in(far_1_1692_0[0]), .out(far_1_1692_1[0]));    relay_conn far_1_1692_1_b(.in(far_1_1692_0[1]), .out(far_1_1692_1[1]));
    wire [1:0] far_1_1692_2;    relay_conn far_1_1692_2_a(.in(far_1_1692_1[0]), .out(far_1_1692_2[0]));    relay_conn far_1_1692_2_b(.in(far_1_1692_1[1]), .out(far_1_1692_2[1]));
    assign layer_1[672] = ~far_1_1692_2[0]; 
    wire [1:0] far_1_1693_0;    relay_conn far_1_1693_0_a(.in(layer_0[723]), .out(far_1_1693_0[0]));    relay_conn far_1_1693_0_b(.in(layer_0[768]), .out(far_1_1693_0[1]));
    assign layer_1[673] = ~(far_1_1693_0[0] | far_1_1693_0[1]); 
    assign layer_1[674] = layer_0[400] & ~layer_0[392]; 
    wire [1:0] far_1_1695_0;    relay_conn far_1_1695_0_a(.in(layer_0[26]), .out(far_1_1695_0[0]));    relay_conn far_1_1695_0_b(.in(layer_0[80]), .out(far_1_1695_0[1]));
    assign layer_1[675] = far_1_1695_0[0] & far_1_1695_0[1]; 
    wire [1:0] far_1_1696_0;    relay_conn far_1_1696_0_a(.in(layer_0[372]), .out(far_1_1696_0[0]));    relay_conn far_1_1696_0_b(.in(layer_0[314]), .out(far_1_1696_0[1]));
    assign layer_1[676] = ~far_1_1696_0[1]; 
    wire [1:0] far_1_1697_0;    relay_conn far_1_1697_0_a(.in(layer_0[1019]), .out(far_1_1697_0[0]));    relay_conn far_1_1697_0_b(.in(layer_0[916]), .out(far_1_1697_0[1]));
    wire [1:0] far_1_1697_1;    relay_conn far_1_1697_1_a(.in(far_1_1697_0[0]), .out(far_1_1697_1[0]));    relay_conn far_1_1697_1_b(.in(far_1_1697_0[1]), .out(far_1_1697_1[1]));
    wire [1:0] far_1_1697_2;    relay_conn far_1_1697_2_a(.in(far_1_1697_1[0]), .out(far_1_1697_2[0]));    relay_conn far_1_1697_2_b(.in(far_1_1697_1[1]), .out(far_1_1697_2[1]));
    assign layer_1[677] = ~(far_1_1697_2[0] & far_1_1697_2[1]); 
    wire [1:0] far_1_1698_0;    relay_conn far_1_1698_0_a(.in(layer_0[241]), .out(far_1_1698_0[0]));    relay_conn far_1_1698_0_b(.in(layer_0[360]), .out(far_1_1698_0[1]));
    wire [1:0] far_1_1698_1;    relay_conn far_1_1698_1_a(.in(far_1_1698_0[0]), .out(far_1_1698_1[0]));    relay_conn far_1_1698_1_b(.in(far_1_1698_0[1]), .out(far_1_1698_1[1]));
    wire [1:0] far_1_1698_2;    relay_conn far_1_1698_2_a(.in(far_1_1698_1[0]), .out(far_1_1698_2[0]));    relay_conn far_1_1698_2_b(.in(far_1_1698_1[1]), .out(far_1_1698_2[1]));
    assign layer_1[678] = far_1_1698_2[1]; 
    wire [1:0] far_1_1699_0;    relay_conn far_1_1699_0_a(.in(layer_0[299]), .out(far_1_1699_0[0]));    relay_conn far_1_1699_0_b(.in(layer_0[175]), .out(far_1_1699_0[1]));
    wire [1:0] far_1_1699_1;    relay_conn far_1_1699_1_a(.in(far_1_1699_0[0]), .out(far_1_1699_1[0]));    relay_conn far_1_1699_1_b(.in(far_1_1699_0[1]), .out(far_1_1699_1[1]));
    wire [1:0] far_1_1699_2;    relay_conn far_1_1699_2_a(.in(far_1_1699_1[0]), .out(far_1_1699_2[0]));    relay_conn far_1_1699_2_b(.in(far_1_1699_1[1]), .out(far_1_1699_2[1]));
    assign layer_1[679] = ~far_1_1699_2[0] | (far_1_1699_2[0] & far_1_1699_2[1]); 
    wire [1:0] far_1_1700_0;    relay_conn far_1_1700_0_a(.in(layer_0[732]), .out(far_1_1700_0[0]));    relay_conn far_1_1700_0_b(.in(layer_0[768]), .out(far_1_1700_0[1]));
    assign layer_1[680] = ~far_1_1700_0[1] | (far_1_1700_0[0] & far_1_1700_0[1]); 
    wire [1:0] far_1_1701_0;    relay_conn far_1_1701_0_a(.in(layer_0[351]), .out(far_1_1701_0[0]));    relay_conn far_1_1701_0_b(.in(layer_0[237]), .out(far_1_1701_0[1]));
    wire [1:0] far_1_1701_1;    relay_conn far_1_1701_1_a(.in(far_1_1701_0[0]), .out(far_1_1701_1[0]));    relay_conn far_1_1701_1_b(.in(far_1_1701_0[1]), .out(far_1_1701_1[1]));
    wire [1:0] far_1_1701_2;    relay_conn far_1_1701_2_a(.in(far_1_1701_1[0]), .out(far_1_1701_2[0]));    relay_conn far_1_1701_2_b(.in(far_1_1701_1[1]), .out(far_1_1701_2[1]));
    assign layer_1[681] = far_1_1701_2[0]; 
    wire [1:0] far_1_1702_0;    relay_conn far_1_1702_0_a(.in(layer_0[84]), .out(far_1_1702_0[0]));    relay_conn far_1_1702_0_b(.in(layer_0[170]), .out(far_1_1702_0[1]));
    wire [1:0] far_1_1702_1;    relay_conn far_1_1702_1_a(.in(far_1_1702_0[0]), .out(far_1_1702_1[0]));    relay_conn far_1_1702_1_b(.in(far_1_1702_0[1]), .out(far_1_1702_1[1]));
    assign layer_1[682] = far_1_1702_1[1]; 
    wire [1:0] far_1_1703_0;    relay_conn far_1_1703_0_a(.in(layer_0[719]), .out(far_1_1703_0[0]));    relay_conn far_1_1703_0_b(.in(layer_0[837]), .out(far_1_1703_0[1]));
    wire [1:0] far_1_1703_1;    relay_conn far_1_1703_1_a(.in(far_1_1703_0[0]), .out(far_1_1703_1[0]));    relay_conn far_1_1703_1_b(.in(far_1_1703_0[1]), .out(far_1_1703_1[1]));
    wire [1:0] far_1_1703_2;    relay_conn far_1_1703_2_a(.in(far_1_1703_1[0]), .out(far_1_1703_2[0]));    relay_conn far_1_1703_2_b(.in(far_1_1703_1[1]), .out(far_1_1703_2[1]));
    assign layer_1[683] = ~(far_1_1703_2[0] & far_1_1703_2[1]); 
    wire [1:0] far_1_1704_0;    relay_conn far_1_1704_0_a(.in(layer_0[459]), .out(far_1_1704_0[0]));    relay_conn far_1_1704_0_b(.in(layer_0[336]), .out(far_1_1704_0[1]));
    wire [1:0] far_1_1704_1;    relay_conn far_1_1704_1_a(.in(far_1_1704_0[0]), .out(far_1_1704_1[0]));    relay_conn far_1_1704_1_b(.in(far_1_1704_0[1]), .out(far_1_1704_1[1]));
    wire [1:0] far_1_1704_2;    relay_conn far_1_1704_2_a(.in(far_1_1704_1[0]), .out(far_1_1704_2[0]));    relay_conn far_1_1704_2_b(.in(far_1_1704_1[1]), .out(far_1_1704_2[1]));
    assign layer_1[684] = ~far_1_1704_2[0]; 
    assign layer_1[685] = ~(layer_0[348] | layer_0[354]); 
    assign layer_1[686] = ~layer_0[954]; 
    assign layer_1[687] = ~(layer_0[156] | layer_0[185]); 
    wire [1:0] far_1_1708_0;    relay_conn far_1_1708_0_a(.in(layer_0[539]), .out(far_1_1708_0[0]));    relay_conn far_1_1708_0_b(.in(layer_0[504]), .out(far_1_1708_0[1]));
    assign layer_1[688] = ~far_1_1708_0[1]; 
    wire [1:0] far_1_1709_0;    relay_conn far_1_1709_0_a(.in(layer_0[942]), .out(far_1_1709_0[0]));    relay_conn far_1_1709_0_b(.in(layer_0[889]), .out(far_1_1709_0[1]));
    assign layer_1[689] = ~(far_1_1709_0[0] | far_1_1709_0[1]); 
    assign layer_1[690] = layer_0[623] & layer_0[630]; 
    wire [1:0] far_1_1711_0;    relay_conn far_1_1711_0_a(.in(layer_0[193]), .out(far_1_1711_0[0]));    relay_conn far_1_1711_0_b(.in(layer_0[149]), .out(far_1_1711_0[1]));
    assign layer_1[691] = ~far_1_1711_0[0] | (far_1_1711_0[0] & far_1_1711_0[1]); 
    wire [1:0] far_1_1712_0;    relay_conn far_1_1712_0_a(.in(layer_0[977]), .out(far_1_1712_0[0]));    relay_conn far_1_1712_0_b(.in(layer_0[909]), .out(far_1_1712_0[1]));
    wire [1:0] far_1_1712_1;    relay_conn far_1_1712_1_a(.in(far_1_1712_0[0]), .out(far_1_1712_1[0]));    relay_conn far_1_1712_1_b(.in(far_1_1712_0[1]), .out(far_1_1712_1[1]));
    assign layer_1[692] = far_1_1712_1[0] & far_1_1712_1[1]; 
    wire [1:0] far_1_1713_0;    relay_conn far_1_1713_0_a(.in(layer_0[799]), .out(far_1_1713_0[0]));    relay_conn far_1_1713_0_b(.in(layer_0[707]), .out(far_1_1713_0[1]));
    wire [1:0] far_1_1713_1;    relay_conn far_1_1713_1_a(.in(far_1_1713_0[0]), .out(far_1_1713_1[0]));    relay_conn far_1_1713_1_b(.in(far_1_1713_0[1]), .out(far_1_1713_1[1]));
    assign layer_1[693] = ~far_1_1713_1[0]; 
    assign layer_1[694] = layer_0[1011]; 
    assign layer_1[695] = layer_0[75] & layer_0[65]; 
    wire [1:0] far_1_1716_0;    relay_conn far_1_1716_0_a(.in(layer_0[246]), .out(far_1_1716_0[0]));    relay_conn far_1_1716_0_b(.in(layer_0[353]), .out(far_1_1716_0[1]));
    wire [1:0] far_1_1716_1;    relay_conn far_1_1716_1_a(.in(far_1_1716_0[0]), .out(far_1_1716_1[0]));    relay_conn far_1_1716_1_b(.in(far_1_1716_0[1]), .out(far_1_1716_1[1]));
    wire [1:0] far_1_1716_2;    relay_conn far_1_1716_2_a(.in(far_1_1716_1[0]), .out(far_1_1716_2[0]));    relay_conn far_1_1716_2_b(.in(far_1_1716_1[1]), .out(far_1_1716_2[1]));
    assign layer_1[696] = far_1_1716_2[0]; 
    wire [1:0] far_1_1717_0;    relay_conn far_1_1717_0_a(.in(layer_0[671]), .out(far_1_1717_0[0]));    relay_conn far_1_1717_0_b(.in(layer_0[736]), .out(far_1_1717_0[1]));
    wire [1:0] far_1_1717_1;    relay_conn far_1_1717_1_a(.in(far_1_1717_0[0]), .out(far_1_1717_1[0]));    relay_conn far_1_1717_1_b(.in(far_1_1717_0[1]), .out(far_1_1717_1[1]));
    assign layer_1[697] = far_1_1717_1[1] & ~far_1_1717_1[0]; 
    wire [1:0] far_1_1718_0;    relay_conn far_1_1718_0_a(.in(layer_0[80]), .out(far_1_1718_0[0]));    relay_conn far_1_1718_0_b(.in(layer_0[131]), .out(far_1_1718_0[1]));
    assign layer_1[698] = far_1_1718_0[1]; 
    wire [1:0] far_1_1719_0;    relay_conn far_1_1719_0_a(.in(layer_0[849]), .out(far_1_1719_0[0]));    relay_conn far_1_1719_0_b(.in(layer_0[816]), .out(far_1_1719_0[1]));
    assign layer_1[699] = ~(far_1_1719_0[0] & far_1_1719_0[1]); 
    wire [1:0] far_1_1720_0;    relay_conn far_1_1720_0_a(.in(layer_0[169]), .out(far_1_1720_0[0]));    relay_conn far_1_1720_0_b(.in(layer_0[65]), .out(far_1_1720_0[1]));
    wire [1:0] far_1_1720_1;    relay_conn far_1_1720_1_a(.in(far_1_1720_0[0]), .out(far_1_1720_1[0]));    relay_conn far_1_1720_1_b(.in(far_1_1720_0[1]), .out(far_1_1720_1[1]));
    wire [1:0] far_1_1720_2;    relay_conn far_1_1720_2_a(.in(far_1_1720_1[0]), .out(far_1_1720_2[0]));    relay_conn far_1_1720_2_b(.in(far_1_1720_1[1]), .out(far_1_1720_2[1]));
    assign layer_1[700] = far_1_1720_2[0] | far_1_1720_2[1]; 
    wire [1:0] far_1_1721_0;    relay_conn far_1_1721_0_a(.in(layer_0[762]), .out(far_1_1721_0[0]));    relay_conn far_1_1721_0_b(.in(layer_0[849]), .out(far_1_1721_0[1]));
    wire [1:0] far_1_1721_1;    relay_conn far_1_1721_1_a(.in(far_1_1721_0[0]), .out(far_1_1721_1[0]));    relay_conn far_1_1721_1_b(.in(far_1_1721_0[1]), .out(far_1_1721_1[1]));
    assign layer_1[701] = ~far_1_1721_1[1] | (far_1_1721_1[0] & far_1_1721_1[1]); 
    assign layer_1[702] = layer_0[855] & ~layer_0[854]; 
    wire [1:0] far_1_1723_0;    relay_conn far_1_1723_0_a(.in(layer_0[891]), .out(far_1_1723_0[0]));    relay_conn far_1_1723_0_b(.in(layer_0[958]), .out(far_1_1723_0[1]));
    wire [1:0] far_1_1723_1;    relay_conn far_1_1723_1_a(.in(far_1_1723_0[0]), .out(far_1_1723_1[0]));    relay_conn far_1_1723_1_b(.in(far_1_1723_0[1]), .out(far_1_1723_1[1]));
    assign layer_1[703] = far_1_1723_1[1] & ~far_1_1723_1[0]; 
    wire [1:0] far_1_1724_0;    relay_conn far_1_1724_0_a(.in(layer_0[95]), .out(far_1_1724_0[0]));    relay_conn far_1_1724_0_b(.in(layer_0[157]), .out(far_1_1724_0[1]));
    assign layer_1[704] = far_1_1724_0[0] & ~far_1_1724_0[1]; 
    wire [1:0] far_1_1725_0;    relay_conn far_1_1725_0_a(.in(layer_0[497]), .out(far_1_1725_0[0]));    relay_conn far_1_1725_0_b(.in(layer_0[559]), .out(far_1_1725_0[1]));
    assign layer_1[705] = ~far_1_1725_0[0]; 
    wire [1:0] far_1_1726_0;    relay_conn far_1_1726_0_a(.in(layer_0[111]), .out(far_1_1726_0[0]));    relay_conn far_1_1726_0_b(.in(layer_0[160]), .out(far_1_1726_0[1]));
    assign layer_1[706] = ~far_1_1726_0[1] | (far_1_1726_0[0] & far_1_1726_0[1]); 
    wire [1:0] far_1_1727_0;    relay_conn far_1_1727_0_a(.in(layer_0[949]), .out(far_1_1727_0[0]));    relay_conn far_1_1727_0_b(.in(layer_0[837]), .out(far_1_1727_0[1]));
    wire [1:0] far_1_1727_1;    relay_conn far_1_1727_1_a(.in(far_1_1727_0[0]), .out(far_1_1727_1[0]));    relay_conn far_1_1727_1_b(.in(far_1_1727_0[1]), .out(far_1_1727_1[1]));
    wire [1:0] far_1_1727_2;    relay_conn far_1_1727_2_a(.in(far_1_1727_1[0]), .out(far_1_1727_2[0]));    relay_conn far_1_1727_2_b(.in(far_1_1727_1[1]), .out(far_1_1727_2[1]));
    assign layer_1[707] = ~far_1_1727_2[1] | (far_1_1727_2[0] & far_1_1727_2[1]); 
    wire [1:0] far_1_1728_0;    relay_conn far_1_1728_0_a(.in(layer_0[957]), .out(far_1_1728_0[0]));    relay_conn far_1_1728_0_b(.in(layer_0[849]), .out(far_1_1728_0[1]));
    wire [1:0] far_1_1728_1;    relay_conn far_1_1728_1_a(.in(far_1_1728_0[0]), .out(far_1_1728_1[0]));    relay_conn far_1_1728_1_b(.in(far_1_1728_0[1]), .out(far_1_1728_1[1]));
    wire [1:0] far_1_1728_2;    relay_conn far_1_1728_2_a(.in(far_1_1728_1[0]), .out(far_1_1728_2[0]));    relay_conn far_1_1728_2_b(.in(far_1_1728_1[1]), .out(far_1_1728_2[1]));
    assign layer_1[708] = ~far_1_1728_2[1]; 
    wire [1:0] far_1_1729_0;    relay_conn far_1_1729_0_a(.in(layer_0[636]), .out(far_1_1729_0[0]));    relay_conn far_1_1729_0_b(.in(layer_0[599]), .out(far_1_1729_0[1]));
    assign layer_1[709] = ~far_1_1729_0[1] | (far_1_1729_0[0] & far_1_1729_0[1]); 
    assign layer_1[710] = layer_0[512]; 
    wire [1:0] far_1_1731_0;    relay_conn far_1_1731_0_a(.in(layer_0[815]), .out(far_1_1731_0[0]));    relay_conn far_1_1731_0_b(.in(layer_0[735]), .out(far_1_1731_0[1]));
    wire [1:0] far_1_1731_1;    relay_conn far_1_1731_1_a(.in(far_1_1731_0[0]), .out(far_1_1731_1[0]));    relay_conn far_1_1731_1_b(.in(far_1_1731_0[1]), .out(far_1_1731_1[1]));
    assign layer_1[711] = far_1_1731_1[0] ^ far_1_1731_1[1]; 
    wire [1:0] far_1_1732_0;    relay_conn far_1_1732_0_a(.in(layer_0[735]), .out(far_1_1732_0[0]));    relay_conn far_1_1732_0_b(.in(layer_0[698]), .out(far_1_1732_0[1]));
    assign layer_1[712] = far_1_1732_0[0] & far_1_1732_0[1]; 
    assign layer_1[713] = ~layer_0[51]; 
    assign layer_1[714] = ~(layer_0[62] & layer_0[49]); 
    wire [1:0] far_1_1735_0;    relay_conn far_1_1735_0_a(.in(layer_0[433]), .out(far_1_1735_0[0]));    relay_conn far_1_1735_0_b(.in(layer_0[395]), .out(far_1_1735_0[1]));
    assign layer_1[715] = far_1_1735_0[1] & ~far_1_1735_0[0]; 
    assign layer_1[716] = ~(layer_0[7] | layer_0[11]); 
    wire [1:0] far_1_1737_0;    relay_conn far_1_1737_0_a(.in(layer_0[676]), .out(far_1_1737_0[0]));    relay_conn far_1_1737_0_b(.in(layer_0[617]), .out(far_1_1737_0[1]));
    assign layer_1[717] = far_1_1737_0[0] & ~far_1_1737_0[1]; 
    assign layer_1[718] = ~(layer_0[938] | layer_0[942]); 
    wire [1:0] far_1_1739_0;    relay_conn far_1_1739_0_a(.in(layer_0[43]), .out(far_1_1739_0[0]));    relay_conn far_1_1739_0_b(.in(layer_0[91]), .out(far_1_1739_0[1]));
    assign layer_1[719] = ~far_1_1739_0[0]; 
    assign layer_1[720] = ~(layer_0[445] & layer_0[444]); 
    wire [1:0] far_1_1741_0;    relay_conn far_1_1741_0_a(.in(layer_0[120]), .out(far_1_1741_0[0]));    relay_conn far_1_1741_0_b(.in(layer_0[208]), .out(far_1_1741_0[1]));
    wire [1:0] far_1_1741_1;    relay_conn far_1_1741_1_a(.in(far_1_1741_0[0]), .out(far_1_1741_1[0]));    relay_conn far_1_1741_1_b(.in(far_1_1741_0[1]), .out(far_1_1741_1[1]));
    assign layer_1[721] = far_1_1741_1[1]; 
    wire [1:0] far_1_1742_0;    relay_conn far_1_1742_0_a(.in(layer_0[178]), .out(far_1_1742_0[0]));    relay_conn far_1_1742_0_b(.in(layer_0[93]), .out(far_1_1742_0[1]));
    wire [1:0] far_1_1742_1;    relay_conn far_1_1742_1_a(.in(far_1_1742_0[0]), .out(far_1_1742_1[0]));    relay_conn far_1_1742_1_b(.in(far_1_1742_0[1]), .out(far_1_1742_1[1]));
    assign layer_1[722] = ~far_1_1742_1[1]; 
    wire [1:0] far_1_1743_0;    relay_conn far_1_1743_0_a(.in(layer_0[368]), .out(far_1_1743_0[0]));    relay_conn far_1_1743_0_b(.in(layer_0[456]), .out(far_1_1743_0[1]));
    wire [1:0] far_1_1743_1;    relay_conn far_1_1743_1_a(.in(far_1_1743_0[0]), .out(far_1_1743_1[0]));    relay_conn far_1_1743_1_b(.in(far_1_1743_0[1]), .out(far_1_1743_1[1]));
    assign layer_1[723] = ~far_1_1743_1[1] | (far_1_1743_1[0] & far_1_1743_1[1]); 
    wire [1:0] far_1_1744_0;    relay_conn far_1_1744_0_a(.in(layer_0[887]), .out(far_1_1744_0[0]));    relay_conn far_1_1744_0_b(.in(layer_0[781]), .out(far_1_1744_0[1]));
    wire [1:0] far_1_1744_1;    relay_conn far_1_1744_1_a(.in(far_1_1744_0[0]), .out(far_1_1744_1[0]));    relay_conn far_1_1744_1_b(.in(far_1_1744_0[1]), .out(far_1_1744_1[1]));
    wire [1:0] far_1_1744_2;    relay_conn far_1_1744_2_a(.in(far_1_1744_1[0]), .out(far_1_1744_2[0]));    relay_conn far_1_1744_2_b(.in(far_1_1744_1[1]), .out(far_1_1744_2[1]));
    assign layer_1[724] = far_1_1744_2[0] & ~far_1_1744_2[1]; 
    wire [1:0] far_1_1745_0;    relay_conn far_1_1745_0_a(.in(layer_0[128]), .out(far_1_1745_0[0]));    relay_conn far_1_1745_0_b(.in(layer_0[182]), .out(far_1_1745_0[1]));
    assign layer_1[725] = ~(far_1_1745_0[0] ^ far_1_1745_0[1]); 
    assign layer_1[726] = layer_0[415] & layer_0[386]; 
    assign layer_1[727] = layer_0[996] ^ layer_0[1019]; 
    assign layer_1[728] = layer_0[521] & layer_0[514]; 
    wire [1:0] far_1_1749_0;    relay_conn far_1_1749_0_a(.in(layer_0[780]), .out(far_1_1749_0[0]));    relay_conn far_1_1749_0_b(.in(layer_0[891]), .out(far_1_1749_0[1]));
    wire [1:0] far_1_1749_1;    relay_conn far_1_1749_1_a(.in(far_1_1749_0[0]), .out(far_1_1749_1[0]));    relay_conn far_1_1749_1_b(.in(far_1_1749_0[1]), .out(far_1_1749_1[1]));
    wire [1:0] far_1_1749_2;    relay_conn far_1_1749_2_a(.in(far_1_1749_1[0]), .out(far_1_1749_2[0]));    relay_conn far_1_1749_2_b(.in(far_1_1749_1[1]), .out(far_1_1749_2[1]));
    assign layer_1[729] = far_1_1749_2[0] & far_1_1749_2[1]; 
    assign layer_1[730] = layer_0[874]; 
    wire [1:0] far_1_1751_0;    relay_conn far_1_1751_0_a(.in(layer_0[444]), .out(far_1_1751_0[0]));    relay_conn far_1_1751_0_b(.in(layer_0[329]), .out(far_1_1751_0[1]));
    wire [1:0] far_1_1751_1;    relay_conn far_1_1751_1_a(.in(far_1_1751_0[0]), .out(far_1_1751_1[0]));    relay_conn far_1_1751_1_b(.in(far_1_1751_0[1]), .out(far_1_1751_1[1]));
    wire [1:0] far_1_1751_2;    relay_conn far_1_1751_2_a(.in(far_1_1751_1[0]), .out(far_1_1751_2[0]));    relay_conn far_1_1751_2_b(.in(far_1_1751_1[1]), .out(far_1_1751_2[1]));
    assign layer_1[731] = far_1_1751_2[0] & ~far_1_1751_2[1]; 
    wire [1:0] far_1_1752_0;    relay_conn far_1_1752_0_a(.in(layer_0[395]), .out(far_1_1752_0[0]));    relay_conn far_1_1752_0_b(.in(layer_0[476]), .out(far_1_1752_0[1]));
    wire [1:0] far_1_1752_1;    relay_conn far_1_1752_1_a(.in(far_1_1752_0[0]), .out(far_1_1752_1[0]));    relay_conn far_1_1752_1_b(.in(far_1_1752_0[1]), .out(far_1_1752_1[1]));
    assign layer_1[732] = ~(far_1_1752_1[0] & far_1_1752_1[1]); 
    assign layer_1[733] = layer_0[62] & ~layer_0[57]; 
    wire [1:0] far_1_1754_0;    relay_conn far_1_1754_0_a(.in(layer_0[357]), .out(far_1_1754_0[0]));    relay_conn far_1_1754_0_b(.in(layer_0[395]), .out(far_1_1754_0[1]));
    assign layer_1[734] = far_1_1754_0[1] & ~far_1_1754_0[0]; 
    wire [1:0] far_1_1755_0;    relay_conn far_1_1755_0_a(.in(layer_0[514]), .out(far_1_1755_0[0]));    relay_conn far_1_1755_0_b(.in(layer_0[476]), .out(far_1_1755_0[1]));
    assign layer_1[735] = far_1_1755_0[1] & ~far_1_1755_0[0]; 
    assign layer_1[736] = layer_0[359] & ~layer_0[363]; 
    wire [1:0] far_1_1757_0;    relay_conn far_1_1757_0_a(.in(layer_0[301]), .out(far_1_1757_0[0]));    relay_conn far_1_1757_0_b(.in(layer_0[400]), .out(far_1_1757_0[1]));
    wire [1:0] far_1_1757_1;    relay_conn far_1_1757_1_a(.in(far_1_1757_0[0]), .out(far_1_1757_1[0]));    relay_conn far_1_1757_1_b(.in(far_1_1757_0[1]), .out(far_1_1757_1[1]));
    wire [1:0] far_1_1757_2;    relay_conn far_1_1757_2_a(.in(far_1_1757_1[0]), .out(far_1_1757_2[0]));    relay_conn far_1_1757_2_b(.in(far_1_1757_1[1]), .out(far_1_1757_2[1]));
    assign layer_1[737] = ~(far_1_1757_2[0] ^ far_1_1757_2[1]); 
    wire [1:0] far_1_1758_0;    relay_conn far_1_1758_0_a(.in(layer_0[233]), .out(far_1_1758_0[0]));    relay_conn far_1_1758_0_b(.in(layer_0[293]), .out(far_1_1758_0[1]));
    assign layer_1[738] = ~(far_1_1758_0[0] | far_1_1758_0[1]); 
    wire [1:0] far_1_1759_0;    relay_conn far_1_1759_0_a(.in(layer_0[329]), .out(far_1_1759_0[0]));    relay_conn far_1_1759_0_b(.in(layer_0[456]), .out(far_1_1759_0[1]));
    wire [1:0] far_1_1759_1;    relay_conn far_1_1759_1_a(.in(far_1_1759_0[0]), .out(far_1_1759_1[0]));    relay_conn far_1_1759_1_b(.in(far_1_1759_0[1]), .out(far_1_1759_1[1]));
    wire [1:0] far_1_1759_2;    relay_conn far_1_1759_2_a(.in(far_1_1759_1[0]), .out(far_1_1759_2[0]));    relay_conn far_1_1759_2_b(.in(far_1_1759_1[1]), .out(far_1_1759_2[1]));
    assign layer_1[739] = ~far_1_1759_2[1]; 
    assign layer_1[740] = layer_0[867] ^ layer_0[860]; 
    wire [1:0] far_1_1761_0;    relay_conn far_1_1761_0_a(.in(layer_0[867]), .out(far_1_1761_0[0]));    relay_conn far_1_1761_0_b(.in(layer_0[824]), .out(far_1_1761_0[1]));
    assign layer_1[741] = ~(far_1_1761_0[0] ^ far_1_1761_0[1]); 
    wire [1:0] far_1_1762_0;    relay_conn far_1_1762_0_a(.in(layer_0[587]), .out(far_1_1762_0[0]));    relay_conn far_1_1762_0_b(.in(layer_0[685]), .out(far_1_1762_0[1]));
    wire [1:0] far_1_1762_1;    relay_conn far_1_1762_1_a(.in(far_1_1762_0[0]), .out(far_1_1762_1[0]));    relay_conn far_1_1762_1_b(.in(far_1_1762_0[1]), .out(far_1_1762_1[1]));
    wire [1:0] far_1_1762_2;    relay_conn far_1_1762_2_a(.in(far_1_1762_1[0]), .out(far_1_1762_2[0]));    relay_conn far_1_1762_2_b(.in(far_1_1762_1[1]), .out(far_1_1762_2[1]));
    assign layer_1[742] = ~far_1_1762_2[0]; 
    wire [1:0] far_1_1763_0;    relay_conn far_1_1763_0_a(.in(layer_0[628]), .out(far_1_1763_0[0]));    relay_conn far_1_1763_0_b(.in(layer_0[686]), .out(far_1_1763_0[1]));
    assign layer_1[743] = far_1_1763_0[0] & ~far_1_1763_0[1]; 
    wire [1:0] far_1_1764_0;    relay_conn far_1_1764_0_a(.in(layer_0[174]), .out(far_1_1764_0[0]));    relay_conn far_1_1764_0_b(.in(layer_0[208]), .out(far_1_1764_0[1]));
    assign layer_1[744] = far_1_1764_0[0]; 
    assign layer_1[745] = layer_0[35]; 
    wire [1:0] far_1_1766_0;    relay_conn far_1_1766_0_a(.in(layer_0[590]), .out(far_1_1766_0[0]));    relay_conn far_1_1766_0_b(.in(layer_0[669]), .out(far_1_1766_0[1]));
    wire [1:0] far_1_1766_1;    relay_conn far_1_1766_1_a(.in(far_1_1766_0[0]), .out(far_1_1766_1[0]));    relay_conn far_1_1766_1_b(.in(far_1_1766_0[1]), .out(far_1_1766_1[1]));
    assign layer_1[746] = far_1_1766_1[0] & ~far_1_1766_1[1]; 
    wire [1:0] far_1_1767_0;    relay_conn far_1_1767_0_a(.in(layer_0[147]), .out(far_1_1767_0[0]));    relay_conn far_1_1767_0_b(.in(layer_0[240]), .out(far_1_1767_0[1]));
    wire [1:0] far_1_1767_1;    relay_conn far_1_1767_1_a(.in(far_1_1767_0[0]), .out(far_1_1767_1[0]));    relay_conn far_1_1767_1_b(.in(far_1_1767_0[1]), .out(far_1_1767_1[1]));
    assign layer_1[747] = ~far_1_1767_1[0]; 
    wire [1:0] far_1_1768_0;    relay_conn far_1_1768_0_a(.in(layer_0[849]), .out(far_1_1768_0[0]));    relay_conn far_1_1768_0_b(.in(layer_0[741]), .out(far_1_1768_0[1]));
    wire [1:0] far_1_1768_1;    relay_conn far_1_1768_1_a(.in(far_1_1768_0[0]), .out(far_1_1768_1[0]));    relay_conn far_1_1768_1_b(.in(far_1_1768_0[1]), .out(far_1_1768_1[1]));
    wire [1:0] far_1_1768_2;    relay_conn far_1_1768_2_a(.in(far_1_1768_1[0]), .out(far_1_1768_2[0]));    relay_conn far_1_1768_2_b(.in(far_1_1768_1[1]), .out(far_1_1768_2[1]));
    assign layer_1[748] = far_1_1768_2[1]; 
    assign layer_1[749] = ~layer_0[21]; 
    wire [1:0] far_1_1770_0;    relay_conn far_1_1770_0_a(.in(layer_0[756]), .out(far_1_1770_0[0]));    relay_conn far_1_1770_0_b(.in(layer_0[860]), .out(far_1_1770_0[1]));
    wire [1:0] far_1_1770_1;    relay_conn far_1_1770_1_a(.in(far_1_1770_0[0]), .out(far_1_1770_1[0]));    relay_conn far_1_1770_1_b(.in(far_1_1770_0[1]), .out(far_1_1770_1[1]));
    wire [1:0] far_1_1770_2;    relay_conn far_1_1770_2_a(.in(far_1_1770_1[0]), .out(far_1_1770_2[0]));    relay_conn far_1_1770_2_b(.in(far_1_1770_1[1]), .out(far_1_1770_2[1]));
    assign layer_1[750] = far_1_1770_2[0] | far_1_1770_2[1]; 
    wire [1:0] far_1_1771_0;    relay_conn far_1_1771_0_a(.in(layer_0[6]), .out(far_1_1771_0[0]));    relay_conn far_1_1771_0_b(.in(layer_0[99]), .out(far_1_1771_0[1]));
    wire [1:0] far_1_1771_1;    relay_conn far_1_1771_1_a(.in(far_1_1771_0[0]), .out(far_1_1771_1[0]));    relay_conn far_1_1771_1_b(.in(far_1_1771_0[1]), .out(far_1_1771_1[1]));
    assign layer_1[751] = far_1_1771_1[1] & ~far_1_1771_1[0]; 
    wire [1:0] far_1_1772_0;    relay_conn far_1_1772_0_a(.in(layer_0[237]), .out(far_1_1772_0[0]));    relay_conn far_1_1772_0_b(.in(layer_0[272]), .out(far_1_1772_0[1]));
    assign layer_1[752] = far_1_1772_0[0] & ~far_1_1772_0[1]; 
    wire [1:0] far_1_1773_0;    relay_conn far_1_1773_0_a(.in(layer_0[314]), .out(far_1_1773_0[0]));    relay_conn far_1_1773_0_b(.in(layer_0[422]), .out(far_1_1773_0[1]));
    wire [1:0] far_1_1773_1;    relay_conn far_1_1773_1_a(.in(far_1_1773_0[0]), .out(far_1_1773_1[0]));    relay_conn far_1_1773_1_b(.in(far_1_1773_0[1]), .out(far_1_1773_1[1]));
    wire [1:0] far_1_1773_2;    relay_conn far_1_1773_2_a(.in(far_1_1773_1[0]), .out(far_1_1773_2[0]));    relay_conn far_1_1773_2_b(.in(far_1_1773_1[1]), .out(far_1_1773_2[1]));
    assign layer_1[753] = far_1_1773_2[0]; 
    wire [1:0] far_1_1774_0;    relay_conn far_1_1774_0_a(.in(layer_0[429]), .out(far_1_1774_0[0]));    relay_conn far_1_1774_0_b(.in(layer_0[313]), .out(far_1_1774_0[1]));
    wire [1:0] far_1_1774_1;    relay_conn far_1_1774_1_a(.in(far_1_1774_0[0]), .out(far_1_1774_1[0]));    relay_conn far_1_1774_1_b(.in(far_1_1774_0[1]), .out(far_1_1774_1[1]));
    wire [1:0] far_1_1774_2;    relay_conn far_1_1774_2_a(.in(far_1_1774_1[0]), .out(far_1_1774_2[0]));    relay_conn far_1_1774_2_b(.in(far_1_1774_1[1]), .out(far_1_1774_2[1]));
    assign layer_1[754] = far_1_1774_2[0] ^ far_1_1774_2[1]; 
    wire [1:0] far_1_1775_0;    relay_conn far_1_1775_0_a(.in(layer_0[366]), .out(far_1_1775_0[0]));    relay_conn far_1_1775_0_b(.in(layer_0[299]), .out(far_1_1775_0[1]));
    wire [1:0] far_1_1775_1;    relay_conn far_1_1775_1_a(.in(far_1_1775_0[0]), .out(far_1_1775_1[0]));    relay_conn far_1_1775_1_b(.in(far_1_1775_0[1]), .out(far_1_1775_1[1]));
    assign layer_1[755] = far_1_1775_1[1]; 
    wire [1:0] far_1_1776_0;    relay_conn far_1_1776_0_a(.in(layer_0[205]), .out(far_1_1776_0[0]));    relay_conn far_1_1776_0_b(.in(layer_0[253]), .out(far_1_1776_0[1]));
    assign layer_1[756] = ~far_1_1776_0[0]; 
    wire [1:0] far_1_1777_0;    relay_conn far_1_1777_0_a(.in(layer_0[666]), .out(far_1_1777_0[0]));    relay_conn far_1_1777_0_b(.in(layer_0[579]), .out(far_1_1777_0[1]));
    wire [1:0] far_1_1777_1;    relay_conn far_1_1777_1_a(.in(far_1_1777_0[0]), .out(far_1_1777_1[0]));    relay_conn far_1_1777_1_b(.in(far_1_1777_0[1]), .out(far_1_1777_1[1]));
    assign layer_1[757] = ~(far_1_1777_1[0] | far_1_1777_1[1]); 
    wire [1:0] far_1_1778_0;    relay_conn far_1_1778_0_a(.in(layer_0[860]), .out(far_1_1778_0[0]));    relay_conn far_1_1778_0_b(.in(layer_0[906]), .out(far_1_1778_0[1]));
    assign layer_1[758] = far_1_1778_0[0]; 
    wire [1:0] far_1_1779_0;    relay_conn far_1_1779_0_a(.in(layer_0[887]), .out(far_1_1779_0[0]));    relay_conn far_1_1779_0_b(.in(layer_0[954]), .out(far_1_1779_0[1]));
    wire [1:0] far_1_1779_1;    relay_conn far_1_1779_1_a(.in(far_1_1779_0[0]), .out(far_1_1779_1[0]));    relay_conn far_1_1779_1_b(.in(far_1_1779_0[1]), .out(far_1_1779_1[1]));
    assign layer_1[759] = far_1_1779_1[0] | far_1_1779_1[1]; 
    wire [1:0] far_1_1780_0;    relay_conn far_1_1780_0_a(.in(layer_0[857]), .out(far_1_1780_0[0]));    relay_conn far_1_1780_0_b(.in(layer_0[770]), .out(far_1_1780_0[1]));
    wire [1:0] far_1_1780_1;    relay_conn far_1_1780_1_a(.in(far_1_1780_0[0]), .out(far_1_1780_1[0]));    relay_conn far_1_1780_1_b(.in(far_1_1780_0[1]), .out(far_1_1780_1[1]));
    assign layer_1[760] = ~far_1_1780_1[1] | (far_1_1780_1[0] & far_1_1780_1[1]); 
    wire [1:0] far_1_1781_0;    relay_conn far_1_1781_0_a(.in(layer_0[582]), .out(far_1_1781_0[0]));    relay_conn far_1_1781_0_b(.in(layer_0[621]), .out(far_1_1781_0[1]));
    assign layer_1[761] = far_1_1781_0[0] & far_1_1781_0[1]; 
    wire [1:0] far_1_1782_0;    relay_conn far_1_1782_0_a(.in(layer_0[415]), .out(far_1_1782_0[0]));    relay_conn far_1_1782_0_b(.in(layer_0[314]), .out(far_1_1782_0[1]));
    wire [1:0] far_1_1782_1;    relay_conn far_1_1782_1_a(.in(far_1_1782_0[0]), .out(far_1_1782_1[0]));    relay_conn far_1_1782_1_b(.in(far_1_1782_0[1]), .out(far_1_1782_1[1]));
    wire [1:0] far_1_1782_2;    relay_conn far_1_1782_2_a(.in(far_1_1782_1[0]), .out(far_1_1782_2[0]));    relay_conn far_1_1782_2_b(.in(far_1_1782_1[1]), .out(far_1_1782_2[1]));
    assign layer_1[762] = far_1_1782_2[0] | far_1_1782_2[1]; 
    assign layer_1[763] = ~layer_0[375] | (layer_0[375] & layer_0[396]); 
    assign layer_1[764] = layer_0[45] & ~layer_0[74]; 
    wire [1:0] far_1_1785_0;    relay_conn far_1_1785_0_a(.in(layer_0[430]), .out(far_1_1785_0[0]));    relay_conn far_1_1785_0_b(.in(layer_0[493]), .out(far_1_1785_0[1]));
    assign layer_1[765] = far_1_1785_0[1]; 
    wire [1:0] far_1_1786_0;    relay_conn far_1_1786_0_a(.in(layer_0[756]), .out(far_1_1786_0[0]));    relay_conn far_1_1786_0_b(.in(layer_0[856]), .out(far_1_1786_0[1]));
    wire [1:0] far_1_1786_1;    relay_conn far_1_1786_1_a(.in(far_1_1786_0[0]), .out(far_1_1786_1[0]));    relay_conn far_1_1786_1_b(.in(far_1_1786_0[1]), .out(far_1_1786_1[1]));
    wire [1:0] far_1_1786_2;    relay_conn far_1_1786_2_a(.in(far_1_1786_1[0]), .out(far_1_1786_2[0]));    relay_conn far_1_1786_2_b(.in(far_1_1786_1[1]), .out(far_1_1786_2[1]));
    assign layer_1[766] = far_1_1786_2[0]; 
    wire [1:0] far_1_1787_0;    relay_conn far_1_1787_0_a(.in(layer_0[786]), .out(far_1_1787_0[0]));    relay_conn far_1_1787_0_b(.in(layer_0[690]), .out(far_1_1787_0[1]));
    wire [1:0] far_1_1787_1;    relay_conn far_1_1787_1_a(.in(far_1_1787_0[0]), .out(far_1_1787_1[0]));    relay_conn far_1_1787_1_b(.in(far_1_1787_0[1]), .out(far_1_1787_1[1]));
    wire [1:0] far_1_1787_2;    relay_conn far_1_1787_2_a(.in(far_1_1787_1[0]), .out(far_1_1787_2[0]));    relay_conn far_1_1787_2_b(.in(far_1_1787_1[1]), .out(far_1_1787_2[1]));
    assign layer_1[767] = ~(far_1_1787_2[0] | far_1_1787_2[1]); 
    assign layer_1[768] = ~(layer_0[661] | layer_0[641]); 
    wire [1:0] far_1_1789_0;    relay_conn far_1_1789_0_a(.in(layer_0[397]), .out(far_1_1789_0[0]));    relay_conn far_1_1789_0_b(.in(layer_0[277]), .out(far_1_1789_0[1]));
    wire [1:0] far_1_1789_1;    relay_conn far_1_1789_1_a(.in(far_1_1789_0[0]), .out(far_1_1789_1[0]));    relay_conn far_1_1789_1_b(.in(far_1_1789_0[1]), .out(far_1_1789_1[1]));
    wire [1:0] far_1_1789_2;    relay_conn far_1_1789_2_a(.in(far_1_1789_1[0]), .out(far_1_1789_2[0]));    relay_conn far_1_1789_2_b(.in(far_1_1789_1[1]), .out(far_1_1789_2[1]));
    assign layer_1[769] = ~far_1_1789_2[0] | (far_1_1789_2[0] & far_1_1789_2[1]); 
    assign layer_1[770] = layer_0[834] & ~layer_0[839]; 
    wire [1:0] far_1_1791_0;    relay_conn far_1_1791_0_a(.in(layer_0[663]), .out(far_1_1791_0[0]));    relay_conn far_1_1791_0_b(.in(layer_0[542]), .out(far_1_1791_0[1]));
    wire [1:0] far_1_1791_1;    relay_conn far_1_1791_1_a(.in(far_1_1791_0[0]), .out(far_1_1791_1[0]));    relay_conn far_1_1791_1_b(.in(far_1_1791_0[1]), .out(far_1_1791_1[1]));
    wire [1:0] far_1_1791_2;    relay_conn far_1_1791_2_a(.in(far_1_1791_1[0]), .out(far_1_1791_2[0]));    relay_conn far_1_1791_2_b(.in(far_1_1791_1[1]), .out(far_1_1791_2[1]));
    assign layer_1[771] = ~far_1_1791_2[0]; 
    assign layer_1[772] = layer_0[119]; 
    wire [1:0] far_1_1793_0;    relay_conn far_1_1793_0_a(.in(layer_0[681]), .out(far_1_1793_0[0]));    relay_conn far_1_1793_0_b(.in(layer_0[743]), .out(far_1_1793_0[1]));
    assign layer_1[773] = ~(far_1_1793_0[0] | far_1_1793_0[1]); 
    wire [1:0] far_1_1794_0;    relay_conn far_1_1794_0_a(.in(layer_0[560]), .out(far_1_1794_0[0]));    relay_conn far_1_1794_0_b(.in(layer_0[629]), .out(far_1_1794_0[1]));
    wire [1:0] far_1_1794_1;    relay_conn far_1_1794_1_a(.in(far_1_1794_0[0]), .out(far_1_1794_1[0]));    relay_conn far_1_1794_1_b(.in(far_1_1794_0[1]), .out(far_1_1794_1[1]));
    assign layer_1[774] = far_1_1794_1[1]; 
    wire [1:0] far_1_1795_0;    relay_conn far_1_1795_0_a(.in(layer_0[305]), .out(far_1_1795_0[0]));    relay_conn far_1_1795_0_b(.in(layer_0[419]), .out(far_1_1795_0[1]));
    wire [1:0] far_1_1795_1;    relay_conn far_1_1795_1_a(.in(far_1_1795_0[0]), .out(far_1_1795_1[0]));    relay_conn far_1_1795_1_b(.in(far_1_1795_0[1]), .out(far_1_1795_1[1]));
    wire [1:0] far_1_1795_2;    relay_conn far_1_1795_2_a(.in(far_1_1795_1[0]), .out(far_1_1795_2[0]));    relay_conn far_1_1795_2_b(.in(far_1_1795_1[1]), .out(far_1_1795_2[1]));
    assign layer_1[775] = far_1_1795_2[0] & far_1_1795_2[1]; 
    assign layer_1[776] = layer_0[550] & ~layer_0[557]; 
    wire [1:0] far_1_1797_0;    relay_conn far_1_1797_0_a(.in(layer_0[696]), .out(far_1_1797_0[0]));    relay_conn far_1_1797_0_b(.in(layer_0[786]), .out(far_1_1797_0[1]));
    wire [1:0] far_1_1797_1;    relay_conn far_1_1797_1_a(.in(far_1_1797_0[0]), .out(far_1_1797_1[0]));    relay_conn far_1_1797_1_b(.in(far_1_1797_0[1]), .out(far_1_1797_1[1]));
    assign layer_1[777] = ~(far_1_1797_1[0] & far_1_1797_1[1]); 
    assign layer_1[778] = layer_0[379] | layer_0[404]; 
    assign layer_1[779] = ~layer_0[290] | (layer_0[313] & layer_0[290]); 
    assign layer_1[780] = ~layer_0[824] | (layer_0[855] & layer_0[824]); 
    wire [1:0] far_1_1801_0;    relay_conn far_1_1801_0_a(.in(layer_0[512]), .out(far_1_1801_0[0]));    relay_conn far_1_1801_0_b(.in(layer_0[580]), .out(far_1_1801_0[1]));
    wire [1:0] far_1_1801_1;    relay_conn far_1_1801_1_a(.in(far_1_1801_0[0]), .out(far_1_1801_1[0]));    relay_conn far_1_1801_1_b(.in(far_1_1801_0[1]), .out(far_1_1801_1[1]));
    assign layer_1[781] = far_1_1801_1[0]; 
    assign layer_1[782] = layer_0[676]; 
    wire [1:0] far_1_1803_0;    relay_conn far_1_1803_0_a(.in(layer_0[1002]), .out(far_1_1803_0[0]));    relay_conn far_1_1803_0_b(.in(layer_0[927]), .out(far_1_1803_0[1]));
    wire [1:0] far_1_1803_1;    relay_conn far_1_1803_1_a(.in(far_1_1803_0[0]), .out(far_1_1803_1[0]));    relay_conn far_1_1803_1_b(.in(far_1_1803_0[1]), .out(far_1_1803_1[1]));
    assign layer_1[783] = ~far_1_1803_1[1]; 
    wire [1:0] far_1_1804_0;    relay_conn far_1_1804_0_a(.in(layer_0[563]), .out(far_1_1804_0[0]));    relay_conn far_1_1804_0_b(.in(layer_0[504]), .out(far_1_1804_0[1]));
    assign layer_1[784] = far_1_1804_0[1]; 
    wire [1:0] far_1_1805_0;    relay_conn far_1_1805_0_a(.in(layer_0[81]), .out(far_1_1805_0[0]));    relay_conn far_1_1805_0_b(.in(layer_0[117]), .out(far_1_1805_0[1]));
    assign layer_1[785] = far_1_1805_0[1]; 
    wire [1:0] far_1_1806_0;    relay_conn far_1_1806_0_a(.in(layer_0[65]), .out(far_1_1806_0[0]));    relay_conn far_1_1806_0_b(.in(layer_0[107]), .out(far_1_1806_0[1]));
    assign layer_1[786] = ~far_1_1806_0[0] | (far_1_1806_0[0] & far_1_1806_0[1]); 
    wire [1:0] far_1_1807_0;    relay_conn far_1_1807_0_a(.in(layer_0[348]), .out(far_1_1807_0[0]));    relay_conn far_1_1807_0_b(.in(layer_0[476]), .out(far_1_1807_0[1]));
    wire [1:0] far_1_1807_1;    relay_conn far_1_1807_1_a(.in(far_1_1807_0[0]), .out(far_1_1807_1[0]));    relay_conn far_1_1807_1_b(.in(far_1_1807_0[1]), .out(far_1_1807_1[1]));
    wire [1:0] far_1_1807_2;    relay_conn far_1_1807_2_a(.in(far_1_1807_1[0]), .out(far_1_1807_2[0]));    relay_conn far_1_1807_2_b(.in(far_1_1807_1[1]), .out(far_1_1807_2[1]));
    wire [1:0] far_1_1807_3;    relay_conn far_1_1807_3_a(.in(far_1_1807_2[0]), .out(far_1_1807_3[0]));    relay_conn far_1_1807_3_b(.in(far_1_1807_2[1]), .out(far_1_1807_3[1]));
    assign layer_1[787] = ~far_1_1807_3[0] | (far_1_1807_3[0] & far_1_1807_3[1]); 
    assign layer_1[788] = ~layer_0[714] | (layer_0[714] & layer_0[732]); 
    wire [1:0] far_1_1809_0;    relay_conn far_1_1809_0_a(.in(layer_0[789]), .out(far_1_1809_0[0]));    relay_conn far_1_1809_0_b(.in(layer_0[861]), .out(far_1_1809_0[1]));
    wire [1:0] far_1_1809_1;    relay_conn far_1_1809_1_a(.in(far_1_1809_0[0]), .out(far_1_1809_1[0]));    relay_conn far_1_1809_1_b(.in(far_1_1809_0[1]), .out(far_1_1809_1[1]));
    assign layer_1[789] = ~(far_1_1809_1[0] & far_1_1809_1[1]); 
    assign layer_1[790] = ~layer_0[731]; 
    assign layer_1[791] = ~layer_0[750] | (layer_0[750] & layer_0[781]); 
    wire [1:0] far_1_1812_0;    relay_conn far_1_1812_0_a(.in(layer_0[354]), .out(far_1_1812_0[0]));    relay_conn far_1_1812_0_b(.in(layer_0[230]), .out(far_1_1812_0[1]));
    wire [1:0] far_1_1812_1;    relay_conn far_1_1812_1_a(.in(far_1_1812_0[0]), .out(far_1_1812_1[0]));    relay_conn far_1_1812_1_b(.in(far_1_1812_0[1]), .out(far_1_1812_1[1]));
    wire [1:0] far_1_1812_2;    relay_conn far_1_1812_2_a(.in(far_1_1812_1[0]), .out(far_1_1812_2[0]));    relay_conn far_1_1812_2_b(.in(far_1_1812_1[1]), .out(far_1_1812_2[1]));
    assign layer_1[792] = far_1_1812_2[0] & far_1_1812_2[1]; 
    assign layer_1[793] = ~layer_0[106]; 
    wire [1:0] far_1_1814_0;    relay_conn far_1_1814_0_a(.in(layer_0[367]), .out(far_1_1814_0[0]));    relay_conn far_1_1814_0_b(.in(layer_0[289]), .out(far_1_1814_0[1]));
    wire [1:0] far_1_1814_1;    relay_conn far_1_1814_1_a(.in(far_1_1814_0[0]), .out(far_1_1814_1[0]));    relay_conn far_1_1814_1_b(.in(far_1_1814_0[1]), .out(far_1_1814_1[1]));
    assign layer_1[794] = ~far_1_1814_1[1] | (far_1_1814_1[0] & far_1_1814_1[1]); 
    assign layer_1[795] = ~layer_0[265] | (layer_0[265] & layer_0[251]); 
    assign layer_1[796] = ~layer_0[93]; 
    wire [1:0] far_1_1817_0;    relay_conn far_1_1817_0_a(.in(layer_0[530]), .out(far_1_1817_0[0]));    relay_conn far_1_1817_0_b(.in(layer_0[656]), .out(far_1_1817_0[1]));
    wire [1:0] far_1_1817_1;    relay_conn far_1_1817_1_a(.in(far_1_1817_0[0]), .out(far_1_1817_1[0]));    relay_conn far_1_1817_1_b(.in(far_1_1817_0[1]), .out(far_1_1817_1[1]));
    wire [1:0] far_1_1817_2;    relay_conn far_1_1817_2_a(.in(far_1_1817_1[0]), .out(far_1_1817_2[0]));    relay_conn far_1_1817_2_b(.in(far_1_1817_1[1]), .out(far_1_1817_2[1]));
    assign layer_1[797] = far_1_1817_2[0] | far_1_1817_2[1]; 
    wire [1:0] far_1_1818_0;    relay_conn far_1_1818_0_a(.in(layer_0[484]), .out(far_1_1818_0[0]));    relay_conn far_1_1818_0_b(.in(layer_0[561]), .out(far_1_1818_0[1]));
    wire [1:0] far_1_1818_1;    relay_conn far_1_1818_1_a(.in(far_1_1818_0[0]), .out(far_1_1818_1[0]));    relay_conn far_1_1818_1_b(.in(far_1_1818_0[1]), .out(far_1_1818_1[1]));
    assign layer_1[798] = far_1_1818_1[0] & ~far_1_1818_1[1]; 
    wire [1:0] far_1_1819_0;    relay_conn far_1_1819_0_a(.in(layer_0[443]), .out(far_1_1819_0[0]));    relay_conn far_1_1819_0_b(.in(layer_0[562]), .out(far_1_1819_0[1]));
    wire [1:0] far_1_1819_1;    relay_conn far_1_1819_1_a(.in(far_1_1819_0[0]), .out(far_1_1819_1[0]));    relay_conn far_1_1819_1_b(.in(far_1_1819_0[1]), .out(far_1_1819_1[1]));
    wire [1:0] far_1_1819_2;    relay_conn far_1_1819_2_a(.in(far_1_1819_1[0]), .out(far_1_1819_2[0]));    relay_conn far_1_1819_2_b(.in(far_1_1819_1[1]), .out(far_1_1819_2[1]));
    assign layer_1[799] = ~(far_1_1819_2[0] & far_1_1819_2[1]); 
    wire [1:0] far_1_1820_0;    relay_conn far_1_1820_0_a(.in(layer_0[579]), .out(far_1_1820_0[0]));    relay_conn far_1_1820_0_b(.in(layer_0[530]), .out(far_1_1820_0[1]));
    assign layer_1[800] = far_1_1820_0[0]; 
    wire [1:0] far_1_1821_0;    relay_conn far_1_1821_0_a(.in(layer_0[852]), .out(far_1_1821_0[0]));    relay_conn far_1_1821_0_b(.in(layer_0[748]), .out(far_1_1821_0[1]));
    wire [1:0] far_1_1821_1;    relay_conn far_1_1821_1_a(.in(far_1_1821_0[0]), .out(far_1_1821_1[0]));    relay_conn far_1_1821_1_b(.in(far_1_1821_0[1]), .out(far_1_1821_1[1]));
    wire [1:0] far_1_1821_2;    relay_conn far_1_1821_2_a(.in(far_1_1821_1[0]), .out(far_1_1821_2[0]));    relay_conn far_1_1821_2_b(.in(far_1_1821_1[1]), .out(far_1_1821_2[1]));
    assign layer_1[801] = far_1_1821_2[0]; 
    assign layer_1[802] = layer_0[330] | layer_0[312]; 
    wire [1:0] far_1_1823_0;    relay_conn far_1_1823_0_a(.in(layer_0[471]), .out(far_1_1823_0[0]));    relay_conn far_1_1823_0_b(.in(layer_0[380]), .out(far_1_1823_0[1]));
    wire [1:0] far_1_1823_1;    relay_conn far_1_1823_1_a(.in(far_1_1823_0[0]), .out(far_1_1823_1[0]));    relay_conn far_1_1823_1_b(.in(far_1_1823_0[1]), .out(far_1_1823_1[1]));
    assign layer_1[803] = far_1_1823_1[0] ^ far_1_1823_1[1]; 
    wire [1:0] far_1_1824_0;    relay_conn far_1_1824_0_a(.in(layer_0[172]), .out(far_1_1824_0[0]));    relay_conn far_1_1824_0_b(.in(layer_0[83]), .out(far_1_1824_0[1]));
    wire [1:0] far_1_1824_1;    relay_conn far_1_1824_1_a(.in(far_1_1824_0[0]), .out(far_1_1824_1[0]));    relay_conn far_1_1824_1_b(.in(far_1_1824_0[1]), .out(far_1_1824_1[1]));
    assign layer_1[804] = far_1_1824_1[1] & ~far_1_1824_1[0]; 
    assign layer_1[805] = ~(layer_0[99] | layer_0[119]); 
    wire [1:0] far_1_1826_0;    relay_conn far_1_1826_0_a(.in(layer_0[478]), .out(far_1_1826_0[0]));    relay_conn far_1_1826_0_b(.in(layer_0[562]), .out(far_1_1826_0[1]));
    wire [1:0] far_1_1826_1;    relay_conn far_1_1826_1_a(.in(far_1_1826_0[0]), .out(far_1_1826_1[0]));    relay_conn far_1_1826_1_b(.in(far_1_1826_0[1]), .out(far_1_1826_1[1]));
    assign layer_1[806] = ~far_1_1826_1[0]; 
    wire [1:0] far_1_1827_0;    relay_conn far_1_1827_0_a(.in(layer_0[289]), .out(far_1_1827_0[0]));    relay_conn far_1_1827_0_b(.in(layer_0[397]), .out(far_1_1827_0[1]));
    wire [1:0] far_1_1827_1;    relay_conn far_1_1827_1_a(.in(far_1_1827_0[0]), .out(far_1_1827_1[0]));    relay_conn far_1_1827_1_b(.in(far_1_1827_0[1]), .out(far_1_1827_1[1]));
    wire [1:0] far_1_1827_2;    relay_conn far_1_1827_2_a(.in(far_1_1827_1[0]), .out(far_1_1827_2[0]));    relay_conn far_1_1827_2_b(.in(far_1_1827_1[1]), .out(far_1_1827_2[1]));
    assign layer_1[807] = ~(far_1_1827_2[0] ^ far_1_1827_2[1]); 
    wire [1:0] far_1_1828_0;    relay_conn far_1_1828_0_a(.in(layer_0[849]), .out(far_1_1828_0[0]));    relay_conn far_1_1828_0_b(.in(layer_0[930]), .out(far_1_1828_0[1]));
    wire [1:0] far_1_1828_1;    relay_conn far_1_1828_1_a(.in(far_1_1828_0[0]), .out(far_1_1828_1[0]));    relay_conn far_1_1828_1_b(.in(far_1_1828_0[1]), .out(far_1_1828_1[1]));
    assign layer_1[808] = far_1_1828_1[0] & ~far_1_1828_1[1]; 
    wire [1:0] far_1_1829_0;    relay_conn far_1_1829_0_a(.in(layer_0[562]), .out(far_1_1829_0[0]));    relay_conn far_1_1829_0_b(.in(layer_0[685]), .out(far_1_1829_0[1]));
    wire [1:0] far_1_1829_1;    relay_conn far_1_1829_1_a(.in(far_1_1829_0[0]), .out(far_1_1829_1[0]));    relay_conn far_1_1829_1_b(.in(far_1_1829_0[1]), .out(far_1_1829_1[1]));
    wire [1:0] far_1_1829_2;    relay_conn far_1_1829_2_a(.in(far_1_1829_1[0]), .out(far_1_1829_2[0]));    relay_conn far_1_1829_2_b(.in(far_1_1829_1[1]), .out(far_1_1829_2[1]));
    assign layer_1[809] = ~far_1_1829_2[1]; 
    assign layer_1[810] = ~(layer_0[710] ^ layer_0[732]); 
    assign layer_1[811] = layer_0[21] & layer_0[1]; 
    assign layer_1[812] = ~layer_0[51] | (layer_0[51] & layer_0[21]); 
    wire [1:0] far_1_1833_0;    relay_conn far_1_1833_0_a(.in(layer_0[327]), .out(far_1_1833_0[0]));    relay_conn far_1_1833_0_b(.in(layer_0[240]), .out(far_1_1833_0[1]));
    wire [1:0] far_1_1833_1;    relay_conn far_1_1833_1_a(.in(far_1_1833_0[0]), .out(far_1_1833_1[0]));    relay_conn far_1_1833_1_b(.in(far_1_1833_0[1]), .out(far_1_1833_1[1]));
    assign layer_1[813] = far_1_1833_1[1] & ~far_1_1833_1[0]; 
    wire [1:0] far_1_1834_0;    relay_conn far_1_1834_0_a(.in(layer_0[354]), .out(far_1_1834_0[0]));    relay_conn far_1_1834_0_b(.in(layer_0[318]), .out(far_1_1834_0[1]));
    assign layer_1[814] = far_1_1834_0[1] & ~far_1_1834_0[0]; 
    wire [1:0] far_1_1835_0;    relay_conn far_1_1835_0_a(.in(layer_0[610]), .out(far_1_1835_0[0]));    relay_conn far_1_1835_0_b(.in(layer_0[565]), .out(far_1_1835_0[1]));
    assign layer_1[815] = far_1_1835_0[1] & ~far_1_1835_0[0]; 
    wire [1:0] far_1_1836_0;    relay_conn far_1_1836_0_a(.in(layer_0[772]), .out(far_1_1836_0[0]));    relay_conn far_1_1836_0_b(.in(layer_0[655]), .out(far_1_1836_0[1]));
    wire [1:0] far_1_1836_1;    relay_conn far_1_1836_1_a(.in(far_1_1836_0[0]), .out(far_1_1836_1[0]));    relay_conn far_1_1836_1_b(.in(far_1_1836_0[1]), .out(far_1_1836_1[1]));
    wire [1:0] far_1_1836_2;    relay_conn far_1_1836_2_a(.in(far_1_1836_1[0]), .out(far_1_1836_2[0]));    relay_conn far_1_1836_2_b(.in(far_1_1836_1[1]), .out(far_1_1836_2[1]));
    assign layer_1[816] = far_1_1836_2[1] & ~far_1_1836_2[0]; 
    wire [1:0] far_1_1837_0;    relay_conn far_1_1837_0_a(.in(layer_0[639]), .out(far_1_1837_0[0]));    relay_conn far_1_1837_0_b(.in(layer_0[731]), .out(far_1_1837_0[1]));
    wire [1:0] far_1_1837_1;    relay_conn far_1_1837_1_a(.in(far_1_1837_0[0]), .out(far_1_1837_1[0]));    relay_conn far_1_1837_1_b(.in(far_1_1837_0[1]), .out(far_1_1837_1[1]));
    assign layer_1[817] = far_1_1837_1[1]; 
    wire [1:0] far_1_1838_0;    relay_conn far_1_1838_0_a(.in(layer_0[65]), .out(far_1_1838_0[0]));    relay_conn far_1_1838_0_b(.in(layer_0[128]), .out(far_1_1838_0[1]));
    assign layer_1[818] = ~far_1_1838_0[0]; 
    wire [1:0] far_1_1839_0;    relay_conn far_1_1839_0_a(.in(layer_0[1019]), .out(far_1_1839_0[0]));    relay_conn far_1_1839_0_b(.in(layer_0[954]), .out(far_1_1839_0[1]));
    wire [1:0] far_1_1839_1;    relay_conn far_1_1839_1_a(.in(far_1_1839_0[0]), .out(far_1_1839_1[0]));    relay_conn far_1_1839_1_b(.in(far_1_1839_0[1]), .out(far_1_1839_1[1]));
    assign layer_1[819] = far_1_1839_1[1]; 
    wire [1:0] far_1_1840_0;    relay_conn far_1_1840_0_a(.in(layer_0[512]), .out(far_1_1840_0[0]));    relay_conn far_1_1840_0_b(.in(layer_0[638]), .out(far_1_1840_0[1]));
    wire [1:0] far_1_1840_1;    relay_conn far_1_1840_1_a(.in(far_1_1840_0[0]), .out(far_1_1840_1[0]));    relay_conn far_1_1840_1_b(.in(far_1_1840_0[1]), .out(far_1_1840_1[1]));
    wire [1:0] far_1_1840_2;    relay_conn far_1_1840_2_a(.in(far_1_1840_1[0]), .out(far_1_1840_2[0]));    relay_conn far_1_1840_2_b(.in(far_1_1840_1[1]), .out(far_1_1840_2[1]));
    assign layer_1[820] = far_1_1840_2[0] & ~far_1_1840_2[1]; 
    assign layer_1[821] = ~layer_0[973] | (layer_0[973] & layer_0[967]); 
    wire [1:0] far_1_1842_0;    relay_conn far_1_1842_0_a(.in(layer_0[223]), .out(far_1_1842_0[0]));    relay_conn far_1_1842_0_b(.in(layer_0[124]), .out(far_1_1842_0[1]));
    wire [1:0] far_1_1842_1;    relay_conn far_1_1842_1_a(.in(far_1_1842_0[0]), .out(far_1_1842_1[0]));    relay_conn far_1_1842_1_b(.in(far_1_1842_0[1]), .out(far_1_1842_1[1]));
    wire [1:0] far_1_1842_2;    relay_conn far_1_1842_2_a(.in(far_1_1842_1[0]), .out(far_1_1842_2[0]));    relay_conn far_1_1842_2_b(.in(far_1_1842_1[1]), .out(far_1_1842_2[1]));
    assign layer_1[822] = far_1_1842_2[0] | far_1_1842_2[1]; 
    assign layer_1[823] = ~layer_0[218] | (layer_0[218] & layer_0[231]); 
    assign layer_1[824] = ~layer_0[852]; 
    wire [1:0] far_1_1845_0;    relay_conn far_1_1845_0_a(.in(layer_0[62]), .out(far_1_1845_0[0]));    relay_conn far_1_1845_0_b(.in(layer_0[185]), .out(far_1_1845_0[1]));
    wire [1:0] far_1_1845_1;    relay_conn far_1_1845_1_a(.in(far_1_1845_0[0]), .out(far_1_1845_1[0]));    relay_conn far_1_1845_1_b(.in(far_1_1845_0[1]), .out(far_1_1845_1[1]));
    wire [1:0] far_1_1845_2;    relay_conn far_1_1845_2_a(.in(far_1_1845_1[0]), .out(far_1_1845_2[0]));    relay_conn far_1_1845_2_b(.in(far_1_1845_1[1]), .out(far_1_1845_2[1]));
    assign layer_1[825] = far_1_1845_2[0]; 
    wire [1:0] far_1_1846_0;    relay_conn far_1_1846_0_a(.in(layer_0[1019]), .out(far_1_1846_0[0]));    relay_conn far_1_1846_0_b(.in(layer_0[916]), .out(far_1_1846_0[1]));
    wire [1:0] far_1_1846_1;    relay_conn far_1_1846_1_a(.in(far_1_1846_0[0]), .out(far_1_1846_1[0]));    relay_conn far_1_1846_1_b(.in(far_1_1846_0[1]), .out(far_1_1846_1[1]));
    wire [1:0] far_1_1846_2;    relay_conn far_1_1846_2_a(.in(far_1_1846_1[0]), .out(far_1_1846_2[0]));    relay_conn far_1_1846_2_b(.in(far_1_1846_1[1]), .out(far_1_1846_2[1]));
    assign layer_1[826] = far_1_1846_2[0] & ~far_1_1846_2[1]; 
    assign layer_1[827] = layer_0[768] | layer_0[777]; 
    assign layer_1[828] = layer_0[915]; 
    wire [1:0] far_1_1849_0;    relay_conn far_1_1849_0_a(.in(layer_0[906]), .out(far_1_1849_0[0]));    relay_conn far_1_1849_0_b(.in(layer_0[837]), .out(far_1_1849_0[1]));
    wire [1:0] far_1_1849_1;    relay_conn far_1_1849_1_a(.in(far_1_1849_0[0]), .out(far_1_1849_1[0]));    relay_conn far_1_1849_1_b(.in(far_1_1849_0[1]), .out(far_1_1849_1[1]));
    assign layer_1[829] = ~far_1_1849_1[1]; 
    wire [1:0] far_1_1850_0;    relay_conn far_1_1850_0_a(.in(layer_0[604]), .out(far_1_1850_0[0]));    relay_conn far_1_1850_0_b(.in(layer_0[481]), .out(far_1_1850_0[1]));
    wire [1:0] far_1_1850_1;    relay_conn far_1_1850_1_a(.in(far_1_1850_0[0]), .out(far_1_1850_1[0]));    relay_conn far_1_1850_1_b(.in(far_1_1850_0[1]), .out(far_1_1850_1[1]));
    wire [1:0] far_1_1850_2;    relay_conn far_1_1850_2_a(.in(far_1_1850_1[0]), .out(far_1_1850_2[0]));    relay_conn far_1_1850_2_b(.in(far_1_1850_1[1]), .out(far_1_1850_2[1]));
    assign layer_1[830] = ~far_1_1850_2[0] | (far_1_1850_2[0] & far_1_1850_2[1]); 
    wire [1:0] far_1_1851_0;    relay_conn far_1_1851_0_a(.in(layer_0[329]), .out(far_1_1851_0[0]));    relay_conn far_1_1851_0_b(.in(layer_0[372]), .out(far_1_1851_0[1]));
    assign layer_1[831] = ~far_1_1851_0[0]; 
    wire [1:0] far_1_1852_0;    relay_conn far_1_1852_0_a(.in(layer_0[400]), .out(far_1_1852_0[0]));    relay_conn far_1_1852_0_b(.in(layer_0[444]), .out(far_1_1852_0[1]));
    assign layer_1[832] = ~far_1_1852_0[1] | (far_1_1852_0[0] & far_1_1852_0[1]); 
    wire [1:0] far_1_1853_0;    relay_conn far_1_1853_0_a(.in(layer_0[118]), .out(far_1_1853_0[0]));    relay_conn far_1_1853_0_b(.in(layer_0[37]), .out(far_1_1853_0[1]));
    wire [1:0] far_1_1853_1;    relay_conn far_1_1853_1_a(.in(far_1_1853_0[0]), .out(far_1_1853_1[0]));    relay_conn far_1_1853_1_b(.in(far_1_1853_0[1]), .out(far_1_1853_1[1]));
    assign layer_1[833] = ~far_1_1853_1[1] | (far_1_1853_1[0] & far_1_1853_1[1]); 
    wire [1:0] far_1_1854_0;    relay_conn far_1_1854_0_a(.in(layer_0[939]), .out(far_1_1854_0[0]));    relay_conn far_1_1854_0_b(.in(layer_0[859]), .out(far_1_1854_0[1]));
    wire [1:0] far_1_1854_1;    relay_conn far_1_1854_1_a(.in(far_1_1854_0[0]), .out(far_1_1854_1[0]));    relay_conn far_1_1854_1_b(.in(far_1_1854_0[1]), .out(far_1_1854_1[1]));
    assign layer_1[834] = ~far_1_1854_1[0] | (far_1_1854_1[0] & far_1_1854_1[1]); 
    wire [1:0] far_1_1855_0;    relay_conn far_1_1855_0_a(.in(layer_0[284]), .out(far_1_1855_0[0]));    relay_conn far_1_1855_0_b(.in(layer_0[359]), .out(far_1_1855_0[1]));
    wire [1:0] far_1_1855_1;    relay_conn far_1_1855_1_a(.in(far_1_1855_0[0]), .out(far_1_1855_1[0]));    relay_conn far_1_1855_1_b(.in(far_1_1855_0[1]), .out(far_1_1855_1[1]));
    assign layer_1[835] = far_1_1855_1[1] & ~far_1_1855_1[0]; 
    wire [1:0] far_1_1856_0;    relay_conn far_1_1856_0_a(.in(layer_0[272]), .out(far_1_1856_0[0]));    relay_conn far_1_1856_0_b(.in(layer_0[170]), .out(far_1_1856_0[1]));
    wire [1:0] far_1_1856_1;    relay_conn far_1_1856_1_a(.in(far_1_1856_0[0]), .out(far_1_1856_1[0]));    relay_conn far_1_1856_1_b(.in(far_1_1856_0[1]), .out(far_1_1856_1[1]));
    wire [1:0] far_1_1856_2;    relay_conn far_1_1856_2_a(.in(far_1_1856_1[0]), .out(far_1_1856_2[0]));    relay_conn far_1_1856_2_b(.in(far_1_1856_1[1]), .out(far_1_1856_2[1]));
    assign layer_1[836] = far_1_1856_2[0] & far_1_1856_2[1]; 
    wire [1:0] far_1_1857_0;    relay_conn far_1_1857_0_a(.in(layer_0[395]), .out(far_1_1857_0[0]));    relay_conn far_1_1857_0_b(.in(layer_0[466]), .out(far_1_1857_0[1]));
    wire [1:0] far_1_1857_1;    relay_conn far_1_1857_1_a(.in(far_1_1857_0[0]), .out(far_1_1857_1[0]));    relay_conn far_1_1857_1_b(.in(far_1_1857_0[1]), .out(far_1_1857_1[1]));
    assign layer_1[837] = ~(far_1_1857_1[0] & far_1_1857_1[1]); 
    assign layer_1[838] = layer_0[283] | layer_0[313]; 
    wire [1:0] far_1_1859_0;    relay_conn far_1_1859_0_a(.in(layer_0[791]), .out(far_1_1859_0[0]));    relay_conn far_1_1859_0_b(.in(layer_0[705]), .out(far_1_1859_0[1]));
    wire [1:0] far_1_1859_1;    relay_conn far_1_1859_1_a(.in(far_1_1859_0[0]), .out(far_1_1859_1[0]));    relay_conn far_1_1859_1_b(.in(far_1_1859_0[1]), .out(far_1_1859_1[1]));
    assign layer_1[839] = ~(far_1_1859_1[0] & far_1_1859_1[1]); 
    assign layer_1[840] = layer_0[91] & ~layer_0[65]; 
    wire [1:0] far_1_1861_0;    relay_conn far_1_1861_0_a(.in(layer_0[318]), .out(far_1_1861_0[0]));    relay_conn far_1_1861_0_b(.in(layer_0[241]), .out(far_1_1861_0[1]));
    wire [1:0] far_1_1861_1;    relay_conn far_1_1861_1_a(.in(far_1_1861_0[0]), .out(far_1_1861_1[0]));    relay_conn far_1_1861_1_b(.in(far_1_1861_0[1]), .out(far_1_1861_1[1]));
    assign layer_1[841] = far_1_1861_1[0] & ~far_1_1861_1[1]; 
    wire [1:0] far_1_1862_0;    relay_conn far_1_1862_0_a(.in(layer_0[598]), .out(far_1_1862_0[0]));    relay_conn far_1_1862_0_b(.in(layer_0[721]), .out(far_1_1862_0[1]));
    wire [1:0] far_1_1862_1;    relay_conn far_1_1862_1_a(.in(far_1_1862_0[0]), .out(far_1_1862_1[0]));    relay_conn far_1_1862_1_b(.in(far_1_1862_0[1]), .out(far_1_1862_1[1]));
    wire [1:0] far_1_1862_2;    relay_conn far_1_1862_2_a(.in(far_1_1862_1[0]), .out(far_1_1862_2[0]));    relay_conn far_1_1862_2_b(.in(far_1_1862_1[1]), .out(far_1_1862_2[1]));
    assign layer_1[842] = ~far_1_1862_2[0] | (far_1_1862_2[0] & far_1_1862_2[1]); 
    wire [1:0] far_1_1863_0;    relay_conn far_1_1863_0_a(.in(layer_0[310]), .out(far_1_1863_0[0]));    relay_conn far_1_1863_0_b(.in(layer_0[392]), .out(far_1_1863_0[1]));
    wire [1:0] far_1_1863_1;    relay_conn far_1_1863_1_a(.in(far_1_1863_0[0]), .out(far_1_1863_1[0]));    relay_conn far_1_1863_1_b(.in(far_1_1863_0[1]), .out(far_1_1863_1[1]));
    assign layer_1[843] = far_1_1863_1[1] & ~far_1_1863_1[0]; 
    wire [1:0] far_1_1864_0;    relay_conn far_1_1864_0_a(.in(layer_0[459]), .out(far_1_1864_0[0]));    relay_conn far_1_1864_0_b(.in(layer_0[522]), .out(far_1_1864_0[1]));
    assign layer_1[844] = ~far_1_1864_0[1] | (far_1_1864_0[0] & far_1_1864_0[1]); 
    wire [1:0] far_1_1865_0;    relay_conn far_1_1865_0_a(.in(layer_0[862]), .out(far_1_1865_0[0]));    relay_conn far_1_1865_0_b(.in(layer_0[908]), .out(far_1_1865_0[1]));
    assign layer_1[845] = ~far_1_1865_0[1] | (far_1_1865_0[0] & far_1_1865_0[1]); 
    wire [1:0] far_1_1866_0;    relay_conn far_1_1866_0_a(.in(layer_0[349]), .out(far_1_1866_0[0]));    relay_conn far_1_1866_0_b(.in(layer_0[477]), .out(far_1_1866_0[1]));
    wire [1:0] far_1_1866_1;    relay_conn far_1_1866_1_a(.in(far_1_1866_0[0]), .out(far_1_1866_1[0]));    relay_conn far_1_1866_1_b(.in(far_1_1866_0[1]), .out(far_1_1866_1[1]));
    wire [1:0] far_1_1866_2;    relay_conn far_1_1866_2_a(.in(far_1_1866_1[0]), .out(far_1_1866_2[0]));    relay_conn far_1_1866_2_b(.in(far_1_1866_1[1]), .out(far_1_1866_2[1]));
    wire [1:0] far_1_1866_3;    relay_conn far_1_1866_3_a(.in(far_1_1866_2[0]), .out(far_1_1866_3[0]));    relay_conn far_1_1866_3_b(.in(far_1_1866_2[1]), .out(far_1_1866_3[1]));
    assign layer_1[846] = ~far_1_1866_3[1] | (far_1_1866_3[0] & far_1_1866_3[1]); 
    assign layer_1[847] = layer_0[194]; 
    assign layer_1[848] = layer_0[988]; 
    wire [1:0] far_1_1869_0;    relay_conn far_1_1869_0_a(.in(layer_0[597]), .out(far_1_1869_0[0]));    relay_conn far_1_1869_0_b(.in(layer_0[682]), .out(far_1_1869_0[1]));
    wire [1:0] far_1_1869_1;    relay_conn far_1_1869_1_a(.in(far_1_1869_0[0]), .out(far_1_1869_1[0]));    relay_conn far_1_1869_1_b(.in(far_1_1869_0[1]), .out(far_1_1869_1[1]));
    assign layer_1[849] = far_1_1869_1[0]; 
    wire [1:0] far_1_1870_0;    relay_conn far_1_1870_0_a(.in(layer_0[109]), .out(far_1_1870_0[0]));    relay_conn far_1_1870_0_b(.in(layer_0[232]), .out(far_1_1870_0[1]));
    wire [1:0] far_1_1870_1;    relay_conn far_1_1870_1_a(.in(far_1_1870_0[0]), .out(far_1_1870_1[0]));    relay_conn far_1_1870_1_b(.in(far_1_1870_0[1]), .out(far_1_1870_1[1]));
    wire [1:0] far_1_1870_2;    relay_conn far_1_1870_2_a(.in(far_1_1870_1[0]), .out(far_1_1870_2[0]));    relay_conn far_1_1870_2_b(.in(far_1_1870_1[1]), .out(far_1_1870_2[1]));
    assign layer_1[850] = far_1_1870_2[0] & far_1_1870_2[1]; 
    assign layer_1[851] = layer_0[604] ^ layer_0[607]; 
    assign layer_1[852] = ~(layer_0[328] | layer_0[307]); 
    wire [1:0] far_1_1873_0;    relay_conn far_1_1873_0_a(.in(layer_0[382]), .out(far_1_1873_0[0]));    relay_conn far_1_1873_0_b(.in(layer_0[258]), .out(far_1_1873_0[1]));
    wire [1:0] far_1_1873_1;    relay_conn far_1_1873_1_a(.in(far_1_1873_0[0]), .out(far_1_1873_1[0]));    relay_conn far_1_1873_1_b(.in(far_1_1873_0[1]), .out(far_1_1873_1[1]));
    wire [1:0] far_1_1873_2;    relay_conn far_1_1873_2_a(.in(far_1_1873_1[0]), .out(far_1_1873_2[0]));    relay_conn far_1_1873_2_b(.in(far_1_1873_1[1]), .out(far_1_1873_2[1]));
    assign layer_1[853] = ~far_1_1873_2[0]; 
    wire [1:0] far_1_1874_0;    relay_conn far_1_1874_0_a(.in(layer_0[313]), .out(far_1_1874_0[0]));    relay_conn far_1_1874_0_b(.in(layer_0[242]), .out(far_1_1874_0[1]));
    wire [1:0] far_1_1874_1;    relay_conn far_1_1874_1_a(.in(far_1_1874_0[0]), .out(far_1_1874_1[0]));    relay_conn far_1_1874_1_b(.in(far_1_1874_0[1]), .out(far_1_1874_1[1]));
    assign layer_1[854] = far_1_1874_1[0]; 
    wire [1:0] far_1_1875_0;    relay_conn far_1_1875_0_a(.in(layer_0[86]), .out(far_1_1875_0[0]));    relay_conn far_1_1875_0_b(.in(layer_0[194]), .out(far_1_1875_0[1]));
    wire [1:0] far_1_1875_1;    relay_conn far_1_1875_1_a(.in(far_1_1875_0[0]), .out(far_1_1875_1[0]));    relay_conn far_1_1875_1_b(.in(far_1_1875_0[1]), .out(far_1_1875_1[1]));
    wire [1:0] far_1_1875_2;    relay_conn far_1_1875_2_a(.in(far_1_1875_1[0]), .out(far_1_1875_2[0]));    relay_conn far_1_1875_2_b(.in(far_1_1875_1[1]), .out(far_1_1875_2[1]));
    assign layer_1[855] = far_1_1875_2[1] & ~far_1_1875_2[0]; 
    wire [1:0] far_1_1876_0;    relay_conn far_1_1876_0_a(.in(layer_0[768]), .out(far_1_1876_0[0]));    relay_conn far_1_1876_0_b(.in(layer_0[701]), .out(far_1_1876_0[1]));
    wire [1:0] far_1_1876_1;    relay_conn far_1_1876_1_a(.in(far_1_1876_0[0]), .out(far_1_1876_1[0]));    relay_conn far_1_1876_1_b(.in(far_1_1876_0[1]), .out(far_1_1876_1[1]));
    assign layer_1[856] = far_1_1876_1[1] & ~far_1_1876_1[0]; 
    wire [1:0] far_1_1877_0;    relay_conn far_1_1877_0_a(.in(layer_0[777]), .out(far_1_1877_0[0]));    relay_conn far_1_1877_0_b(.in(layer_0[686]), .out(far_1_1877_0[1]));
    wire [1:0] far_1_1877_1;    relay_conn far_1_1877_1_a(.in(far_1_1877_0[0]), .out(far_1_1877_1[0]));    relay_conn far_1_1877_1_b(.in(far_1_1877_0[1]), .out(far_1_1877_1[1]));
    assign layer_1[857] = ~(far_1_1877_1[0] ^ far_1_1877_1[1]); 
    wire [1:0] far_1_1878_0;    relay_conn far_1_1878_0_a(.in(layer_0[361]), .out(far_1_1878_0[0]));    relay_conn far_1_1878_0_b(.in(layer_0[276]), .out(far_1_1878_0[1]));
    wire [1:0] far_1_1878_1;    relay_conn far_1_1878_1_a(.in(far_1_1878_0[0]), .out(far_1_1878_1[0]));    relay_conn far_1_1878_1_b(.in(far_1_1878_0[1]), .out(far_1_1878_1[1]));
    assign layer_1[858] = far_1_1878_1[1]; 
    assign layer_1[859] = ~(layer_0[832] & layer_0[810]); 
    wire [1:0] far_1_1880_0;    relay_conn far_1_1880_0_a(.in(layer_0[65]), .out(far_1_1880_0[0]));    relay_conn far_1_1880_0_b(.in(layer_0[123]), .out(far_1_1880_0[1]));
    assign layer_1[860] = ~far_1_1880_0[0] | (far_1_1880_0[0] & far_1_1880_0[1]); 
    wire [1:0] far_1_1881_0;    relay_conn far_1_1881_0_a(.in(layer_0[530]), .out(far_1_1881_0[0]));    relay_conn far_1_1881_0_b(.in(layer_0[442]), .out(far_1_1881_0[1]));
    wire [1:0] far_1_1881_1;    relay_conn far_1_1881_1_a(.in(far_1_1881_0[0]), .out(far_1_1881_1[0]));    relay_conn far_1_1881_1_b(.in(far_1_1881_0[1]), .out(far_1_1881_1[1]));
    assign layer_1[861] = ~(far_1_1881_1[0] ^ far_1_1881_1[1]); 
    wire [1:0] far_1_1882_0;    relay_conn far_1_1882_0_a(.in(layer_0[305]), .out(far_1_1882_0[0]));    relay_conn far_1_1882_0_b(.in(layer_0[354]), .out(far_1_1882_0[1]));
    assign layer_1[862] = ~far_1_1882_0[0] | (far_1_1882_0[0] & far_1_1882_0[1]); 
    wire [1:0] far_1_1883_0;    relay_conn far_1_1883_0_a(.in(layer_0[889]), .out(far_1_1883_0[0]));    relay_conn far_1_1883_0_b(.in(layer_0[826]), .out(far_1_1883_0[1]));
    assign layer_1[863] = far_1_1883_0[0] & far_1_1883_0[1]; 
    assign layer_1[864] = layer_0[444]; 
    assign layer_1[865] = layer_0[956] & ~layer_0[927]; 
    wire [1:0] far_1_1886_0;    relay_conn far_1_1886_0_a(.in(layer_0[702]), .out(far_1_1886_0[0]));    relay_conn far_1_1886_0_b(.in(layer_0[815]), .out(far_1_1886_0[1]));
    wire [1:0] far_1_1886_1;    relay_conn far_1_1886_1_a(.in(far_1_1886_0[0]), .out(far_1_1886_1[0]));    relay_conn far_1_1886_1_b(.in(far_1_1886_0[1]), .out(far_1_1886_1[1]));
    wire [1:0] far_1_1886_2;    relay_conn far_1_1886_2_a(.in(far_1_1886_1[0]), .out(far_1_1886_2[0]));    relay_conn far_1_1886_2_b(.in(far_1_1886_1[1]), .out(far_1_1886_2[1]));
    assign layer_1[866] = ~far_1_1886_2[0]; 
    assign layer_1[867] = ~(layer_0[362] | layer_0[385]); 
    wire [1:0] far_1_1888_0;    relay_conn far_1_1888_0_a(.in(layer_0[265]), .out(far_1_1888_0[0]));    relay_conn far_1_1888_0_b(.in(layer_0[377]), .out(far_1_1888_0[1]));
    wire [1:0] far_1_1888_1;    relay_conn far_1_1888_1_a(.in(far_1_1888_0[0]), .out(far_1_1888_1[0]));    relay_conn far_1_1888_1_b(.in(far_1_1888_0[1]), .out(far_1_1888_1[1]));
    wire [1:0] far_1_1888_2;    relay_conn far_1_1888_2_a(.in(far_1_1888_1[0]), .out(far_1_1888_2[0]));    relay_conn far_1_1888_2_b(.in(far_1_1888_1[1]), .out(far_1_1888_2[1]));
    assign layer_1[868] = far_1_1888_2[0] ^ far_1_1888_2[1]; 
    wire [1:0] far_1_1889_0;    relay_conn far_1_1889_0_a(.in(layer_0[443]), .out(far_1_1889_0[0]));    relay_conn far_1_1889_0_b(.in(layer_0[377]), .out(far_1_1889_0[1]));
    wire [1:0] far_1_1889_1;    relay_conn far_1_1889_1_a(.in(far_1_1889_0[0]), .out(far_1_1889_1[0]));    relay_conn far_1_1889_1_b(.in(far_1_1889_0[1]), .out(far_1_1889_1[1]));
    assign layer_1[869] = far_1_1889_1[0] ^ far_1_1889_1[1]; 
    wire [1:0] far_1_1890_0;    relay_conn far_1_1890_0_a(.in(layer_0[579]), .out(far_1_1890_0[0]));    relay_conn far_1_1890_0_b(.in(layer_0[676]), .out(far_1_1890_0[1]));
    wire [1:0] far_1_1890_1;    relay_conn far_1_1890_1_a(.in(far_1_1890_0[0]), .out(far_1_1890_1[0]));    relay_conn far_1_1890_1_b(.in(far_1_1890_0[1]), .out(far_1_1890_1[1]));
    wire [1:0] far_1_1890_2;    relay_conn far_1_1890_2_a(.in(far_1_1890_1[0]), .out(far_1_1890_2[0]));    relay_conn far_1_1890_2_b(.in(far_1_1890_1[1]), .out(far_1_1890_2[1]));
    assign layer_1[870] = far_1_1890_2[0]; 
    wire [1:0] far_1_1891_0;    relay_conn far_1_1891_0_a(.in(layer_0[344]), .out(far_1_1891_0[0]));    relay_conn far_1_1891_0_b(.in(layer_0[252]), .out(far_1_1891_0[1]));
    wire [1:0] far_1_1891_1;    relay_conn far_1_1891_1_a(.in(far_1_1891_0[0]), .out(far_1_1891_1[0]));    relay_conn far_1_1891_1_b(.in(far_1_1891_0[1]), .out(far_1_1891_1[1]));
    assign layer_1[871] = far_1_1891_1[1] & ~far_1_1891_1[0]; 
    wire [1:0] far_1_1892_0;    relay_conn far_1_1892_0_a(.in(layer_0[376]), .out(far_1_1892_0[0]));    relay_conn far_1_1892_0_b(.in(layer_0[484]), .out(far_1_1892_0[1]));
    wire [1:0] far_1_1892_1;    relay_conn far_1_1892_1_a(.in(far_1_1892_0[0]), .out(far_1_1892_1[0]));    relay_conn far_1_1892_1_b(.in(far_1_1892_0[1]), .out(far_1_1892_1[1]));
    wire [1:0] far_1_1892_2;    relay_conn far_1_1892_2_a(.in(far_1_1892_1[0]), .out(far_1_1892_2[0]));    relay_conn far_1_1892_2_b(.in(far_1_1892_1[1]), .out(far_1_1892_2[1]));
    assign layer_1[872] = far_1_1892_2[0]; 
    assign layer_1[873] = layer_0[694] & layer_0[702]; 
    assign layer_1[874] = layer_0[299] & layer_0[280]; 
    assign layer_1[875] = layer_0[893] & layer_0[884]; 
    assign layer_1[876] = layer_0[979] & ~layer_0[950]; 
    wire [1:0] far_1_1897_0;    relay_conn far_1_1897_0_a(.in(layer_0[330]), .out(far_1_1897_0[0]));    relay_conn far_1_1897_0_b(.in(layer_0[441]), .out(far_1_1897_0[1]));
    wire [1:0] far_1_1897_1;    relay_conn far_1_1897_1_a(.in(far_1_1897_0[0]), .out(far_1_1897_1[0]));    relay_conn far_1_1897_1_b(.in(far_1_1897_0[1]), .out(far_1_1897_1[1]));
    wire [1:0] far_1_1897_2;    relay_conn far_1_1897_2_a(.in(far_1_1897_1[0]), .out(far_1_1897_2[0]));    relay_conn far_1_1897_2_b(.in(far_1_1897_1[1]), .out(far_1_1897_2[1]));
    assign layer_1[877] = far_1_1897_2[0]; 
    wire [1:0] far_1_1898_0;    relay_conn far_1_1898_0_a(.in(layer_0[253]), .out(far_1_1898_0[0]));    relay_conn far_1_1898_0_b(.in(layer_0[178]), .out(far_1_1898_0[1]));
    wire [1:0] far_1_1898_1;    relay_conn far_1_1898_1_a(.in(far_1_1898_0[0]), .out(far_1_1898_1[0]));    relay_conn far_1_1898_1_b(.in(far_1_1898_0[1]), .out(far_1_1898_1[1]));
    assign layer_1[878] = ~far_1_1898_1[0]; 
    assign layer_1[879] = layer_0[577] & ~layer_0[599]; 
    wire [1:0] far_1_1900_0;    relay_conn far_1_1900_0_a(.in(layer_0[577]), .out(far_1_1900_0[0]));    relay_conn far_1_1900_0_b(.in(layer_0[544]), .out(far_1_1900_0[1]));
    assign layer_1[880] = ~far_1_1900_0[1] | (far_1_1900_0[0] & far_1_1900_0[1]); 
    assign layer_1[881] = layer_0[607] & ~layer_0[614]; 
    wire [1:0] far_1_1902_0;    relay_conn far_1_1902_0_a(.in(layer_0[726]), .out(far_1_1902_0[0]));    relay_conn far_1_1902_0_b(.in(layer_0[843]), .out(far_1_1902_0[1]));
    wire [1:0] far_1_1902_1;    relay_conn far_1_1902_1_a(.in(far_1_1902_0[0]), .out(far_1_1902_1[0]));    relay_conn far_1_1902_1_b(.in(far_1_1902_0[1]), .out(far_1_1902_1[1]));
    wire [1:0] far_1_1902_2;    relay_conn far_1_1902_2_a(.in(far_1_1902_1[0]), .out(far_1_1902_2[0]));    relay_conn far_1_1902_2_b(.in(far_1_1902_1[1]), .out(far_1_1902_2[1]));
    assign layer_1[882] = far_1_1902_2[0] & ~far_1_1902_2[1]; 
    wire [1:0] far_1_1903_0;    relay_conn far_1_1903_0_a(.in(layer_0[884]), .out(far_1_1903_0[0]));    relay_conn far_1_1903_0_b(.in(layer_0[1011]), .out(far_1_1903_0[1]));
    wire [1:0] far_1_1903_1;    relay_conn far_1_1903_1_a(.in(far_1_1903_0[0]), .out(far_1_1903_1[0]));    relay_conn far_1_1903_1_b(.in(far_1_1903_0[1]), .out(far_1_1903_1[1]));
    wire [1:0] far_1_1903_2;    relay_conn far_1_1903_2_a(.in(far_1_1903_1[0]), .out(far_1_1903_2[0]));    relay_conn far_1_1903_2_b(.in(far_1_1903_1[1]), .out(far_1_1903_2[1]));
    assign layer_1[883] = ~far_1_1903_2[1]; 
    assign layer_1[884] = ~(layer_0[612] | layer_0[607]); 
    wire [1:0] far_1_1905_0;    relay_conn far_1_1905_0_a(.in(layer_0[339]), .out(far_1_1905_0[0]));    relay_conn far_1_1905_0_b(.in(layer_0[392]), .out(far_1_1905_0[1]));
    assign layer_1[885] = ~far_1_1905_0[1]; 
    wire [1:0] far_1_1906_0;    relay_conn far_1_1906_0_a(.in(layer_0[157]), .out(far_1_1906_0[0]));    relay_conn far_1_1906_0_b(.in(layer_0[190]), .out(far_1_1906_0[1]));
    assign layer_1[886] = far_1_1906_0[0] | far_1_1906_0[1]; 
    wire [1:0] far_1_1907_0;    relay_conn far_1_1907_0_a(.in(layer_0[156]), .out(far_1_1907_0[0]));    relay_conn far_1_1907_0_b(.in(layer_0[123]), .out(far_1_1907_0[1]));
    assign layer_1[887] = far_1_1907_0[1] & ~far_1_1907_0[0]; 
    assign layer_1[888] = ~(layer_0[908] & layer_0[877]); 
    wire [1:0] far_1_1909_0;    relay_conn far_1_1909_0_a(.in(layer_0[356]), .out(far_1_1909_0[0]));    relay_conn far_1_1909_0_b(.in(layer_0[242]), .out(far_1_1909_0[1]));
    wire [1:0] far_1_1909_1;    relay_conn far_1_1909_1_a(.in(far_1_1909_0[0]), .out(far_1_1909_1[0]));    relay_conn far_1_1909_1_b(.in(far_1_1909_0[1]), .out(far_1_1909_1[1]));
    wire [1:0] far_1_1909_2;    relay_conn far_1_1909_2_a(.in(far_1_1909_1[0]), .out(far_1_1909_2[0]));    relay_conn far_1_1909_2_b(.in(far_1_1909_1[1]), .out(far_1_1909_2[1]));
    assign layer_1[889] = ~(far_1_1909_2[0] | far_1_1909_2[1]); 
    wire [1:0] far_1_1910_0;    relay_conn far_1_1910_0_a(.in(layer_0[702]), .out(far_1_1910_0[0]));    relay_conn far_1_1910_0_b(.in(layer_0[617]), .out(far_1_1910_0[1]));
    wire [1:0] far_1_1910_1;    relay_conn far_1_1910_1_a(.in(far_1_1910_0[0]), .out(far_1_1910_1[0]));    relay_conn far_1_1910_1_b(.in(far_1_1910_0[1]), .out(far_1_1910_1[1]));
    assign layer_1[890] = ~far_1_1910_1[0]; 
    wire [1:0] far_1_1911_0;    relay_conn far_1_1911_0_a(.in(layer_0[1006]), .out(far_1_1911_0[0]));    relay_conn far_1_1911_0_b(.in(layer_0[894]), .out(far_1_1911_0[1]));
    wire [1:0] far_1_1911_1;    relay_conn far_1_1911_1_a(.in(far_1_1911_0[0]), .out(far_1_1911_1[0]));    relay_conn far_1_1911_1_b(.in(far_1_1911_0[1]), .out(far_1_1911_1[1]));
    wire [1:0] far_1_1911_2;    relay_conn far_1_1911_2_a(.in(far_1_1911_1[0]), .out(far_1_1911_2[0]));    relay_conn far_1_1911_2_b(.in(far_1_1911_1[1]), .out(far_1_1911_2[1]));
    assign layer_1[891] = far_1_1911_2[0] & far_1_1911_2[1]; 
    wire [1:0] far_1_1912_0;    relay_conn far_1_1912_0_a(.in(layer_0[630]), .out(far_1_1912_0[0]));    relay_conn far_1_1912_0_b(.in(layer_0[554]), .out(far_1_1912_0[1]));
    wire [1:0] far_1_1912_1;    relay_conn far_1_1912_1_a(.in(far_1_1912_0[0]), .out(far_1_1912_1[0]));    relay_conn far_1_1912_1_b(.in(far_1_1912_0[1]), .out(far_1_1912_1[1]));
    assign layer_1[892] = far_1_1912_1[0] & far_1_1912_1[1]; 
    wire [1:0] far_1_1913_0;    relay_conn far_1_1913_0_a(.in(layer_0[970]), .out(far_1_1913_0[0]));    relay_conn far_1_1913_0_b(.in(layer_0[873]), .out(far_1_1913_0[1]));
    wire [1:0] far_1_1913_1;    relay_conn far_1_1913_1_a(.in(far_1_1913_0[0]), .out(far_1_1913_1[0]));    relay_conn far_1_1913_1_b(.in(far_1_1913_0[1]), .out(far_1_1913_1[1]));
    wire [1:0] far_1_1913_2;    relay_conn far_1_1913_2_a(.in(far_1_1913_1[0]), .out(far_1_1913_2[0]));    relay_conn far_1_1913_2_b(.in(far_1_1913_1[1]), .out(far_1_1913_2[1]));
    assign layer_1[893] = ~(far_1_1913_2[0] & far_1_1913_2[1]); 
    assign layer_1[894] = ~layer_0[100] | (layer_0[100] & layer_0[81]); 
    assign layer_1[895] = layer_0[984] & layer_0[997]; 
    wire [1:0] far_1_1916_0;    relay_conn far_1_1916_0_a(.in(layer_0[410]), .out(far_1_1916_0[0]));    relay_conn far_1_1916_0_b(.in(layer_0[506]), .out(far_1_1916_0[1]));
    wire [1:0] far_1_1916_1;    relay_conn far_1_1916_1_a(.in(far_1_1916_0[0]), .out(far_1_1916_1[0]));    relay_conn far_1_1916_1_b(.in(far_1_1916_0[1]), .out(far_1_1916_1[1]));
    wire [1:0] far_1_1916_2;    relay_conn far_1_1916_2_a(.in(far_1_1916_1[0]), .out(far_1_1916_2[0]));    relay_conn far_1_1916_2_b(.in(far_1_1916_1[1]), .out(far_1_1916_2[1]));
    assign layer_1[896] = ~far_1_1916_2[0]; 
    assign layer_1[897] = ~layer_0[503]; 
    wire [1:0] far_1_1918_0;    relay_conn far_1_1918_0_a(.in(layer_0[678]), .out(far_1_1918_0[0]));    relay_conn far_1_1918_0_b(.in(layer_0[607]), .out(far_1_1918_0[1]));
    wire [1:0] far_1_1918_1;    relay_conn far_1_1918_1_a(.in(far_1_1918_0[0]), .out(far_1_1918_1[0]));    relay_conn far_1_1918_1_b(.in(far_1_1918_0[1]), .out(far_1_1918_1[1]));
    assign layer_1[898] = far_1_1918_1[0] & ~far_1_1918_1[1]; 
    wire [1:0] far_1_1919_0;    relay_conn far_1_1919_0_a(.in(layer_0[367]), .out(far_1_1919_0[0]));    relay_conn far_1_1919_0_b(.in(layer_0[282]), .out(far_1_1919_0[1]));
    wire [1:0] far_1_1919_1;    relay_conn far_1_1919_1_a(.in(far_1_1919_0[0]), .out(far_1_1919_1[0]));    relay_conn far_1_1919_1_b(.in(far_1_1919_0[1]), .out(far_1_1919_1[1]));
    assign layer_1[899] = ~far_1_1919_1[0]; 
    assign layer_1[900] = ~layer_0[339]; 
    wire [1:0] far_1_1921_0;    relay_conn far_1_1921_0_a(.in(layer_0[66]), .out(far_1_1921_0[0]));    relay_conn far_1_1921_0_b(.in(layer_0[150]), .out(far_1_1921_0[1]));
    wire [1:0] far_1_1921_1;    relay_conn far_1_1921_1_a(.in(far_1_1921_0[0]), .out(far_1_1921_1[0]));    relay_conn far_1_1921_1_b(.in(far_1_1921_0[1]), .out(far_1_1921_1[1]));
    assign layer_1[901] = ~far_1_1921_1[0] | (far_1_1921_1[0] & far_1_1921_1[1]); 
    wire [1:0] far_1_1922_0;    relay_conn far_1_1922_0_a(.in(layer_0[777]), .out(far_1_1922_0[0]));    relay_conn far_1_1922_0_b(.in(layer_0[888]), .out(far_1_1922_0[1]));
    wire [1:0] far_1_1922_1;    relay_conn far_1_1922_1_a(.in(far_1_1922_0[0]), .out(far_1_1922_1[0]));    relay_conn far_1_1922_1_b(.in(far_1_1922_0[1]), .out(far_1_1922_1[1]));
    wire [1:0] far_1_1922_2;    relay_conn far_1_1922_2_a(.in(far_1_1922_1[0]), .out(far_1_1922_2[0]));    relay_conn far_1_1922_2_b(.in(far_1_1922_1[1]), .out(far_1_1922_2[1]));
    assign layer_1[902] = ~far_1_1922_2[1] | (far_1_1922_2[0] & far_1_1922_2[1]); 
    wire [1:0] far_1_1923_0;    relay_conn far_1_1923_0_a(.in(layer_0[195]), .out(far_1_1923_0[0]));    relay_conn far_1_1923_0_b(.in(layer_0[303]), .out(far_1_1923_0[1]));
    wire [1:0] far_1_1923_1;    relay_conn far_1_1923_1_a(.in(far_1_1923_0[0]), .out(far_1_1923_1[0]));    relay_conn far_1_1923_1_b(.in(far_1_1923_0[1]), .out(far_1_1923_1[1]));
    wire [1:0] far_1_1923_2;    relay_conn far_1_1923_2_a(.in(far_1_1923_1[0]), .out(far_1_1923_2[0]));    relay_conn far_1_1923_2_b(.in(far_1_1923_1[1]), .out(far_1_1923_2[1]));
    assign layer_1[903] = far_1_1923_2[0] & ~far_1_1923_2[1]; 
    assign layer_1[904] = ~layer_0[937]; 
    wire [1:0] far_1_1925_0;    relay_conn far_1_1925_0_a(.in(layer_0[480]), .out(far_1_1925_0[0]));    relay_conn far_1_1925_0_b(.in(layer_0[438]), .out(far_1_1925_0[1]));
    assign layer_1[905] = far_1_1925_0[0]; 
    wire [1:0] far_1_1926_0;    relay_conn far_1_1926_0_a(.in(layer_0[285]), .out(far_1_1926_0[0]));    relay_conn far_1_1926_0_b(.in(layer_0[381]), .out(far_1_1926_0[1]));
    wire [1:0] far_1_1926_1;    relay_conn far_1_1926_1_a(.in(far_1_1926_0[0]), .out(far_1_1926_1[0]));    relay_conn far_1_1926_1_b(.in(far_1_1926_0[1]), .out(far_1_1926_1[1]));
    wire [1:0] far_1_1926_2;    relay_conn far_1_1926_2_a(.in(far_1_1926_1[0]), .out(far_1_1926_2[0]));    relay_conn far_1_1926_2_b(.in(far_1_1926_1[1]), .out(far_1_1926_2[1]));
    assign layer_1[906] = ~far_1_1926_2[1]; 
    assign layer_1[907] = layer_0[152] | layer_0[172]; 
    wire [1:0] far_1_1928_0;    relay_conn far_1_1928_0_a(.in(layer_0[487]), .out(far_1_1928_0[0]));    relay_conn far_1_1928_0_b(.in(layer_0[400]), .out(far_1_1928_0[1]));
    wire [1:0] far_1_1928_1;    relay_conn far_1_1928_1_a(.in(far_1_1928_0[0]), .out(far_1_1928_1[0]));    relay_conn far_1_1928_1_b(.in(far_1_1928_0[1]), .out(far_1_1928_1[1]));
    assign layer_1[908] = far_1_1928_1[1]; 
    assign layer_1[909] = ~layer_0[985] | (layer_0[985] & layer_0[954]); 
    assign layer_1[910] = layer_0[849] | layer_0[874]; 
    wire [1:0] far_1_1931_0;    relay_conn far_1_1931_0_a(.in(layer_0[841]), .out(far_1_1931_0[0]));    relay_conn far_1_1931_0_b(.in(layer_0[891]), .out(far_1_1931_0[1]));
    assign layer_1[911] = far_1_1931_0[0] & far_1_1931_0[1]; 
    wire [1:0] far_1_1932_0;    relay_conn far_1_1932_0_a(.in(layer_0[946]), .out(far_1_1932_0[0]));    relay_conn far_1_1932_0_b(.in(layer_0[1002]), .out(far_1_1932_0[1]));
    assign layer_1[912] = far_1_1932_0[1] & ~far_1_1932_0[0]; 
    wire [1:0] far_1_1933_0;    relay_conn far_1_1933_0_a(.in(layer_0[251]), .out(far_1_1933_0[0]));    relay_conn far_1_1933_0_b(.in(layer_0[356]), .out(far_1_1933_0[1]));
    wire [1:0] far_1_1933_1;    relay_conn far_1_1933_1_a(.in(far_1_1933_0[0]), .out(far_1_1933_1[0]));    relay_conn far_1_1933_1_b(.in(far_1_1933_0[1]), .out(far_1_1933_1[1]));
    wire [1:0] far_1_1933_2;    relay_conn far_1_1933_2_a(.in(far_1_1933_1[0]), .out(far_1_1933_2[0]));    relay_conn far_1_1933_2_b(.in(far_1_1933_1[1]), .out(far_1_1933_2[1]));
    assign layer_1[913] = ~far_1_1933_2[0]; 
    wire [1:0] far_1_1934_0;    relay_conn far_1_1934_0_a(.in(layer_0[565]), .out(far_1_1934_0[0]));    relay_conn far_1_1934_0_b(.in(layer_0[509]), .out(far_1_1934_0[1]));
    assign layer_1[914] = ~(far_1_1934_0[0] ^ far_1_1934_0[1]); 
    wire [1:0] far_1_1935_0;    relay_conn far_1_1935_0_a(.in(layer_0[791]), .out(far_1_1935_0[0]));    relay_conn far_1_1935_0_b(.in(layer_0[886]), .out(far_1_1935_0[1]));
    wire [1:0] far_1_1935_1;    relay_conn far_1_1935_1_a(.in(far_1_1935_0[0]), .out(far_1_1935_1[0]));    relay_conn far_1_1935_1_b(.in(far_1_1935_0[1]), .out(far_1_1935_1[1]));
    assign layer_1[915] = ~far_1_1935_1[0]; 
    assign layer_1[916] = layer_0[697]; 
    wire [1:0] far_1_1937_0;    relay_conn far_1_1937_0_a(.in(layer_0[307]), .out(far_1_1937_0[0]));    relay_conn far_1_1937_0_b(.in(layer_0[407]), .out(far_1_1937_0[1]));
    wire [1:0] far_1_1937_1;    relay_conn far_1_1937_1_a(.in(far_1_1937_0[0]), .out(far_1_1937_1[0]));    relay_conn far_1_1937_1_b(.in(far_1_1937_0[1]), .out(far_1_1937_1[1]));
    wire [1:0] far_1_1937_2;    relay_conn far_1_1937_2_a(.in(far_1_1937_1[0]), .out(far_1_1937_2[0]));    relay_conn far_1_1937_2_b(.in(far_1_1937_1[1]), .out(far_1_1937_2[1]));
    assign layer_1[917] = ~far_1_1937_2[0]; 
    wire [1:0] far_1_1938_0;    relay_conn far_1_1938_0_a(.in(layer_0[293]), .out(far_1_1938_0[0]));    relay_conn far_1_1938_0_b(.in(layer_0[243]), .out(far_1_1938_0[1]));
    assign layer_1[918] = ~far_1_1938_0[1]; 
    assign layer_1[919] = ~(layer_0[485] | layer_0[497]); 
    wire [1:0] far_1_1940_0;    relay_conn far_1_1940_0_a(.in(layer_0[960]), .out(far_1_1940_0[0]));    relay_conn far_1_1940_0_b(.in(layer_0[854]), .out(far_1_1940_0[1]));
    wire [1:0] far_1_1940_1;    relay_conn far_1_1940_1_a(.in(far_1_1940_0[0]), .out(far_1_1940_1[0]));    relay_conn far_1_1940_1_b(.in(far_1_1940_0[1]), .out(far_1_1940_1[1]));
    wire [1:0] far_1_1940_2;    relay_conn far_1_1940_2_a(.in(far_1_1940_1[0]), .out(far_1_1940_2[0]));    relay_conn far_1_1940_2_b(.in(far_1_1940_1[1]), .out(far_1_1940_2[1]));
    assign layer_1[920] = far_1_1940_2[0] & ~far_1_1940_2[1]; 
    wire [1:0] far_1_1941_0;    relay_conn far_1_1941_0_a(.in(layer_0[1011]), .out(far_1_1941_0[0]));    relay_conn far_1_1941_0_b(.in(layer_0[942]), .out(far_1_1941_0[1]));
    wire [1:0] far_1_1941_1;    relay_conn far_1_1941_1_a(.in(far_1_1941_0[0]), .out(far_1_1941_1[0]));    relay_conn far_1_1941_1_b(.in(far_1_1941_0[1]), .out(far_1_1941_1[1]));
    assign layer_1[921] = ~far_1_1941_1[0] | (far_1_1941_1[0] & far_1_1941_1[1]); 
    wire [1:0] far_1_1942_0;    relay_conn far_1_1942_0_a(.in(layer_0[314]), .out(far_1_1942_0[0]));    relay_conn far_1_1942_0_b(.in(layer_0[354]), .out(far_1_1942_0[1]));
    assign layer_1[922] = far_1_1942_0[0] & far_1_1942_0[1]; 
    wire [1:0] far_1_1943_0;    relay_conn far_1_1943_0_a(.in(layer_0[623]), .out(far_1_1943_0[0]));    relay_conn far_1_1943_0_b(.in(layer_0[553]), .out(far_1_1943_0[1]));
    wire [1:0] far_1_1943_1;    relay_conn far_1_1943_1_a(.in(far_1_1943_0[0]), .out(far_1_1943_1[0]));    relay_conn far_1_1943_1_b(.in(far_1_1943_0[1]), .out(far_1_1943_1[1]));
    assign layer_1[923] = far_1_1943_1[0] | far_1_1943_1[1]; 
    assign layer_1[924] = ~layer_0[67] | (layer_0[91] & layer_0[67]); 
    wire [1:0] far_1_1945_0;    relay_conn far_1_1945_0_a(.in(layer_0[701]), .out(far_1_1945_0[0]));    relay_conn far_1_1945_0_b(.in(layer_0[768]), .out(far_1_1945_0[1]));
    wire [1:0] far_1_1945_1;    relay_conn far_1_1945_1_a(.in(far_1_1945_0[0]), .out(far_1_1945_1[0]));    relay_conn far_1_1945_1_b(.in(far_1_1945_0[1]), .out(far_1_1945_1[1]));
    assign layer_1[925] = ~(far_1_1945_1[0] ^ far_1_1945_1[1]); 
    wire [1:0] far_1_1946_0;    relay_conn far_1_1946_0_a(.in(layer_0[918]), .out(far_1_1946_0[0]));    relay_conn far_1_1946_0_b(.in(layer_0[881]), .out(far_1_1946_0[1]));
    assign layer_1[926] = far_1_1946_0[0] | far_1_1946_0[1]; 
    wire [1:0] far_1_1947_0;    relay_conn far_1_1947_0_a(.in(layer_0[397]), .out(far_1_1947_0[0]));    relay_conn far_1_1947_0_b(.in(layer_0[522]), .out(far_1_1947_0[1]));
    wire [1:0] far_1_1947_1;    relay_conn far_1_1947_1_a(.in(far_1_1947_0[0]), .out(far_1_1947_1[0]));    relay_conn far_1_1947_1_b(.in(far_1_1947_0[1]), .out(far_1_1947_1[1]));
    wire [1:0] far_1_1947_2;    relay_conn far_1_1947_2_a(.in(far_1_1947_1[0]), .out(far_1_1947_2[0]));    relay_conn far_1_1947_2_b(.in(far_1_1947_1[1]), .out(far_1_1947_2[1]));
    assign layer_1[927] = far_1_1947_2[1] & ~far_1_1947_2[0]; 
    assign layer_1[928] = layer_0[906] & layer_0[919]; 
    assign layer_1[929] = ~layer_0[816]; 
    wire [1:0] far_1_1950_0;    relay_conn far_1_1950_0_a(.in(layer_0[304]), .out(far_1_1950_0[0]));    relay_conn far_1_1950_0_b(.in(layer_0[402]), .out(far_1_1950_0[1]));
    wire [1:0] far_1_1950_1;    relay_conn far_1_1950_1_a(.in(far_1_1950_0[0]), .out(far_1_1950_1[0]));    relay_conn far_1_1950_1_b(.in(far_1_1950_0[1]), .out(far_1_1950_1[1]));
    wire [1:0] far_1_1950_2;    relay_conn far_1_1950_2_a(.in(far_1_1950_1[0]), .out(far_1_1950_2[0]));    relay_conn far_1_1950_2_b(.in(far_1_1950_1[1]), .out(far_1_1950_2[1]));
    assign layer_1[930] = ~(far_1_1950_2[0] ^ far_1_1950_2[1]); 
    wire [1:0] far_1_1951_0;    relay_conn far_1_1951_0_a(.in(layer_0[173]), .out(far_1_1951_0[0]));    relay_conn far_1_1951_0_b(.in(layer_0[261]), .out(far_1_1951_0[1]));
    wire [1:0] far_1_1951_1;    relay_conn far_1_1951_1_a(.in(far_1_1951_0[0]), .out(far_1_1951_1[0]));    relay_conn far_1_1951_1_b(.in(far_1_1951_0[1]), .out(far_1_1951_1[1]));
    assign layer_1[931] = far_1_1951_1[1]; 
    assign layer_1[932] = ~layer_0[141] | (layer_0[141] & layer_0[148]); 
    assign layer_1[933] = layer_0[43] ^ layer_0[61]; 
    wire [1:0] far_1_1954_0;    relay_conn far_1_1954_0_a(.in(layer_0[976]), .out(far_1_1954_0[0]));    relay_conn far_1_1954_0_b(.in(layer_0[849]), .out(far_1_1954_0[1]));
    wire [1:0] far_1_1954_1;    relay_conn far_1_1954_1_a(.in(far_1_1954_0[0]), .out(far_1_1954_1[0]));    relay_conn far_1_1954_1_b(.in(far_1_1954_0[1]), .out(far_1_1954_1[1]));
    wire [1:0] far_1_1954_2;    relay_conn far_1_1954_2_a(.in(far_1_1954_1[0]), .out(far_1_1954_2[0]));    relay_conn far_1_1954_2_b(.in(far_1_1954_1[1]), .out(far_1_1954_2[1]));
    assign layer_1[934] = ~(far_1_1954_2[0] ^ far_1_1954_2[1]); 
    wire [1:0] far_1_1955_0;    relay_conn far_1_1955_0_a(.in(layer_0[392]), .out(far_1_1955_0[0]));    relay_conn far_1_1955_0_b(.in(layer_0[512]), .out(far_1_1955_0[1]));
    wire [1:0] far_1_1955_1;    relay_conn far_1_1955_1_a(.in(far_1_1955_0[0]), .out(far_1_1955_1[0]));    relay_conn far_1_1955_1_b(.in(far_1_1955_0[1]), .out(far_1_1955_1[1]));
    wire [1:0] far_1_1955_2;    relay_conn far_1_1955_2_a(.in(far_1_1955_1[0]), .out(far_1_1955_2[0]));    relay_conn far_1_1955_2_b(.in(far_1_1955_1[1]), .out(far_1_1955_2[1]));
    assign layer_1[935] = far_1_1955_2[0]; 
    wire [1:0] far_1_1956_0;    relay_conn far_1_1956_0_a(.in(layer_0[775]), .out(far_1_1956_0[0]));    relay_conn far_1_1956_0_b(.in(layer_0[843]), .out(far_1_1956_0[1]));
    wire [1:0] far_1_1956_1;    relay_conn far_1_1956_1_a(.in(far_1_1956_0[0]), .out(far_1_1956_1[0]));    relay_conn far_1_1956_1_b(.in(far_1_1956_0[1]), .out(far_1_1956_1[1]));
    assign layer_1[936] = far_1_1956_1[0] ^ far_1_1956_1[1]; 
    wire [1:0] far_1_1957_0;    relay_conn far_1_1957_0_a(.in(layer_0[676]), .out(far_1_1957_0[0]));    relay_conn far_1_1957_0_b(.in(layer_0[559]), .out(far_1_1957_0[1]));
    wire [1:0] far_1_1957_1;    relay_conn far_1_1957_1_a(.in(far_1_1957_0[0]), .out(far_1_1957_1[0]));    relay_conn far_1_1957_1_b(.in(far_1_1957_0[1]), .out(far_1_1957_1[1]));
    wire [1:0] far_1_1957_2;    relay_conn far_1_1957_2_a(.in(far_1_1957_1[0]), .out(far_1_1957_2[0]));    relay_conn far_1_1957_2_b(.in(far_1_1957_1[1]), .out(far_1_1957_2[1]));
    assign layer_1[937] = far_1_1957_2[1] & ~far_1_1957_2[0]; 
    wire [1:0] far_1_1958_0;    relay_conn far_1_1958_0_a(.in(layer_0[614]), .out(far_1_1958_0[0]));    relay_conn far_1_1958_0_b(.in(layer_0[669]), .out(far_1_1958_0[1]));
    assign layer_1[938] = ~far_1_1958_0[0] | (far_1_1958_0[0] & far_1_1958_0[1]); 
    assign layer_1[939] = ~(layer_0[909] ^ layer_0[917]); 
    wire [1:0] far_1_1960_0;    relay_conn far_1_1960_0_a(.in(layer_0[312]), .out(far_1_1960_0[0]));    relay_conn far_1_1960_0_b(.in(layer_0[192]), .out(far_1_1960_0[1]));
    wire [1:0] far_1_1960_1;    relay_conn far_1_1960_1_a(.in(far_1_1960_0[0]), .out(far_1_1960_1[0]));    relay_conn far_1_1960_1_b(.in(far_1_1960_0[1]), .out(far_1_1960_1[1]));
    wire [1:0] far_1_1960_2;    relay_conn far_1_1960_2_a(.in(far_1_1960_1[0]), .out(far_1_1960_2[0]));    relay_conn far_1_1960_2_b(.in(far_1_1960_1[1]), .out(far_1_1960_2[1]));
    assign layer_1[940] = ~(far_1_1960_2[0] & far_1_1960_2[1]); 
    wire [1:0] far_1_1961_0;    relay_conn far_1_1961_0_a(.in(layer_0[682]), .out(far_1_1961_0[0]));    relay_conn far_1_1961_0_b(.in(layer_0[573]), .out(far_1_1961_0[1]));
    wire [1:0] far_1_1961_1;    relay_conn far_1_1961_1_a(.in(far_1_1961_0[0]), .out(far_1_1961_1[0]));    relay_conn far_1_1961_1_b(.in(far_1_1961_0[1]), .out(far_1_1961_1[1]));
    wire [1:0] far_1_1961_2;    relay_conn far_1_1961_2_a(.in(far_1_1961_1[0]), .out(far_1_1961_2[0]));    relay_conn far_1_1961_2_b(.in(far_1_1961_1[1]), .out(far_1_1961_2[1]));
    assign layer_1[941] = far_1_1961_2[1]; 
    wire [1:0] far_1_1962_0;    relay_conn far_1_1962_0_a(.in(layer_0[65]), .out(far_1_1962_0[0]));    relay_conn far_1_1962_0_b(.in(layer_0[111]), .out(far_1_1962_0[1]));
    assign layer_1[942] = ~far_1_1962_0[1] | (far_1_1962_0[0] & far_1_1962_0[1]); 
    wire [1:0] far_1_1963_0;    relay_conn far_1_1963_0_a(.in(layer_0[638]), .out(far_1_1963_0[0]));    relay_conn far_1_1963_0_b(.in(layer_0[553]), .out(far_1_1963_0[1]));
    wire [1:0] far_1_1963_1;    relay_conn far_1_1963_1_a(.in(far_1_1963_0[0]), .out(far_1_1963_1[0]));    relay_conn far_1_1963_1_b(.in(far_1_1963_0[1]), .out(far_1_1963_1[1]));
    assign layer_1[943] = far_1_1963_1[1] & ~far_1_1963_1[0]; 
    wire [1:0] far_1_1964_0;    relay_conn far_1_1964_0_a(.in(layer_0[68]), .out(far_1_1964_0[0]));    relay_conn far_1_1964_0_b(.in(layer_0[134]), .out(far_1_1964_0[1]));
    wire [1:0] far_1_1964_1;    relay_conn far_1_1964_1_a(.in(far_1_1964_0[0]), .out(far_1_1964_1[0]));    relay_conn far_1_1964_1_b(.in(far_1_1964_0[1]), .out(far_1_1964_1[1]));
    assign layer_1[944] = ~far_1_1964_1[1]; 
    wire [1:0] far_1_1965_0;    relay_conn far_1_1965_0_a(.in(layer_0[614]), .out(far_1_1965_0[0]));    relay_conn far_1_1965_0_b(.in(layer_0[710]), .out(far_1_1965_0[1]));
    wire [1:0] far_1_1965_1;    relay_conn far_1_1965_1_a(.in(far_1_1965_0[0]), .out(far_1_1965_1[0]));    relay_conn far_1_1965_1_b(.in(far_1_1965_0[1]), .out(far_1_1965_1[1]));
    wire [1:0] far_1_1965_2;    relay_conn far_1_1965_2_a(.in(far_1_1965_1[0]), .out(far_1_1965_2[0]));    relay_conn far_1_1965_2_b(.in(far_1_1965_1[1]), .out(far_1_1965_2[1]));
    assign layer_1[945] = ~(far_1_1965_2[0] | far_1_1965_2[1]); 
    wire [1:0] far_1_1966_0;    relay_conn far_1_1966_0_a(.in(layer_0[530]), .out(far_1_1966_0[0]));    relay_conn far_1_1966_0_b(.in(layer_0[438]), .out(far_1_1966_0[1]));
    wire [1:0] far_1_1966_1;    relay_conn far_1_1966_1_a(.in(far_1_1966_0[0]), .out(far_1_1966_1[0]));    relay_conn far_1_1966_1_b(.in(far_1_1966_0[1]), .out(far_1_1966_1[1]));
    assign layer_1[946] = far_1_1966_1[0] | far_1_1966_1[1]; 
    wire [1:0] far_1_1967_0;    relay_conn far_1_1967_0_a(.in(layer_0[450]), .out(far_1_1967_0[0]));    relay_conn far_1_1967_0_b(.in(layer_0[559]), .out(far_1_1967_0[1]));
    wire [1:0] far_1_1967_1;    relay_conn far_1_1967_1_a(.in(far_1_1967_0[0]), .out(far_1_1967_1[0]));    relay_conn far_1_1967_1_b(.in(far_1_1967_0[1]), .out(far_1_1967_1[1]));
    wire [1:0] far_1_1967_2;    relay_conn far_1_1967_2_a(.in(far_1_1967_1[0]), .out(far_1_1967_2[0]));    relay_conn far_1_1967_2_b(.in(far_1_1967_1[1]), .out(far_1_1967_2[1]));
    assign layer_1[947] = far_1_1967_2[0]; 
    wire [1:0] far_1_1968_0;    relay_conn far_1_1968_0_a(.in(layer_0[114]), .out(far_1_1968_0[0]));    relay_conn far_1_1968_0_b(.in(layer_0[242]), .out(far_1_1968_0[1]));
    wire [1:0] far_1_1968_1;    relay_conn far_1_1968_1_a(.in(far_1_1968_0[0]), .out(far_1_1968_1[0]));    relay_conn far_1_1968_1_b(.in(far_1_1968_0[1]), .out(far_1_1968_1[1]));
    wire [1:0] far_1_1968_2;    relay_conn far_1_1968_2_a(.in(far_1_1968_1[0]), .out(far_1_1968_2[0]));    relay_conn far_1_1968_2_b(.in(far_1_1968_1[1]), .out(far_1_1968_2[1]));
    wire [1:0] far_1_1968_3;    relay_conn far_1_1968_3_a(.in(far_1_1968_2[0]), .out(far_1_1968_3[0]));    relay_conn far_1_1968_3_b(.in(far_1_1968_2[1]), .out(far_1_1968_3[1]));
    assign layer_1[948] = far_1_1968_3[0] ^ far_1_1968_3[1]; 
    wire [1:0] far_1_1969_0;    relay_conn far_1_1969_0_a(.in(layer_0[302]), .out(far_1_1969_0[0]));    relay_conn far_1_1969_0_b(.in(layer_0[210]), .out(far_1_1969_0[1]));
    wire [1:0] far_1_1969_1;    relay_conn far_1_1969_1_a(.in(far_1_1969_0[0]), .out(far_1_1969_1[0]));    relay_conn far_1_1969_1_b(.in(far_1_1969_0[1]), .out(far_1_1969_1[1]));
    assign layer_1[949] = far_1_1969_1[1]; 
    wire [1:0] far_1_1970_0;    relay_conn far_1_1970_0_a(.in(layer_0[656]), .out(far_1_1970_0[0]));    relay_conn far_1_1970_0_b(.in(layer_0[543]), .out(far_1_1970_0[1]));
    wire [1:0] far_1_1970_1;    relay_conn far_1_1970_1_a(.in(far_1_1970_0[0]), .out(far_1_1970_1[0]));    relay_conn far_1_1970_1_b(.in(far_1_1970_0[1]), .out(far_1_1970_1[1]));
    wire [1:0] far_1_1970_2;    relay_conn far_1_1970_2_a(.in(far_1_1970_1[0]), .out(far_1_1970_2[0]));    relay_conn far_1_1970_2_b(.in(far_1_1970_1[1]), .out(far_1_1970_2[1]));
    assign layer_1[950] = far_1_1970_2[0] | far_1_1970_2[1]; 
    wire [1:0] far_1_1971_0;    relay_conn far_1_1971_0_a(.in(layer_0[98]), .out(far_1_1971_0[0]));    relay_conn far_1_1971_0_b(.in(layer_0[62]), .out(far_1_1971_0[1]));
    assign layer_1[951] = ~(far_1_1971_0[0] & far_1_1971_0[1]); 
    wire [1:0] far_1_1972_0;    relay_conn far_1_1972_0_a(.in(layer_0[1007]), .out(far_1_1972_0[0]));    relay_conn far_1_1972_0_b(.in(layer_0[973]), .out(far_1_1972_0[1]));
    assign layer_1[952] = ~far_1_1972_0[1]; 
    wire [1:0] far_1_1973_0;    relay_conn far_1_1973_0_a(.in(layer_0[140]), .out(far_1_1973_0[0]));    relay_conn far_1_1973_0_b(.in(layer_0[210]), .out(far_1_1973_0[1]));
    wire [1:0] far_1_1973_1;    relay_conn far_1_1973_1_a(.in(far_1_1973_0[0]), .out(far_1_1973_1[0]));    relay_conn far_1_1973_1_b(.in(far_1_1973_0[1]), .out(far_1_1973_1[1]));
    assign layer_1[953] = far_1_1973_1[0] | far_1_1973_1[1]; 
    wire [1:0] far_1_1974_0;    relay_conn far_1_1974_0_a(.in(layer_0[21]), .out(far_1_1974_0[0]));    relay_conn far_1_1974_0_b(.in(layer_0[91]), .out(far_1_1974_0[1]));
    wire [1:0] far_1_1974_1;    relay_conn far_1_1974_1_a(.in(far_1_1974_0[0]), .out(far_1_1974_1[0]));    relay_conn far_1_1974_1_b(.in(far_1_1974_0[1]), .out(far_1_1974_1[1]));
    assign layer_1[954] = ~(far_1_1974_1[0] | far_1_1974_1[1]); 
    wire [1:0] far_1_1975_0;    relay_conn far_1_1975_0_a(.in(layer_0[515]), .out(far_1_1975_0[0]));    relay_conn far_1_1975_0_b(.in(layer_0[413]), .out(far_1_1975_0[1]));
    wire [1:0] far_1_1975_1;    relay_conn far_1_1975_1_a(.in(far_1_1975_0[0]), .out(far_1_1975_1[0]));    relay_conn far_1_1975_1_b(.in(far_1_1975_0[1]), .out(far_1_1975_1[1]));
    wire [1:0] far_1_1975_2;    relay_conn far_1_1975_2_a(.in(far_1_1975_1[0]), .out(far_1_1975_2[0]));    relay_conn far_1_1975_2_b(.in(far_1_1975_1[1]), .out(far_1_1975_2[1]));
    assign layer_1[955] = ~(far_1_1975_2[0] | far_1_1975_2[1]); 
    wire [1:0] far_1_1976_0;    relay_conn far_1_1976_0_a(.in(layer_0[891]), .out(far_1_1976_0[0]));    relay_conn far_1_1976_0_b(.in(layer_0[1002]), .out(far_1_1976_0[1]));
    wire [1:0] far_1_1976_1;    relay_conn far_1_1976_1_a(.in(far_1_1976_0[0]), .out(far_1_1976_1[0]));    relay_conn far_1_1976_1_b(.in(far_1_1976_0[1]), .out(far_1_1976_1[1]));
    wire [1:0] far_1_1976_2;    relay_conn far_1_1976_2_a(.in(far_1_1976_1[0]), .out(far_1_1976_2[0]));    relay_conn far_1_1976_2_b(.in(far_1_1976_1[1]), .out(far_1_1976_2[1]));
    assign layer_1[956] = far_1_1976_2[0] | far_1_1976_2[1]; 
    wire [1:0] far_1_1977_0;    relay_conn far_1_1977_0_a(.in(layer_0[584]), .out(far_1_1977_0[0]));    relay_conn far_1_1977_0_b(.in(layer_0[656]), .out(far_1_1977_0[1]));
    wire [1:0] far_1_1977_1;    relay_conn far_1_1977_1_a(.in(far_1_1977_0[0]), .out(far_1_1977_1[0]));    relay_conn far_1_1977_1_b(.in(far_1_1977_0[1]), .out(far_1_1977_1[1]));
    assign layer_1[957] = ~(far_1_1977_1[0] ^ far_1_1977_1[1]); 
    wire [1:0] far_1_1978_0;    relay_conn far_1_1978_0_a(.in(layer_0[610]), .out(far_1_1978_0[0]));    relay_conn far_1_1978_0_b(.in(layer_0[735]), .out(far_1_1978_0[1]));
    wire [1:0] far_1_1978_1;    relay_conn far_1_1978_1_a(.in(far_1_1978_0[0]), .out(far_1_1978_1[0]));    relay_conn far_1_1978_1_b(.in(far_1_1978_0[1]), .out(far_1_1978_1[1]));
    wire [1:0] far_1_1978_2;    relay_conn far_1_1978_2_a(.in(far_1_1978_1[0]), .out(far_1_1978_2[0]));    relay_conn far_1_1978_2_b(.in(far_1_1978_1[1]), .out(far_1_1978_2[1]));
    assign layer_1[958] = far_1_1978_2[0] & far_1_1978_2[1]; 
    wire [1:0] far_1_1979_0;    relay_conn far_1_1979_0_a(.in(layer_0[741]), .out(far_1_1979_0[0]));    relay_conn far_1_1979_0_b(.in(layer_0[806]), .out(far_1_1979_0[1]));
    wire [1:0] far_1_1979_1;    relay_conn far_1_1979_1_a(.in(far_1_1979_0[0]), .out(far_1_1979_1[0]));    relay_conn far_1_1979_1_b(.in(far_1_1979_0[1]), .out(far_1_1979_1[1]));
    assign layer_1[959] = ~far_1_1979_1[0]; 
    assign layer_1[960] = layer_0[908] ^ layer_0[916]; 
    wire [1:0] far_1_1981_0;    relay_conn far_1_1981_0_a(.in(layer_0[321]), .out(far_1_1981_0[0]));    relay_conn far_1_1981_0_b(.in(layer_0[241]), .out(far_1_1981_0[1]));
    wire [1:0] far_1_1981_1;    relay_conn far_1_1981_1_a(.in(far_1_1981_0[0]), .out(far_1_1981_1[0]));    relay_conn far_1_1981_1_b(.in(far_1_1981_0[1]), .out(far_1_1981_1[1]));
    assign layer_1[961] = far_1_1981_1[1]; 
    wire [1:0] far_1_1982_0;    relay_conn far_1_1982_0_a(.in(layer_0[117]), .out(far_1_1982_0[0]));    relay_conn far_1_1982_0_b(.in(layer_0[219]), .out(far_1_1982_0[1]));
    wire [1:0] far_1_1982_1;    relay_conn far_1_1982_1_a(.in(far_1_1982_0[0]), .out(far_1_1982_1[0]));    relay_conn far_1_1982_1_b(.in(far_1_1982_0[1]), .out(far_1_1982_1[1]));
    wire [1:0] far_1_1982_2;    relay_conn far_1_1982_2_a(.in(far_1_1982_1[0]), .out(far_1_1982_2[0]));    relay_conn far_1_1982_2_b(.in(far_1_1982_1[1]), .out(far_1_1982_2[1]));
    assign layer_1[962] = ~far_1_1982_2[0]; 
    assign layer_1[963] = layer_0[676] & ~layer_0[651]; 
    wire [1:0] far_1_1984_0;    relay_conn far_1_1984_0_a(.in(layer_0[821]), .out(far_1_1984_0[0]));    relay_conn far_1_1984_0_b(.in(layer_0[773]), .out(far_1_1984_0[1]));
    assign layer_1[964] = ~far_1_1984_0[0] | (far_1_1984_0[0] & far_1_1984_0[1]); 
    wire [1:0] far_1_1985_0;    relay_conn far_1_1985_0_a(.in(layer_0[500]), .out(far_1_1985_0[0]));    relay_conn far_1_1985_0_b(.in(layer_0[412]), .out(far_1_1985_0[1]));
    wire [1:0] far_1_1985_1;    relay_conn far_1_1985_1_a(.in(far_1_1985_0[0]), .out(far_1_1985_1[0]));    relay_conn far_1_1985_1_b(.in(far_1_1985_0[1]), .out(far_1_1985_1[1]));
    assign layer_1[965] = ~far_1_1985_1[0]; 
    wire [1:0] far_1_1986_0;    relay_conn far_1_1986_0_a(.in(layer_0[242]), .out(far_1_1986_0[0]));    relay_conn far_1_1986_0_b(.in(layer_0[336]), .out(far_1_1986_0[1]));
    wire [1:0] far_1_1986_1;    relay_conn far_1_1986_1_a(.in(far_1_1986_0[0]), .out(far_1_1986_1[0]));    relay_conn far_1_1986_1_b(.in(far_1_1986_0[1]), .out(far_1_1986_1[1]));
    assign layer_1[966] = far_1_1986_1[1]; 
    assign layer_1[967] = layer_0[679] | layer_0[669]; 
    wire [1:0] far_1_1988_0;    relay_conn far_1_1988_0_a(.in(layer_0[584]), .out(far_1_1988_0[0]));    relay_conn far_1_1988_0_b(.in(layer_0[543]), .out(far_1_1988_0[1]));
    assign layer_1[968] = ~(far_1_1988_0[0] & far_1_1988_0[1]); 
    assign layer_1[969] = ~layer_0[98]; 
    wire [1:0] far_1_1990_0;    relay_conn far_1_1990_0_a(.in(layer_0[1002]), .out(far_1_1990_0[0]));    relay_conn far_1_1990_0_b(.in(layer_0[897]), .out(far_1_1990_0[1]));
    wire [1:0] far_1_1990_1;    relay_conn far_1_1990_1_a(.in(far_1_1990_0[0]), .out(far_1_1990_1[0]));    relay_conn far_1_1990_1_b(.in(far_1_1990_0[1]), .out(far_1_1990_1[1]));
    wire [1:0] far_1_1990_2;    relay_conn far_1_1990_2_a(.in(far_1_1990_1[0]), .out(far_1_1990_2[0]));    relay_conn far_1_1990_2_b(.in(far_1_1990_1[1]), .out(far_1_1990_2[1]));
    assign layer_1[970] = ~far_1_1990_2[1] | (far_1_1990_2[0] & far_1_1990_2[1]); 
    assign layer_1[971] = layer_0[419] ^ layer_0[443]; 
    wire [1:0] far_1_1992_0;    relay_conn far_1_1992_0_a(.in(layer_0[391]), .out(far_1_1992_0[0]));    relay_conn far_1_1992_0_b(.in(layer_0[504]), .out(far_1_1992_0[1]));
    wire [1:0] far_1_1992_1;    relay_conn far_1_1992_1_a(.in(far_1_1992_0[0]), .out(far_1_1992_1[0]));    relay_conn far_1_1992_1_b(.in(far_1_1992_0[1]), .out(far_1_1992_1[1]));
    wire [1:0] far_1_1992_2;    relay_conn far_1_1992_2_a(.in(far_1_1992_1[0]), .out(far_1_1992_2[0]));    relay_conn far_1_1992_2_b(.in(far_1_1992_1[1]), .out(far_1_1992_2[1]));
    assign layer_1[972] = far_1_1992_2[0] | far_1_1992_2[1]; 
    wire [1:0] far_1_1993_0;    relay_conn far_1_1993_0_a(.in(layer_0[614]), .out(far_1_1993_0[0]));    relay_conn far_1_1993_0_b(.in(layer_0[659]), .out(far_1_1993_0[1]));
    assign layer_1[973] = far_1_1993_0[0] & far_1_1993_0[1]; 
    wire [1:0] far_1_1994_0;    relay_conn far_1_1994_0_a(.in(layer_0[219]), .out(far_1_1994_0[0]));    relay_conn far_1_1994_0_b(.in(layer_0[143]), .out(far_1_1994_0[1]));
    wire [1:0] far_1_1994_1;    relay_conn far_1_1994_1_a(.in(far_1_1994_0[0]), .out(far_1_1994_1[0]));    relay_conn far_1_1994_1_b(.in(far_1_1994_0[1]), .out(far_1_1994_1[1]));
    assign layer_1[974] = ~(far_1_1994_1[0] & far_1_1994_1[1]); 
    wire [1:0] far_1_1995_0;    relay_conn far_1_1995_0_a(.in(layer_0[847]), .out(far_1_1995_0[0]));    relay_conn far_1_1995_0_b(.in(layer_0[798]), .out(far_1_1995_0[1]));
    assign layer_1[975] = ~(far_1_1995_0[0] & far_1_1995_0[1]); 
    assign layer_1[976] = ~(layer_0[824] & layer_0[852]); 
    wire [1:0] far_1_1997_0;    relay_conn far_1_1997_0_a(.in(layer_0[163]), .out(far_1_1997_0[0]));    relay_conn far_1_1997_0_b(.in(layer_0[246]), .out(far_1_1997_0[1]));
    wire [1:0] far_1_1997_1;    relay_conn far_1_1997_1_a(.in(far_1_1997_0[0]), .out(far_1_1997_1[0]));    relay_conn far_1_1997_1_b(.in(far_1_1997_0[1]), .out(far_1_1997_1[1]));
    assign layer_1[977] = ~(far_1_1997_1[0] ^ far_1_1997_1[1]); 
    wire [1:0] far_1_1998_0;    relay_conn far_1_1998_0_a(.in(layer_0[220]), .out(far_1_1998_0[0]));    relay_conn far_1_1998_0_b(.in(layer_0[109]), .out(far_1_1998_0[1]));
    wire [1:0] far_1_1998_1;    relay_conn far_1_1998_1_a(.in(far_1_1998_0[0]), .out(far_1_1998_1[0]));    relay_conn far_1_1998_1_b(.in(far_1_1998_0[1]), .out(far_1_1998_1[1]));
    wire [1:0] far_1_1998_2;    relay_conn far_1_1998_2_a(.in(far_1_1998_1[0]), .out(far_1_1998_2[0]));    relay_conn far_1_1998_2_b(.in(far_1_1998_1[1]), .out(far_1_1998_2[1]));
    assign layer_1[978] = far_1_1998_2[0] & far_1_1998_2[1]; 
    assign layer_1[979] = layer_0[116]; 
    wire [1:0] far_1_2000_0;    relay_conn far_1_2000_0_a(.in(layer_0[590]), .out(far_1_2000_0[0]));    relay_conn far_1_2000_0_b(.in(layer_0[495]), .out(far_1_2000_0[1]));
    wire [1:0] far_1_2000_1;    relay_conn far_1_2000_1_a(.in(far_1_2000_0[0]), .out(far_1_2000_1[0]));    relay_conn far_1_2000_1_b(.in(far_1_2000_0[1]), .out(far_1_2000_1[1]));
    assign layer_1[980] = far_1_2000_1[0] | far_1_2000_1[1]; 
    wire [1:0] far_1_2001_0;    relay_conn far_1_2001_0_a(.in(layer_0[663]), .out(far_1_2001_0[0]));    relay_conn far_1_2001_0_b(.in(layer_0[731]), .out(far_1_2001_0[1]));
    wire [1:0] far_1_2001_1;    relay_conn far_1_2001_1_a(.in(far_1_2001_0[0]), .out(far_1_2001_1[0]));    relay_conn far_1_2001_1_b(.in(far_1_2001_0[1]), .out(far_1_2001_1[1]));
    assign layer_1[981] = ~(far_1_2001_1[0] & far_1_2001_1[1]); 
    assign layer_1[982] = layer_0[659]; 
    assign layer_1[983] = ~(layer_0[894] ^ layer_0[865]); 
    wire [1:0] far_1_2004_0;    relay_conn far_1_2004_0_a(.in(layer_0[110]), .out(far_1_2004_0[0]));    relay_conn far_1_2004_0_b(.in(layer_0[64]), .out(far_1_2004_0[1]));
    assign layer_1[984] = far_1_2004_0[1] & ~far_1_2004_0[0]; 
    wire [1:0] far_1_2005_0;    relay_conn far_1_2005_0_a(.in(layer_0[923]), .out(far_1_2005_0[0]));    relay_conn far_1_2005_0_b(.in(layer_0[956]), .out(far_1_2005_0[1]));
    assign layer_1[985] = far_1_2005_0[1]; 
    wire [1:0] far_1_2006_0;    relay_conn far_1_2006_0_a(.in(layer_0[923]), .out(far_1_2006_0[0]));    relay_conn far_1_2006_0_b(.in(layer_0[855]), .out(far_1_2006_0[1]));
    wire [1:0] far_1_2006_1;    relay_conn far_1_2006_1_a(.in(far_1_2006_0[0]), .out(far_1_2006_1[0]));    relay_conn far_1_2006_1_b(.in(far_1_2006_0[1]), .out(far_1_2006_1[1]));
    assign layer_1[986] = far_1_2006_1[0] & far_1_2006_1[1]; 
    assign layer_1[987] = layer_0[131] | layer_0[107]; 
    wire [1:0] far_1_2008_0;    relay_conn far_1_2008_0_a(.in(layer_0[867]), .out(far_1_2008_0[0]));    relay_conn far_1_2008_0_b(.in(layer_0[983]), .out(far_1_2008_0[1]));
    wire [1:0] far_1_2008_1;    relay_conn far_1_2008_1_a(.in(far_1_2008_0[0]), .out(far_1_2008_1[0]));    relay_conn far_1_2008_1_b(.in(far_1_2008_0[1]), .out(far_1_2008_1[1]));
    wire [1:0] far_1_2008_2;    relay_conn far_1_2008_2_a(.in(far_1_2008_1[0]), .out(far_1_2008_2[0]));    relay_conn far_1_2008_2_b(.in(far_1_2008_1[1]), .out(far_1_2008_2[1]));
    assign layer_1[988] = ~(far_1_2008_2[0] & far_1_2008_2[1]); 
    wire [1:0] far_1_2009_0;    relay_conn far_1_2009_0_a(.in(layer_0[323]), .out(far_1_2009_0[0]));    relay_conn far_1_2009_0_b(.in(layer_0[446]), .out(far_1_2009_0[1]));
    wire [1:0] far_1_2009_1;    relay_conn far_1_2009_1_a(.in(far_1_2009_0[0]), .out(far_1_2009_1[0]));    relay_conn far_1_2009_1_b(.in(far_1_2009_0[1]), .out(far_1_2009_1[1]));
    wire [1:0] far_1_2009_2;    relay_conn far_1_2009_2_a(.in(far_1_2009_1[0]), .out(far_1_2009_2[0]));    relay_conn far_1_2009_2_b(.in(far_1_2009_1[1]), .out(far_1_2009_2[1]));
    assign layer_1[989] = ~far_1_2009_2[1] | (far_1_2009_2[0] & far_1_2009_2[1]); 
    assign layer_1[990] = ~(layer_0[91] | layer_0[119]); 
    wire [1:0] far_1_2011_0;    relay_conn far_1_2011_0_a(.in(layer_0[91]), .out(far_1_2011_0[0]));    relay_conn far_1_2011_0_b(.in(layer_0[21]), .out(far_1_2011_0[1]));
    wire [1:0] far_1_2011_1;    relay_conn far_1_2011_1_a(.in(far_1_2011_0[0]), .out(far_1_2011_1[0]));    relay_conn far_1_2011_1_b(.in(far_1_2011_0[1]), .out(far_1_2011_1[1]));
    assign layer_1[991] = far_1_2011_1[1]; 
    assign layer_1[992] = layer_0[362] & ~layer_0[373]; 
    assign layer_1[993] = layer_0[283] & ~layer_0[301]; 
    wire [1:0] far_1_2014_0;    relay_conn far_1_2014_0_a(.in(layer_0[484]), .out(far_1_2014_0[0]));    relay_conn far_1_2014_0_b(.in(layer_0[543]), .out(far_1_2014_0[1]));
    assign layer_1[994] = ~(far_1_2014_0[0] & far_1_2014_0[1]); 
    wire [1:0] far_1_2015_0;    relay_conn far_1_2015_0_a(.in(layer_0[208]), .out(far_1_2015_0[0]));    relay_conn far_1_2015_0_b(.in(layer_0[256]), .out(far_1_2015_0[1]));
    assign layer_1[995] = far_1_2015_0[1] & ~far_1_2015_0[0]; 
    wire [1:0] far_1_2016_0;    relay_conn far_1_2016_0_a(.in(layer_0[560]), .out(far_1_2016_0[0]));    relay_conn far_1_2016_0_b(.in(layer_0[659]), .out(far_1_2016_0[1]));
    wire [1:0] far_1_2016_1;    relay_conn far_1_2016_1_a(.in(far_1_2016_0[0]), .out(far_1_2016_1[0]));    relay_conn far_1_2016_1_b(.in(far_1_2016_0[1]), .out(far_1_2016_1[1]));
    wire [1:0] far_1_2016_2;    relay_conn far_1_2016_2_a(.in(far_1_2016_1[0]), .out(far_1_2016_2[0]));    relay_conn far_1_2016_2_b(.in(far_1_2016_1[1]), .out(far_1_2016_2[1]));
    assign layer_1[996] = far_1_2016_2[1] & ~far_1_2016_2[0]; 
    wire [1:0] far_1_2017_0;    relay_conn far_1_2017_0_a(.in(layer_0[419]), .out(far_1_2017_0[0]));    relay_conn far_1_2017_0_b(.in(layer_0[355]), .out(far_1_2017_0[1]));
    wire [1:0] far_1_2017_1;    relay_conn far_1_2017_1_a(.in(far_1_2017_0[0]), .out(far_1_2017_1[0]));    relay_conn far_1_2017_1_b(.in(far_1_2017_0[1]), .out(far_1_2017_1[1]));
    assign layer_1[997] = far_1_2017_1[0] & ~far_1_2017_1[1]; 
    wire [1:0] far_1_2018_0;    relay_conn far_1_2018_0_a(.in(layer_0[381]), .out(far_1_2018_0[0]));    relay_conn far_1_2018_0_b(.in(layer_0[430]), .out(far_1_2018_0[1]));
    assign layer_1[998] = far_1_2018_0[1]; 
    wire [1:0] far_1_2019_0;    relay_conn far_1_2019_0_a(.in(layer_0[365]), .out(far_1_2019_0[0]));    relay_conn far_1_2019_0_b(.in(layer_0[438]), .out(far_1_2019_0[1]));
    wire [1:0] far_1_2019_1;    relay_conn far_1_2019_1_a(.in(far_1_2019_0[0]), .out(far_1_2019_1[0]));    relay_conn far_1_2019_1_b(.in(far_1_2019_0[1]), .out(far_1_2019_1[1]));
    assign layer_1[999] = far_1_2019_1[0] & ~far_1_2019_1[1]; 
    wire [1:0] far_1_2020_0;    relay_conn far_1_2020_0_a(.in(layer_0[339]), .out(far_1_2020_0[0]));    relay_conn far_1_2020_0_b(.in(layer_0[232]), .out(far_1_2020_0[1]));
    wire [1:0] far_1_2020_1;    relay_conn far_1_2020_1_a(.in(far_1_2020_0[0]), .out(far_1_2020_1[0]));    relay_conn far_1_2020_1_b(.in(far_1_2020_0[1]), .out(far_1_2020_1[1]));
    wire [1:0] far_1_2020_2;    relay_conn far_1_2020_2_a(.in(far_1_2020_1[0]), .out(far_1_2020_2[0]));    relay_conn far_1_2020_2_b(.in(far_1_2020_1[1]), .out(far_1_2020_2[1]));
    assign layer_1[1000] = ~far_1_2020_2[0]; 
    wire [1:0] far_1_2021_0;    relay_conn far_1_2021_0_a(.in(layer_0[10]), .out(far_1_2021_0[0]));    relay_conn far_1_2021_0_b(.in(layer_0[96]), .out(far_1_2021_0[1]));
    wire [1:0] far_1_2021_1;    relay_conn far_1_2021_1_a(.in(far_1_2021_0[0]), .out(far_1_2021_1[0]));    relay_conn far_1_2021_1_b(.in(far_1_2021_0[1]), .out(far_1_2021_1[1]));
    assign layer_1[1001] = ~(far_1_2021_1[0] & far_1_2021_1[1]); 
    wire [1:0] far_1_2022_0;    relay_conn far_1_2022_0_a(.in(layer_0[806]), .out(far_1_2022_0[0]));    relay_conn far_1_2022_0_b(.in(layer_0[930]), .out(far_1_2022_0[1]));
    wire [1:0] far_1_2022_1;    relay_conn far_1_2022_1_a(.in(far_1_2022_0[0]), .out(far_1_2022_1[0]));    relay_conn far_1_2022_1_b(.in(far_1_2022_0[1]), .out(far_1_2022_1[1]));
    wire [1:0] far_1_2022_2;    relay_conn far_1_2022_2_a(.in(far_1_2022_1[0]), .out(far_1_2022_2[0]));    relay_conn far_1_2022_2_b(.in(far_1_2022_1[1]), .out(far_1_2022_2[1]));
    assign layer_1[1002] = ~(far_1_2022_2[0] | far_1_2022_2[1]); 
    assign layer_1[1003] = ~layer_0[446] | (layer_0[446] & layer_0[471]); 
    wire [1:0] far_1_2024_0;    relay_conn far_1_2024_0_a(.in(layer_0[150]), .out(far_1_2024_0[0]));    relay_conn far_1_2024_0_b(.in(layer_0[204]), .out(far_1_2024_0[1]));
    assign layer_1[1004] = ~far_1_2024_0[0] | (far_1_2024_0[0] & far_1_2024_0[1]); 
    wire [1:0] far_1_2025_0;    relay_conn far_1_2025_0_a(.in(layer_0[314]), .out(far_1_2025_0[0]));    relay_conn far_1_2025_0_b(.in(layer_0[361]), .out(far_1_2025_0[1]));
    assign layer_1[1005] = ~far_1_2025_0[0] | (far_1_2025_0[0] & far_1_2025_0[1]); 
    assign layer_1[1006] = layer_0[442] ^ layer_0[472]; 
    wire [1:0] far_1_2027_0;    relay_conn far_1_2027_0_a(.in(layer_0[585]), .out(far_1_2027_0[0]));    relay_conn far_1_2027_0_b(.in(layer_0[468]), .out(far_1_2027_0[1]));
    wire [1:0] far_1_2027_1;    relay_conn far_1_2027_1_a(.in(far_1_2027_0[0]), .out(far_1_2027_1[0]));    relay_conn far_1_2027_1_b(.in(far_1_2027_0[1]), .out(far_1_2027_1[1]));
    wire [1:0] far_1_2027_2;    relay_conn far_1_2027_2_a(.in(far_1_2027_1[0]), .out(far_1_2027_2[0]));    relay_conn far_1_2027_2_b(.in(far_1_2027_1[1]), .out(far_1_2027_2[1]));
    assign layer_1[1007] = far_1_2027_2[1] & ~far_1_2027_2[0]; 
    wire [1:0] far_1_2028_0;    relay_conn far_1_2028_0_a(.in(layer_0[372]), .out(far_1_2028_0[0]));    relay_conn far_1_2028_0_b(.in(layer_0[463]), .out(far_1_2028_0[1]));
    wire [1:0] far_1_2028_1;    relay_conn far_1_2028_1_a(.in(far_1_2028_0[0]), .out(far_1_2028_1[0]));    relay_conn far_1_2028_1_b(.in(far_1_2028_0[1]), .out(far_1_2028_1[1]));
    assign layer_1[1008] = far_1_2028_1[0] & far_1_2028_1[1]; 
    wire [1:0] far_1_2029_0;    relay_conn far_1_2029_0_a(.in(layer_0[429]), .out(far_1_2029_0[0]));    relay_conn far_1_2029_0_b(.in(layer_0[313]), .out(far_1_2029_0[1]));
    wire [1:0] far_1_2029_1;    relay_conn far_1_2029_1_a(.in(far_1_2029_0[0]), .out(far_1_2029_1[0]));    relay_conn far_1_2029_1_b(.in(far_1_2029_0[1]), .out(far_1_2029_1[1]));
    wire [1:0] far_1_2029_2;    relay_conn far_1_2029_2_a(.in(far_1_2029_1[0]), .out(far_1_2029_2[0]));    relay_conn far_1_2029_2_b(.in(far_1_2029_1[1]), .out(far_1_2029_2[1]));
    assign layer_1[1009] = ~(far_1_2029_2[0] ^ far_1_2029_2[1]); 
    wire [1:0] far_1_2030_0;    relay_conn far_1_2030_0_a(.in(layer_0[539]), .out(far_1_2030_0[0]));    relay_conn far_1_2030_0_b(.in(layer_0[485]), .out(far_1_2030_0[1]));
    assign layer_1[1010] = far_1_2030_0[0]; 
    assign layer_1[1011] = layer_0[91] & layer_0[65]; 
    wire [1:0] far_1_2032_0;    relay_conn far_1_2032_0_a(.in(layer_0[367]), .out(far_1_2032_0[0]));    relay_conn far_1_2032_0_b(.in(layer_0[265]), .out(far_1_2032_0[1]));
    wire [1:0] far_1_2032_1;    relay_conn far_1_2032_1_a(.in(far_1_2032_0[0]), .out(far_1_2032_1[0]));    relay_conn far_1_2032_1_b(.in(far_1_2032_0[1]), .out(far_1_2032_1[1]));
    wire [1:0] far_1_2032_2;    relay_conn far_1_2032_2_a(.in(far_1_2032_1[0]), .out(far_1_2032_2[0]));    relay_conn far_1_2032_2_b(.in(far_1_2032_1[1]), .out(far_1_2032_2[1]));
    assign layer_1[1012] = ~(far_1_2032_2[0] | far_1_2032_2[1]); 
    wire [1:0] far_1_2033_0;    relay_conn far_1_2033_0_a(.in(layer_0[877]), .out(far_1_2033_0[0]));    relay_conn far_1_2033_0_b(.in(layer_0[924]), .out(far_1_2033_0[1]));
    assign layer_1[1013] = ~(far_1_2033_0[0] & far_1_2033_0[1]); 
    wire [1:0] far_1_2034_0;    relay_conn far_1_2034_0_a(.in(layer_0[377]), .out(far_1_2034_0[0]));    relay_conn far_1_2034_0_b(.in(layer_0[453]), .out(far_1_2034_0[1]));
    wire [1:0] far_1_2034_1;    relay_conn far_1_2034_1_a(.in(far_1_2034_0[0]), .out(far_1_2034_1[0]));    relay_conn far_1_2034_1_b(.in(far_1_2034_0[1]), .out(far_1_2034_1[1]));
    assign layer_1[1014] = ~(far_1_2034_1[0] ^ far_1_2034_1[1]); 
    wire [1:0] far_1_2035_0;    relay_conn far_1_2035_0_a(.in(layer_0[258]), .out(far_1_2035_0[0]));    relay_conn far_1_2035_0_b(.in(layer_0[172]), .out(far_1_2035_0[1]));
    wire [1:0] far_1_2035_1;    relay_conn far_1_2035_1_a(.in(far_1_2035_0[0]), .out(far_1_2035_1[0]));    relay_conn far_1_2035_1_b(.in(far_1_2035_0[1]), .out(far_1_2035_1[1]));
    assign layer_1[1015] = far_1_2035_1[0]; 
    wire [1:0] far_1_2036_0;    relay_conn far_1_2036_0_a(.in(layer_0[873]), .out(far_1_2036_0[0]));    relay_conn far_1_2036_0_b(.in(layer_0[785]), .out(far_1_2036_0[1]));
    wire [1:0] far_1_2036_1;    relay_conn far_1_2036_1_a(.in(far_1_2036_0[0]), .out(far_1_2036_1[0]));    relay_conn far_1_2036_1_b(.in(far_1_2036_0[1]), .out(far_1_2036_1[1]));
    assign layer_1[1016] = far_1_2036_1[0] ^ far_1_2036_1[1]; 
    assign layer_1[1017] = layer_0[841] & ~layer_0[857]; 
    assign layer_1[1018] = layer_0[876]; 
    assign layer_1[1019] = layer_0[448] | layer_0[429]; 
    // Layer 2 ============================================================
    wire [1:0] far_2_2040_0;    relay_conn far_2_2040_0_a(.in(layer_1[631]), .out(far_2_2040_0[0]));    relay_conn far_2_2040_0_b(.in(layer_1[743]), .out(far_2_2040_0[1]));
    wire [1:0] far_2_2040_1;    relay_conn far_2_2040_1_a(.in(far_2_2040_0[0]), .out(far_2_2040_1[0]));    relay_conn far_2_2040_1_b(.in(far_2_2040_0[1]), .out(far_2_2040_1[1]));
    wire [1:0] far_2_2040_2;    relay_conn far_2_2040_2_a(.in(far_2_2040_1[0]), .out(far_2_2040_2[0]));    relay_conn far_2_2040_2_b(.in(far_2_2040_1[1]), .out(far_2_2040_2[1]));
    assign layer_2[0] = far_2_2040_2[0] ^ far_2_2040_2[1]; 
    wire [1:0] far_2_2041_0;    relay_conn far_2_2041_0_a(.in(layer_1[303]), .out(far_2_2041_0[0]));    relay_conn far_2_2041_0_b(.in(layer_1[409]), .out(far_2_2041_0[1]));
    wire [1:0] far_2_2041_1;    relay_conn far_2_2041_1_a(.in(far_2_2041_0[0]), .out(far_2_2041_1[0]));    relay_conn far_2_2041_1_b(.in(far_2_2041_0[1]), .out(far_2_2041_1[1]));
    wire [1:0] far_2_2041_2;    relay_conn far_2_2041_2_a(.in(far_2_2041_1[0]), .out(far_2_2041_2[0]));    relay_conn far_2_2041_2_b(.in(far_2_2041_1[1]), .out(far_2_2041_2[1]));
    assign layer_2[1] = far_2_2041_2[0] & ~far_2_2041_2[1]; 
    assign layer_2[2] = layer_1[952]; 
    wire [1:0] far_2_2043_0;    relay_conn far_2_2043_0_a(.in(layer_1[280]), .out(far_2_2043_0[0]));    relay_conn far_2_2043_0_b(.in(layer_1[248]), .out(far_2_2043_0[1]));
    assign layer_2[3] = far_2_2043_0[0] | far_2_2043_0[1]; 
    wire [1:0] far_2_2044_0;    relay_conn far_2_2044_0_a(.in(layer_1[571]), .out(far_2_2044_0[0]));    relay_conn far_2_2044_0_b(.in(layer_1[507]), .out(far_2_2044_0[1]));
    wire [1:0] far_2_2044_1;    relay_conn far_2_2044_1_a(.in(far_2_2044_0[0]), .out(far_2_2044_1[0]));    relay_conn far_2_2044_1_b(.in(far_2_2044_0[1]), .out(far_2_2044_1[1]));
    assign layer_2[4] = ~far_2_2044_1[1] | (far_2_2044_1[0] & far_2_2044_1[1]); 
    wire [1:0] far_2_2045_0;    relay_conn far_2_2045_0_a(.in(layer_1[84]), .out(far_2_2045_0[0]));    relay_conn far_2_2045_0_b(.in(layer_1[21]), .out(far_2_2045_0[1]));
    assign layer_2[5] = far_2_2045_0[0] & far_2_2045_0[1]; 
    wire [1:0] far_2_2046_0;    relay_conn far_2_2046_0_a(.in(layer_1[410]), .out(far_2_2046_0[0]));    relay_conn far_2_2046_0_b(.in(layer_1[445]), .out(far_2_2046_0[1]));
    assign layer_2[6] = far_2_2046_0[1] & ~far_2_2046_0[0]; 
    wire [1:0] far_2_2047_0;    relay_conn far_2_2047_0_a(.in(layer_1[349]), .out(far_2_2047_0[0]));    relay_conn far_2_2047_0_b(.in(layer_1[248]), .out(far_2_2047_0[1]));
    wire [1:0] far_2_2047_1;    relay_conn far_2_2047_1_a(.in(far_2_2047_0[0]), .out(far_2_2047_1[0]));    relay_conn far_2_2047_1_b(.in(far_2_2047_0[1]), .out(far_2_2047_1[1]));
    wire [1:0] far_2_2047_2;    relay_conn far_2_2047_2_a(.in(far_2_2047_1[0]), .out(far_2_2047_2[0]));    relay_conn far_2_2047_2_b(.in(far_2_2047_1[1]), .out(far_2_2047_2[1]));
    assign layer_2[7] = far_2_2047_2[1] & ~far_2_2047_2[0]; 
    assign layer_2[8] = ~(layer_1[627] & layer_1[645]); 
    assign layer_2[9] = ~(layer_1[287] & layer_1[269]); 
    assign layer_2[10] = layer_1[574]; 
    wire [1:0] far_2_2051_0;    relay_conn far_2_2051_0_a(.in(layer_1[409]), .out(far_2_2051_0[0]));    relay_conn far_2_2051_0_b(.in(layer_1[467]), .out(far_2_2051_0[1]));
    assign layer_2[11] = ~far_2_2051_0[1] | (far_2_2051_0[0] & far_2_2051_0[1]); 
    wire [1:0] far_2_2052_0;    relay_conn far_2_2052_0_a(.in(layer_1[86]), .out(far_2_2052_0[0]));    relay_conn far_2_2052_0_b(.in(layer_1[127]), .out(far_2_2052_0[1]));
    assign layer_2[12] = far_2_2052_0[0] & far_2_2052_0[1]; 
    wire [1:0] far_2_2053_0;    relay_conn far_2_2053_0_a(.in(layer_1[219]), .out(far_2_2053_0[0]));    relay_conn far_2_2053_0_b(.in(layer_1[95]), .out(far_2_2053_0[1]));
    wire [1:0] far_2_2053_1;    relay_conn far_2_2053_1_a(.in(far_2_2053_0[0]), .out(far_2_2053_1[0]));    relay_conn far_2_2053_1_b(.in(far_2_2053_0[1]), .out(far_2_2053_1[1]));
    wire [1:0] far_2_2053_2;    relay_conn far_2_2053_2_a(.in(far_2_2053_1[0]), .out(far_2_2053_2[0]));    relay_conn far_2_2053_2_b(.in(far_2_2053_1[1]), .out(far_2_2053_2[1]));
    assign layer_2[13] = ~(far_2_2053_2[0] & far_2_2053_2[1]); 
    assign layer_2[14] = ~(layer_1[64] ^ layer_1[66]); 
    wire [1:0] far_2_2055_0;    relay_conn far_2_2055_0_a(.in(layer_1[608]), .out(far_2_2055_0[0]));    relay_conn far_2_2055_0_b(.in(layer_1[692]), .out(far_2_2055_0[1]));
    wire [1:0] far_2_2055_1;    relay_conn far_2_2055_1_a(.in(far_2_2055_0[0]), .out(far_2_2055_1[0]));    relay_conn far_2_2055_1_b(.in(far_2_2055_0[1]), .out(far_2_2055_1[1]));
    assign layer_2[15] = ~(far_2_2055_1[0] | far_2_2055_1[1]); 
    wire [1:0] far_2_2056_0;    relay_conn far_2_2056_0_a(.in(layer_1[40]), .out(far_2_2056_0[0]));    relay_conn far_2_2056_0_b(.in(layer_1[101]), .out(far_2_2056_0[1]));
    assign layer_2[16] = far_2_2056_0[1]; 
    assign layer_2[17] = layer_1[127] & layer_1[150]; 
    wire [1:0] far_2_2058_0;    relay_conn far_2_2058_0_a(.in(layer_1[383]), .out(far_2_2058_0[0]));    relay_conn far_2_2058_0_b(.in(layer_1[293]), .out(far_2_2058_0[1]));
    wire [1:0] far_2_2058_1;    relay_conn far_2_2058_1_a(.in(far_2_2058_0[0]), .out(far_2_2058_1[0]));    relay_conn far_2_2058_1_b(.in(far_2_2058_0[1]), .out(far_2_2058_1[1]));
    assign layer_2[18] = far_2_2058_1[0] | far_2_2058_1[1]; 
    wire [1:0] far_2_2059_0;    relay_conn far_2_2059_0_a(.in(layer_1[562]), .out(far_2_2059_0[0]));    relay_conn far_2_2059_0_b(.in(layer_1[596]), .out(far_2_2059_0[1]));
    assign layer_2[19] = far_2_2059_0[0] | far_2_2059_0[1]; 
    assign layer_2[20] = ~(layer_1[893] & layer_1[878]); 
    wire [1:0] far_2_2061_0;    relay_conn far_2_2061_0_a(.in(layer_1[421]), .out(far_2_2061_0[0]));    relay_conn far_2_2061_0_b(.in(layer_1[542]), .out(far_2_2061_0[1]));
    wire [1:0] far_2_2061_1;    relay_conn far_2_2061_1_a(.in(far_2_2061_0[0]), .out(far_2_2061_1[0]));    relay_conn far_2_2061_1_b(.in(far_2_2061_0[1]), .out(far_2_2061_1[1]));
    wire [1:0] far_2_2061_2;    relay_conn far_2_2061_2_a(.in(far_2_2061_1[0]), .out(far_2_2061_2[0]));    relay_conn far_2_2061_2_b(.in(far_2_2061_1[1]), .out(far_2_2061_2[1]));
    assign layer_2[21] = ~(far_2_2061_2[0] & far_2_2061_2[1]); 
    assign layer_2[22] = layer_1[234] & layer_1[215]; 
    wire [1:0] far_2_2063_0;    relay_conn far_2_2063_0_a(.in(layer_1[309]), .out(far_2_2063_0[0]));    relay_conn far_2_2063_0_b(.in(layer_1[397]), .out(far_2_2063_0[1]));
    wire [1:0] far_2_2063_1;    relay_conn far_2_2063_1_a(.in(far_2_2063_0[0]), .out(far_2_2063_1[0]));    relay_conn far_2_2063_1_b(.in(far_2_2063_0[1]), .out(far_2_2063_1[1]));
    assign layer_2[23] = ~(far_2_2063_1[0] ^ far_2_2063_1[1]); 
    wire [1:0] far_2_2064_0;    relay_conn far_2_2064_0_a(.in(layer_1[26]), .out(far_2_2064_0[0]));    relay_conn far_2_2064_0_b(.in(layer_1[132]), .out(far_2_2064_0[1]));
    wire [1:0] far_2_2064_1;    relay_conn far_2_2064_1_a(.in(far_2_2064_0[0]), .out(far_2_2064_1[0]));    relay_conn far_2_2064_1_b(.in(far_2_2064_0[1]), .out(far_2_2064_1[1]));
    wire [1:0] far_2_2064_2;    relay_conn far_2_2064_2_a(.in(far_2_2064_1[0]), .out(far_2_2064_2[0]));    relay_conn far_2_2064_2_b(.in(far_2_2064_1[1]), .out(far_2_2064_2[1]));
    assign layer_2[24] = ~far_2_2064_2[0]; 
    assign layer_2[25] = layer_1[584] & layer_1[564]; 
    wire [1:0] far_2_2066_0;    relay_conn far_2_2066_0_a(.in(layer_1[183]), .out(far_2_2066_0[0]));    relay_conn far_2_2066_0_b(.in(layer_1[283]), .out(far_2_2066_0[1]));
    wire [1:0] far_2_2066_1;    relay_conn far_2_2066_1_a(.in(far_2_2066_0[0]), .out(far_2_2066_1[0]));    relay_conn far_2_2066_1_b(.in(far_2_2066_0[1]), .out(far_2_2066_1[1]));
    wire [1:0] far_2_2066_2;    relay_conn far_2_2066_2_a(.in(far_2_2066_1[0]), .out(far_2_2066_2[0]));    relay_conn far_2_2066_2_b(.in(far_2_2066_1[1]), .out(far_2_2066_2[1]));
    assign layer_2[26] = far_2_2066_2[1] & ~far_2_2066_2[0]; 
    assign layer_2[27] = ~layer_1[423] | (layer_1[423] & layer_1[396]); 
    wire [1:0] far_2_2068_0;    relay_conn far_2_2068_0_a(.in(layer_1[932]), .out(far_2_2068_0[0]));    relay_conn far_2_2068_0_b(.in(layer_1[988]), .out(far_2_2068_0[1]));
    assign layer_2[28] = far_2_2068_0[0] | far_2_2068_0[1]; 
    wire [1:0] far_2_2069_0;    relay_conn far_2_2069_0_a(.in(layer_1[609]), .out(far_2_2069_0[0]));    relay_conn far_2_2069_0_b(.in(layer_1[481]), .out(far_2_2069_0[1]));
    wire [1:0] far_2_2069_1;    relay_conn far_2_2069_1_a(.in(far_2_2069_0[0]), .out(far_2_2069_1[0]));    relay_conn far_2_2069_1_b(.in(far_2_2069_0[1]), .out(far_2_2069_1[1]));
    wire [1:0] far_2_2069_2;    relay_conn far_2_2069_2_a(.in(far_2_2069_1[0]), .out(far_2_2069_2[0]));    relay_conn far_2_2069_2_b(.in(far_2_2069_1[1]), .out(far_2_2069_2[1]));
    wire [1:0] far_2_2069_3;    relay_conn far_2_2069_3_a(.in(far_2_2069_2[0]), .out(far_2_2069_3[0]));    relay_conn far_2_2069_3_b(.in(far_2_2069_2[1]), .out(far_2_2069_3[1]));
    assign layer_2[29] = ~far_2_2069_3[0] | (far_2_2069_3[0] & far_2_2069_3[1]); 
    wire [1:0] far_2_2070_0;    relay_conn far_2_2070_0_a(.in(layer_1[41]), .out(far_2_2070_0[0]));    relay_conn far_2_2070_0_b(.in(layer_1[166]), .out(far_2_2070_0[1]));
    wire [1:0] far_2_2070_1;    relay_conn far_2_2070_1_a(.in(far_2_2070_0[0]), .out(far_2_2070_1[0]));    relay_conn far_2_2070_1_b(.in(far_2_2070_0[1]), .out(far_2_2070_1[1]));
    wire [1:0] far_2_2070_2;    relay_conn far_2_2070_2_a(.in(far_2_2070_1[0]), .out(far_2_2070_2[0]));    relay_conn far_2_2070_2_b(.in(far_2_2070_1[1]), .out(far_2_2070_2[1]));
    assign layer_2[30] = far_2_2070_2[0] | far_2_2070_2[1]; 
    wire [1:0] far_2_2071_0;    relay_conn far_2_2071_0_a(.in(layer_1[1002]), .out(far_2_2071_0[0]));    relay_conn far_2_2071_0_b(.in(layer_1[965]), .out(far_2_2071_0[1]));
    assign layer_2[31] = ~(far_2_2071_0[0] | far_2_2071_0[1]); 
    wire [1:0] far_2_2072_0;    relay_conn far_2_2072_0_a(.in(layer_1[500]), .out(far_2_2072_0[0]));    relay_conn far_2_2072_0_b(.in(layer_1[614]), .out(far_2_2072_0[1]));
    wire [1:0] far_2_2072_1;    relay_conn far_2_2072_1_a(.in(far_2_2072_0[0]), .out(far_2_2072_1[0]));    relay_conn far_2_2072_1_b(.in(far_2_2072_0[1]), .out(far_2_2072_1[1]));
    wire [1:0] far_2_2072_2;    relay_conn far_2_2072_2_a(.in(far_2_2072_1[0]), .out(far_2_2072_2[0]));    relay_conn far_2_2072_2_b(.in(far_2_2072_1[1]), .out(far_2_2072_2[1]));
    assign layer_2[32] = ~far_2_2072_2[1] | (far_2_2072_2[0] & far_2_2072_2[1]); 
    wire [1:0] far_2_2073_0;    relay_conn far_2_2073_0_a(.in(layer_1[471]), .out(far_2_2073_0[0]));    relay_conn far_2_2073_0_b(.in(layer_1[352]), .out(far_2_2073_0[1]));
    wire [1:0] far_2_2073_1;    relay_conn far_2_2073_1_a(.in(far_2_2073_0[0]), .out(far_2_2073_1[0]));    relay_conn far_2_2073_1_b(.in(far_2_2073_0[1]), .out(far_2_2073_1[1]));
    wire [1:0] far_2_2073_2;    relay_conn far_2_2073_2_a(.in(far_2_2073_1[0]), .out(far_2_2073_2[0]));    relay_conn far_2_2073_2_b(.in(far_2_2073_1[1]), .out(far_2_2073_2[1]));
    assign layer_2[33] = far_2_2073_2[0] | far_2_2073_2[1]; 
    wire [1:0] far_2_2074_0;    relay_conn far_2_2074_0_a(.in(layer_1[646]), .out(far_2_2074_0[0]));    relay_conn far_2_2074_0_b(.in(layer_1[542]), .out(far_2_2074_0[1]));
    wire [1:0] far_2_2074_1;    relay_conn far_2_2074_1_a(.in(far_2_2074_0[0]), .out(far_2_2074_1[0]));    relay_conn far_2_2074_1_b(.in(far_2_2074_0[1]), .out(far_2_2074_1[1]));
    wire [1:0] far_2_2074_2;    relay_conn far_2_2074_2_a(.in(far_2_2074_1[0]), .out(far_2_2074_2[0]));    relay_conn far_2_2074_2_b(.in(far_2_2074_1[1]), .out(far_2_2074_2[1]));
    assign layer_2[34] = far_2_2074_2[0] & ~far_2_2074_2[1]; 
    assign layer_2[35] = ~(layer_1[138] & layer_1[159]); 
    assign layer_2[36] = ~layer_1[323] | (layer_1[321] & layer_1[323]); 
    wire [1:0] far_2_2077_0;    relay_conn far_2_2077_0_a(.in(layer_1[910]), .out(far_2_2077_0[0]));    relay_conn far_2_2077_0_b(.in(layer_1[815]), .out(far_2_2077_0[1]));
    wire [1:0] far_2_2077_1;    relay_conn far_2_2077_1_a(.in(far_2_2077_0[0]), .out(far_2_2077_1[0]));    relay_conn far_2_2077_1_b(.in(far_2_2077_0[1]), .out(far_2_2077_1[1]));
    assign layer_2[37] = far_2_2077_1[0] & ~far_2_2077_1[1]; 
    wire [1:0] far_2_2078_0;    relay_conn far_2_2078_0_a(.in(layer_1[795]), .out(far_2_2078_0[0]));    relay_conn far_2_2078_0_b(.in(layer_1[757]), .out(far_2_2078_0[1]));
    assign layer_2[38] = ~(far_2_2078_0[0] | far_2_2078_0[1]); 
    wire [1:0] far_2_2079_0;    relay_conn far_2_2079_0_a(.in(layer_1[238]), .out(far_2_2079_0[0]));    relay_conn far_2_2079_0_b(.in(layer_1[360]), .out(far_2_2079_0[1]));
    wire [1:0] far_2_2079_1;    relay_conn far_2_2079_1_a(.in(far_2_2079_0[0]), .out(far_2_2079_1[0]));    relay_conn far_2_2079_1_b(.in(far_2_2079_0[1]), .out(far_2_2079_1[1]));
    wire [1:0] far_2_2079_2;    relay_conn far_2_2079_2_a(.in(far_2_2079_1[0]), .out(far_2_2079_2[0]));    relay_conn far_2_2079_2_b(.in(far_2_2079_1[1]), .out(far_2_2079_2[1]));
    assign layer_2[39] = ~(far_2_2079_2[0] ^ far_2_2079_2[1]); 
    assign layer_2[40] = ~layer_1[962]; 
    assign layer_2[41] = ~(layer_1[2] | layer_1[12]); 
    wire [1:0] far_2_2082_0;    relay_conn far_2_2082_0_a(.in(layer_1[731]), .out(far_2_2082_0[0]));    relay_conn far_2_2082_0_b(.in(layer_1[817]), .out(far_2_2082_0[1]));
    wire [1:0] far_2_2082_1;    relay_conn far_2_2082_1_a(.in(far_2_2082_0[0]), .out(far_2_2082_1[0]));    relay_conn far_2_2082_1_b(.in(far_2_2082_0[1]), .out(far_2_2082_1[1]));
    assign layer_2[42] = ~(far_2_2082_1[0] ^ far_2_2082_1[1]); 
    wire [1:0] far_2_2083_0;    relay_conn far_2_2083_0_a(.in(layer_1[309]), .out(far_2_2083_0[0]));    relay_conn far_2_2083_0_b(.in(layer_1[208]), .out(far_2_2083_0[1]));
    wire [1:0] far_2_2083_1;    relay_conn far_2_2083_1_a(.in(far_2_2083_0[0]), .out(far_2_2083_1[0]));    relay_conn far_2_2083_1_b(.in(far_2_2083_0[1]), .out(far_2_2083_1[1]));
    wire [1:0] far_2_2083_2;    relay_conn far_2_2083_2_a(.in(far_2_2083_1[0]), .out(far_2_2083_2[0]));    relay_conn far_2_2083_2_b(.in(far_2_2083_1[1]), .out(far_2_2083_2[1]));
    assign layer_2[43] = far_2_2083_2[0] & ~far_2_2083_2[1]; 
    assign layer_2[44] = layer_1[355] | layer_1[363]; 
    wire [1:0] far_2_2085_0;    relay_conn far_2_2085_0_a(.in(layer_1[12]), .out(far_2_2085_0[0]));    relay_conn far_2_2085_0_b(.in(layer_1[54]), .out(far_2_2085_0[1]));
    assign layer_2[45] = ~far_2_2085_0[0] | (far_2_2085_0[0] & far_2_2085_0[1]); 
    wire [1:0] far_2_2086_0;    relay_conn far_2_2086_0_a(.in(layer_1[955]), .out(far_2_2086_0[0]));    relay_conn far_2_2086_0_b(.in(layer_1[900]), .out(far_2_2086_0[1]));
    assign layer_2[46] = ~(far_2_2086_0[0] ^ far_2_2086_0[1]); 
    wire [1:0] far_2_2087_0;    relay_conn far_2_2087_0_a(.in(layer_1[219]), .out(far_2_2087_0[0]));    relay_conn far_2_2087_0_b(.in(layer_1[313]), .out(far_2_2087_0[1]));
    wire [1:0] far_2_2087_1;    relay_conn far_2_2087_1_a(.in(far_2_2087_0[0]), .out(far_2_2087_1[0]));    relay_conn far_2_2087_1_b(.in(far_2_2087_0[1]), .out(far_2_2087_1[1]));
    assign layer_2[47] = ~far_2_2087_1[0]; 
    wire [1:0] far_2_2088_0;    relay_conn far_2_2088_0_a(.in(layer_1[644]), .out(far_2_2088_0[0]));    relay_conn far_2_2088_0_b(.in(layer_1[525]), .out(far_2_2088_0[1]));
    wire [1:0] far_2_2088_1;    relay_conn far_2_2088_1_a(.in(far_2_2088_0[0]), .out(far_2_2088_1[0]));    relay_conn far_2_2088_1_b(.in(far_2_2088_0[1]), .out(far_2_2088_1[1]));
    wire [1:0] far_2_2088_2;    relay_conn far_2_2088_2_a(.in(far_2_2088_1[0]), .out(far_2_2088_2[0]));    relay_conn far_2_2088_2_b(.in(far_2_2088_1[1]), .out(far_2_2088_2[1]));
    assign layer_2[48] = far_2_2088_2[0] & ~far_2_2088_2[1]; 
    wire [1:0] far_2_2089_0;    relay_conn far_2_2089_0_a(.in(layer_1[889]), .out(far_2_2089_0[0]));    relay_conn far_2_2089_0_b(.in(layer_1[951]), .out(far_2_2089_0[1]));
    assign layer_2[49] = ~far_2_2089_0[0] | (far_2_2089_0[0] & far_2_2089_0[1]); 
    wire [1:0] far_2_2090_0;    relay_conn far_2_2090_0_a(.in(layer_1[502]), .out(far_2_2090_0[0]));    relay_conn far_2_2090_0_b(.in(layer_1[467]), .out(far_2_2090_0[1]));
    assign layer_2[50] = ~(far_2_2090_0[0] ^ far_2_2090_0[1]); 
    wire [1:0] far_2_2091_0;    relay_conn far_2_2091_0_a(.in(layer_1[338]), .out(far_2_2091_0[0]));    relay_conn far_2_2091_0_b(.in(layer_1[437]), .out(far_2_2091_0[1]));
    wire [1:0] far_2_2091_1;    relay_conn far_2_2091_1_a(.in(far_2_2091_0[0]), .out(far_2_2091_1[0]));    relay_conn far_2_2091_1_b(.in(far_2_2091_0[1]), .out(far_2_2091_1[1]));
    wire [1:0] far_2_2091_2;    relay_conn far_2_2091_2_a(.in(far_2_2091_1[0]), .out(far_2_2091_2[0]));    relay_conn far_2_2091_2_b(.in(far_2_2091_1[1]), .out(far_2_2091_2[1]));
    assign layer_2[51] = ~far_2_2091_2[1] | (far_2_2091_2[0] & far_2_2091_2[1]); 
    wire [1:0] far_2_2092_0;    relay_conn far_2_2092_0_a(.in(layer_1[182]), .out(far_2_2092_0[0]));    relay_conn far_2_2092_0_b(.in(layer_1[309]), .out(far_2_2092_0[1]));
    wire [1:0] far_2_2092_1;    relay_conn far_2_2092_1_a(.in(far_2_2092_0[0]), .out(far_2_2092_1[0]));    relay_conn far_2_2092_1_b(.in(far_2_2092_0[1]), .out(far_2_2092_1[1]));
    wire [1:0] far_2_2092_2;    relay_conn far_2_2092_2_a(.in(far_2_2092_1[0]), .out(far_2_2092_2[0]));    relay_conn far_2_2092_2_b(.in(far_2_2092_1[1]), .out(far_2_2092_2[1]));
    assign layer_2[52] = far_2_2092_2[0] | far_2_2092_2[1]; 
    assign layer_2[53] = ~(layer_1[95] | layer_1[92]); 
    wire [1:0] far_2_2094_0;    relay_conn far_2_2094_0_a(.in(layer_1[786]), .out(far_2_2094_0[0]));    relay_conn far_2_2094_0_b(.in(layer_1[716]), .out(far_2_2094_0[1]));
    wire [1:0] far_2_2094_1;    relay_conn far_2_2094_1_a(.in(far_2_2094_0[0]), .out(far_2_2094_1[0]));    relay_conn far_2_2094_1_b(.in(far_2_2094_0[1]), .out(far_2_2094_1[1]));
    assign layer_2[54] = far_2_2094_1[1]; 
    assign layer_2[55] = layer_1[862]; 
    wire [1:0] far_2_2096_0;    relay_conn far_2_2096_0_a(.in(layer_1[476]), .out(far_2_2096_0[0]));    relay_conn far_2_2096_0_b(.in(layer_1[426]), .out(far_2_2096_0[1]));
    assign layer_2[56] = ~far_2_2096_0[1] | (far_2_2096_0[0] & far_2_2096_0[1]); 
    wire [1:0] far_2_2097_0;    relay_conn far_2_2097_0_a(.in(layer_1[333]), .out(far_2_2097_0[0]));    relay_conn far_2_2097_0_b(.in(layer_1[408]), .out(far_2_2097_0[1]));
    wire [1:0] far_2_2097_1;    relay_conn far_2_2097_1_a(.in(far_2_2097_0[0]), .out(far_2_2097_1[0]));    relay_conn far_2_2097_1_b(.in(far_2_2097_0[1]), .out(far_2_2097_1[1]));
    assign layer_2[57] = ~far_2_2097_1[0]; 
    wire [1:0] far_2_2098_0;    relay_conn far_2_2098_0_a(.in(layer_1[613]), .out(far_2_2098_0[0]));    relay_conn far_2_2098_0_b(.in(layer_1[711]), .out(far_2_2098_0[1]));
    wire [1:0] far_2_2098_1;    relay_conn far_2_2098_1_a(.in(far_2_2098_0[0]), .out(far_2_2098_1[0]));    relay_conn far_2_2098_1_b(.in(far_2_2098_0[1]), .out(far_2_2098_1[1]));
    wire [1:0] far_2_2098_2;    relay_conn far_2_2098_2_a(.in(far_2_2098_1[0]), .out(far_2_2098_2[0]));    relay_conn far_2_2098_2_b(.in(far_2_2098_1[1]), .out(far_2_2098_2[1]));
    assign layer_2[58] = ~far_2_2098_2[0] | (far_2_2098_2[0] & far_2_2098_2[1]); 
    wire [1:0] far_2_2099_0;    relay_conn far_2_2099_0_a(.in(layer_1[130]), .out(far_2_2099_0[0]));    relay_conn far_2_2099_0_b(.in(layer_1[165]), .out(far_2_2099_0[1]));
    assign layer_2[59] = ~far_2_2099_0[0] | (far_2_2099_0[0] & far_2_2099_0[1]); 
    wire [1:0] far_2_2100_0;    relay_conn far_2_2100_0_a(.in(layer_1[743]), .out(far_2_2100_0[0]));    relay_conn far_2_2100_0_b(.in(layer_1[646]), .out(far_2_2100_0[1]));
    wire [1:0] far_2_2100_1;    relay_conn far_2_2100_1_a(.in(far_2_2100_0[0]), .out(far_2_2100_1[0]));    relay_conn far_2_2100_1_b(.in(far_2_2100_0[1]), .out(far_2_2100_1[1]));
    wire [1:0] far_2_2100_2;    relay_conn far_2_2100_2_a(.in(far_2_2100_1[0]), .out(far_2_2100_2[0]));    relay_conn far_2_2100_2_b(.in(far_2_2100_1[1]), .out(far_2_2100_2[1]));
    assign layer_2[60] = far_2_2100_2[0]; 
    wire [1:0] far_2_2101_0;    relay_conn far_2_2101_0_a(.in(layer_1[690]), .out(far_2_2101_0[0]));    relay_conn far_2_2101_0_b(.in(layer_1[582]), .out(far_2_2101_0[1]));
    wire [1:0] far_2_2101_1;    relay_conn far_2_2101_1_a(.in(far_2_2101_0[0]), .out(far_2_2101_1[0]));    relay_conn far_2_2101_1_b(.in(far_2_2101_0[1]), .out(far_2_2101_1[1]));
    wire [1:0] far_2_2101_2;    relay_conn far_2_2101_2_a(.in(far_2_2101_1[0]), .out(far_2_2101_2[0]));    relay_conn far_2_2101_2_b(.in(far_2_2101_1[1]), .out(far_2_2101_2[1]));
    assign layer_2[61] = far_2_2101_2[0] & ~far_2_2101_2[1]; 
    wire [1:0] far_2_2102_0;    relay_conn far_2_2102_0_a(.in(layer_1[98]), .out(far_2_2102_0[0]));    relay_conn far_2_2102_0_b(.in(layer_1[22]), .out(far_2_2102_0[1]));
    wire [1:0] far_2_2102_1;    relay_conn far_2_2102_1_a(.in(far_2_2102_0[0]), .out(far_2_2102_1[0]));    relay_conn far_2_2102_1_b(.in(far_2_2102_0[1]), .out(far_2_2102_1[1]));
    assign layer_2[62] = far_2_2102_1[0] | far_2_2102_1[1]; 
    wire [1:0] far_2_2103_0;    relay_conn far_2_2103_0_a(.in(layer_1[727]), .out(far_2_2103_0[0]));    relay_conn far_2_2103_0_b(.in(layer_1[622]), .out(far_2_2103_0[1]));
    wire [1:0] far_2_2103_1;    relay_conn far_2_2103_1_a(.in(far_2_2103_0[0]), .out(far_2_2103_1[0]));    relay_conn far_2_2103_1_b(.in(far_2_2103_0[1]), .out(far_2_2103_1[1]));
    wire [1:0] far_2_2103_2;    relay_conn far_2_2103_2_a(.in(far_2_2103_1[0]), .out(far_2_2103_2[0]));    relay_conn far_2_2103_2_b(.in(far_2_2103_1[1]), .out(far_2_2103_2[1]));
    assign layer_2[63] = ~far_2_2103_2[0]; 
    wire [1:0] far_2_2104_0;    relay_conn far_2_2104_0_a(.in(layer_1[506]), .out(far_2_2104_0[0]));    relay_conn far_2_2104_0_b(.in(layer_1[391]), .out(far_2_2104_0[1]));
    wire [1:0] far_2_2104_1;    relay_conn far_2_2104_1_a(.in(far_2_2104_0[0]), .out(far_2_2104_1[0]));    relay_conn far_2_2104_1_b(.in(far_2_2104_0[1]), .out(far_2_2104_1[1]));
    wire [1:0] far_2_2104_2;    relay_conn far_2_2104_2_a(.in(far_2_2104_1[0]), .out(far_2_2104_2[0]));    relay_conn far_2_2104_2_b(.in(far_2_2104_1[1]), .out(far_2_2104_2[1]));
    assign layer_2[64] = far_2_2104_2[1] & ~far_2_2104_2[0]; 
    wire [1:0] far_2_2105_0;    relay_conn far_2_2105_0_a(.in(layer_1[0]), .out(far_2_2105_0[0]));    relay_conn far_2_2105_0_b(.in(layer_1[93]), .out(far_2_2105_0[1]));
    wire [1:0] far_2_2105_1;    relay_conn far_2_2105_1_a(.in(far_2_2105_0[0]), .out(far_2_2105_1[0]));    relay_conn far_2_2105_1_b(.in(far_2_2105_0[1]), .out(far_2_2105_1[1]));
    assign layer_2[65] = far_2_2105_1[1] & ~far_2_2105_1[0]; 
    wire [1:0] far_2_2106_0;    relay_conn far_2_2106_0_a(.in(layer_1[662]), .out(far_2_2106_0[0]));    relay_conn far_2_2106_0_b(.in(layer_1[763]), .out(far_2_2106_0[1]));
    wire [1:0] far_2_2106_1;    relay_conn far_2_2106_1_a(.in(far_2_2106_0[0]), .out(far_2_2106_1[0]));    relay_conn far_2_2106_1_b(.in(far_2_2106_0[1]), .out(far_2_2106_1[1]));
    wire [1:0] far_2_2106_2;    relay_conn far_2_2106_2_a(.in(far_2_2106_1[0]), .out(far_2_2106_2[0]));    relay_conn far_2_2106_2_b(.in(far_2_2106_1[1]), .out(far_2_2106_2[1]));
    assign layer_2[66] = ~(far_2_2106_2[0] ^ far_2_2106_2[1]); 
    assign layer_2[67] = ~(layer_1[284] & layer_1[256]); 
    wire [1:0] far_2_2108_0;    relay_conn far_2_2108_0_a(.in(layer_1[917]), .out(far_2_2108_0[0]));    relay_conn far_2_2108_0_b(.in(layer_1[954]), .out(far_2_2108_0[1]));
    assign layer_2[68] = ~(far_2_2108_0[0] ^ far_2_2108_0[1]); 
    wire [1:0] far_2_2109_0;    relay_conn far_2_2109_0_a(.in(layer_1[234]), .out(far_2_2109_0[0]));    relay_conn far_2_2109_0_b(.in(layer_1[278]), .out(far_2_2109_0[1]));
    assign layer_2[69] = ~(far_2_2109_0[0] & far_2_2109_0[1]); 
    assign layer_2[70] = ~layer_1[71]; 
    wire [1:0] far_2_2111_0;    relay_conn far_2_2111_0_a(.in(layer_1[932]), .out(far_2_2111_0[0]));    relay_conn far_2_2111_0_b(.in(layer_1[850]), .out(far_2_2111_0[1]));
    wire [1:0] far_2_2111_1;    relay_conn far_2_2111_1_a(.in(far_2_2111_0[0]), .out(far_2_2111_1[0]));    relay_conn far_2_2111_1_b(.in(far_2_2111_0[1]), .out(far_2_2111_1[1]));
    assign layer_2[71] = far_2_2111_1[0] & ~far_2_2111_1[1]; 
    wire [1:0] far_2_2112_0;    relay_conn far_2_2112_0_a(.in(layer_1[348]), .out(far_2_2112_0[0]));    relay_conn far_2_2112_0_b(.in(layer_1[311]), .out(far_2_2112_0[1]));
    assign layer_2[72] = far_2_2112_0[0] & far_2_2112_0[1]; 
    wire [1:0] far_2_2113_0;    relay_conn far_2_2113_0_a(.in(layer_1[505]), .out(far_2_2113_0[0]));    relay_conn far_2_2113_0_b(.in(layer_1[537]), .out(far_2_2113_0[1]));
    assign layer_2[73] = far_2_2113_0[0] ^ far_2_2113_0[1]; 
    wire [1:0] far_2_2114_0;    relay_conn far_2_2114_0_a(.in(layer_1[338]), .out(far_2_2114_0[0]));    relay_conn far_2_2114_0_b(.in(layer_1[393]), .out(far_2_2114_0[1]));
    assign layer_2[74] = ~far_2_2114_0[0] | (far_2_2114_0[0] & far_2_2114_0[1]); 
    wire [1:0] far_2_2115_0;    relay_conn far_2_2115_0_a(.in(layer_1[688]), .out(far_2_2115_0[0]));    relay_conn far_2_2115_0_b(.in(layer_1[795]), .out(far_2_2115_0[1]));
    wire [1:0] far_2_2115_1;    relay_conn far_2_2115_1_a(.in(far_2_2115_0[0]), .out(far_2_2115_1[0]));    relay_conn far_2_2115_1_b(.in(far_2_2115_0[1]), .out(far_2_2115_1[1]));
    wire [1:0] far_2_2115_2;    relay_conn far_2_2115_2_a(.in(far_2_2115_1[0]), .out(far_2_2115_2[0]));    relay_conn far_2_2115_2_b(.in(far_2_2115_1[1]), .out(far_2_2115_2[1]));
    assign layer_2[75] = far_2_2115_2[0]; 
    wire [1:0] far_2_2116_0;    relay_conn far_2_2116_0_a(.in(layer_1[220]), .out(far_2_2116_0[0]));    relay_conn far_2_2116_0_b(.in(layer_1[118]), .out(far_2_2116_0[1]));
    wire [1:0] far_2_2116_1;    relay_conn far_2_2116_1_a(.in(far_2_2116_0[0]), .out(far_2_2116_1[0]));    relay_conn far_2_2116_1_b(.in(far_2_2116_0[1]), .out(far_2_2116_1[1]));
    wire [1:0] far_2_2116_2;    relay_conn far_2_2116_2_a(.in(far_2_2116_1[0]), .out(far_2_2116_2[0]));    relay_conn far_2_2116_2_b(.in(far_2_2116_1[1]), .out(far_2_2116_2[1]));
    assign layer_2[76] = far_2_2116_2[0] & ~far_2_2116_2[1]; 
    assign layer_2[77] = layer_1[323] | layer_1[316]; 
    wire [1:0] far_2_2118_0;    relay_conn far_2_2118_0_a(.in(layer_1[941]), .out(far_2_2118_0[0]));    relay_conn far_2_2118_0_b(.in(layer_1[994]), .out(far_2_2118_0[1]));
    assign layer_2[78] = far_2_2118_0[0] | far_2_2118_0[1]; 
    wire [1:0] far_2_2119_0;    relay_conn far_2_2119_0_a(.in(layer_1[521]), .out(far_2_2119_0[0]));    relay_conn far_2_2119_0_b(.in(layer_1[408]), .out(far_2_2119_0[1]));
    wire [1:0] far_2_2119_1;    relay_conn far_2_2119_1_a(.in(far_2_2119_0[0]), .out(far_2_2119_1[0]));    relay_conn far_2_2119_1_b(.in(far_2_2119_0[1]), .out(far_2_2119_1[1]));
    wire [1:0] far_2_2119_2;    relay_conn far_2_2119_2_a(.in(far_2_2119_1[0]), .out(far_2_2119_2[0]));    relay_conn far_2_2119_2_b(.in(far_2_2119_1[1]), .out(far_2_2119_2[1]));
    assign layer_2[79] = far_2_2119_2[0] | far_2_2119_2[1]; 
    wire [1:0] far_2_2120_0;    relay_conn far_2_2120_0_a(.in(layer_1[288]), .out(far_2_2120_0[0]));    relay_conn far_2_2120_0_b(.in(layer_1[329]), .out(far_2_2120_0[1]));
    assign layer_2[80] = far_2_2120_0[0] & ~far_2_2120_0[1]; 
    wire [1:0] far_2_2121_0;    relay_conn far_2_2121_0_a(.in(layer_1[537]), .out(far_2_2121_0[0]));    relay_conn far_2_2121_0_b(.in(layer_1[630]), .out(far_2_2121_0[1]));
    wire [1:0] far_2_2121_1;    relay_conn far_2_2121_1_a(.in(far_2_2121_0[0]), .out(far_2_2121_1[0]));    relay_conn far_2_2121_1_b(.in(far_2_2121_0[1]), .out(far_2_2121_1[1]));
    assign layer_2[81] = far_2_2121_1[0] & ~far_2_2121_1[1]; 
    wire [1:0] far_2_2122_0;    relay_conn far_2_2122_0_a(.in(layer_1[137]), .out(far_2_2122_0[0]));    relay_conn far_2_2122_0_b(.in(layer_1[98]), .out(far_2_2122_0[1]));
    assign layer_2[82] = ~far_2_2122_0[0]; 
    assign layer_2[83] = ~(layer_1[416] | layer_1[432]); 
    wire [1:0] far_2_2124_0;    relay_conn far_2_2124_0_a(.in(layer_1[835]), .out(far_2_2124_0[0]));    relay_conn far_2_2124_0_b(.in(layer_1[717]), .out(far_2_2124_0[1]));
    wire [1:0] far_2_2124_1;    relay_conn far_2_2124_1_a(.in(far_2_2124_0[0]), .out(far_2_2124_1[0]));    relay_conn far_2_2124_1_b(.in(far_2_2124_0[1]), .out(far_2_2124_1[1]));
    wire [1:0] far_2_2124_2;    relay_conn far_2_2124_2_a(.in(far_2_2124_1[0]), .out(far_2_2124_2[0]));    relay_conn far_2_2124_2_b(.in(far_2_2124_1[1]), .out(far_2_2124_2[1]));
    assign layer_2[84] = ~(far_2_2124_2[0] & far_2_2124_2[1]); 
    wire [1:0] far_2_2125_0;    relay_conn far_2_2125_0_a(.in(layer_1[701]), .out(far_2_2125_0[0]));    relay_conn far_2_2125_0_b(.in(layer_1[789]), .out(far_2_2125_0[1]));
    wire [1:0] far_2_2125_1;    relay_conn far_2_2125_1_a(.in(far_2_2125_0[0]), .out(far_2_2125_1[0]));    relay_conn far_2_2125_1_b(.in(far_2_2125_0[1]), .out(far_2_2125_1[1]));
    assign layer_2[85] = far_2_2125_1[0]; 
    wire [1:0] far_2_2126_0;    relay_conn far_2_2126_0_a(.in(layer_1[692]), .out(far_2_2126_0[0]));    relay_conn far_2_2126_0_b(.in(layer_1[574]), .out(far_2_2126_0[1]));
    wire [1:0] far_2_2126_1;    relay_conn far_2_2126_1_a(.in(far_2_2126_0[0]), .out(far_2_2126_1[0]));    relay_conn far_2_2126_1_b(.in(far_2_2126_0[1]), .out(far_2_2126_1[1]));
    wire [1:0] far_2_2126_2;    relay_conn far_2_2126_2_a(.in(far_2_2126_1[0]), .out(far_2_2126_2[0]));    relay_conn far_2_2126_2_b(.in(far_2_2126_1[1]), .out(far_2_2126_2[1]));
    assign layer_2[86] = far_2_2126_2[1] & ~far_2_2126_2[0]; 
    wire [1:0] far_2_2127_0;    relay_conn far_2_2127_0_a(.in(layer_1[443]), .out(far_2_2127_0[0]));    relay_conn far_2_2127_0_b(.in(layer_1[364]), .out(far_2_2127_0[1]));
    wire [1:0] far_2_2127_1;    relay_conn far_2_2127_1_a(.in(far_2_2127_0[0]), .out(far_2_2127_1[0]));    relay_conn far_2_2127_1_b(.in(far_2_2127_0[1]), .out(far_2_2127_1[1]));
    assign layer_2[87] = far_2_2127_1[0] & ~far_2_2127_1[1]; 
    wire [1:0] far_2_2128_0;    relay_conn far_2_2128_0_a(.in(layer_1[401]), .out(far_2_2128_0[0]));    relay_conn far_2_2128_0_b(.in(layer_1[446]), .out(far_2_2128_0[1]));
    assign layer_2[88] = ~(far_2_2128_0[0] ^ far_2_2128_0[1]); 
    wire [1:0] far_2_2129_0;    relay_conn far_2_2129_0_a(.in(layer_1[33]), .out(far_2_2129_0[0]));    relay_conn far_2_2129_0_b(.in(layer_1[151]), .out(far_2_2129_0[1]));
    wire [1:0] far_2_2129_1;    relay_conn far_2_2129_1_a(.in(far_2_2129_0[0]), .out(far_2_2129_1[0]));    relay_conn far_2_2129_1_b(.in(far_2_2129_0[1]), .out(far_2_2129_1[1]));
    wire [1:0] far_2_2129_2;    relay_conn far_2_2129_2_a(.in(far_2_2129_1[0]), .out(far_2_2129_2[0]));    relay_conn far_2_2129_2_b(.in(far_2_2129_1[1]), .out(far_2_2129_2[1]));
    assign layer_2[89] = ~far_2_2129_2[1] | (far_2_2129_2[0] & far_2_2129_2[1]); 
    wire [1:0] far_2_2130_0;    relay_conn far_2_2130_0_a(.in(layer_1[374]), .out(far_2_2130_0[0]));    relay_conn far_2_2130_0_b(.in(layer_1[481]), .out(far_2_2130_0[1]));
    wire [1:0] far_2_2130_1;    relay_conn far_2_2130_1_a(.in(far_2_2130_0[0]), .out(far_2_2130_1[0]));    relay_conn far_2_2130_1_b(.in(far_2_2130_0[1]), .out(far_2_2130_1[1]));
    wire [1:0] far_2_2130_2;    relay_conn far_2_2130_2_a(.in(far_2_2130_1[0]), .out(far_2_2130_2[0]));    relay_conn far_2_2130_2_b(.in(far_2_2130_1[1]), .out(far_2_2130_2[1]));
    assign layer_2[90] = ~far_2_2130_2[1]; 
    wire [1:0] far_2_2131_0;    relay_conn far_2_2131_0_a(.in(layer_1[373]), .out(far_2_2131_0[0]));    relay_conn far_2_2131_0_b(.in(layer_1[284]), .out(far_2_2131_0[1]));
    wire [1:0] far_2_2131_1;    relay_conn far_2_2131_1_a(.in(far_2_2131_0[0]), .out(far_2_2131_1[0]));    relay_conn far_2_2131_1_b(.in(far_2_2131_0[1]), .out(far_2_2131_1[1]));
    assign layer_2[91] = far_2_2131_1[0] & ~far_2_2131_1[1]; 
    wire [1:0] far_2_2132_0;    relay_conn far_2_2132_0_a(.in(layer_1[814]), .out(far_2_2132_0[0]));    relay_conn far_2_2132_0_b(.in(layer_1[865]), .out(far_2_2132_0[1]));
    assign layer_2[92] = far_2_2132_0[1] & ~far_2_2132_0[0]; 
    assign layer_2[93] = layer_1[40]; 
    assign layer_2[94] = layer_1[812] & layer_1[796]; 
    wire [1:0] far_2_2135_0;    relay_conn far_2_2135_0_a(.in(layer_1[12]), .out(far_2_2135_0[0]));    relay_conn far_2_2135_0_b(.in(layer_1[65]), .out(far_2_2135_0[1]));
    assign layer_2[95] = far_2_2135_0[1] & ~far_2_2135_0[0]; 
    wire [1:0] far_2_2136_0;    relay_conn far_2_2136_0_a(.in(layer_1[450]), .out(far_2_2136_0[0]));    relay_conn far_2_2136_0_b(.in(layer_1[417]), .out(far_2_2136_0[1]));
    assign layer_2[96] = far_2_2136_0[1] & ~far_2_2136_0[0]; 
    wire [1:0] far_2_2137_0;    relay_conn far_2_2137_0_a(.in(layer_1[687]), .out(far_2_2137_0[0]));    relay_conn far_2_2137_0_b(.in(layer_1[561]), .out(far_2_2137_0[1]));
    wire [1:0] far_2_2137_1;    relay_conn far_2_2137_1_a(.in(far_2_2137_0[0]), .out(far_2_2137_1[0]));    relay_conn far_2_2137_1_b(.in(far_2_2137_0[1]), .out(far_2_2137_1[1]));
    wire [1:0] far_2_2137_2;    relay_conn far_2_2137_2_a(.in(far_2_2137_1[0]), .out(far_2_2137_2[0]));    relay_conn far_2_2137_2_b(.in(far_2_2137_1[1]), .out(far_2_2137_2[1]));
    assign layer_2[97] = ~(far_2_2137_2[0] & far_2_2137_2[1]); 
    wire [1:0] far_2_2138_0;    relay_conn far_2_2138_0_a(.in(layer_1[521]), .out(far_2_2138_0[0]));    relay_conn far_2_2138_0_b(.in(layer_1[559]), .out(far_2_2138_0[1]));
    assign layer_2[98] = ~(far_2_2138_0[0] & far_2_2138_0[1]); 
    wire [1:0] far_2_2139_0;    relay_conn far_2_2139_0_a(.in(layer_1[447]), .out(far_2_2139_0[0]));    relay_conn far_2_2139_0_b(.in(layer_1[505]), .out(far_2_2139_0[1]));
    assign layer_2[99] = ~far_2_2139_0[0]; 
    wire [1:0] far_2_2140_0;    relay_conn far_2_2140_0_a(.in(layer_1[66]), .out(far_2_2140_0[0]));    relay_conn far_2_2140_0_b(.in(layer_1[102]), .out(far_2_2140_0[1]));
    assign layer_2[100] = far_2_2140_0[0] & far_2_2140_0[1]; 
    wire [1:0] far_2_2141_0;    relay_conn far_2_2141_0_a(.in(layer_1[910]), .out(far_2_2141_0[0]));    relay_conn far_2_2141_0_b(.in(layer_1[814]), .out(far_2_2141_0[1]));
    wire [1:0] far_2_2141_1;    relay_conn far_2_2141_1_a(.in(far_2_2141_0[0]), .out(far_2_2141_1[0]));    relay_conn far_2_2141_1_b(.in(far_2_2141_0[1]), .out(far_2_2141_1[1]));
    wire [1:0] far_2_2141_2;    relay_conn far_2_2141_2_a(.in(far_2_2141_1[0]), .out(far_2_2141_2[0]));    relay_conn far_2_2141_2_b(.in(far_2_2141_1[1]), .out(far_2_2141_2[1]));
    assign layer_2[101] = far_2_2141_2[0] | far_2_2141_2[1]; 
    wire [1:0] far_2_2142_0;    relay_conn far_2_2142_0_a(.in(layer_1[765]), .out(far_2_2142_0[0]));    relay_conn far_2_2142_0_b(.in(layer_1[669]), .out(far_2_2142_0[1]));
    wire [1:0] far_2_2142_1;    relay_conn far_2_2142_1_a(.in(far_2_2142_0[0]), .out(far_2_2142_1[0]));    relay_conn far_2_2142_1_b(.in(far_2_2142_0[1]), .out(far_2_2142_1[1]));
    wire [1:0] far_2_2142_2;    relay_conn far_2_2142_2_a(.in(far_2_2142_1[0]), .out(far_2_2142_2[0]));    relay_conn far_2_2142_2_b(.in(far_2_2142_1[1]), .out(far_2_2142_2[1]));
    assign layer_2[102] = far_2_2142_2[0] & far_2_2142_2[1]; 
    wire [1:0] far_2_2143_0;    relay_conn far_2_2143_0_a(.in(layer_1[875]), .out(far_2_2143_0[0]));    relay_conn far_2_2143_0_b(.in(layer_1[998]), .out(far_2_2143_0[1]));
    wire [1:0] far_2_2143_1;    relay_conn far_2_2143_1_a(.in(far_2_2143_0[0]), .out(far_2_2143_1[0]));    relay_conn far_2_2143_1_b(.in(far_2_2143_0[1]), .out(far_2_2143_1[1]));
    wire [1:0] far_2_2143_2;    relay_conn far_2_2143_2_a(.in(far_2_2143_1[0]), .out(far_2_2143_2[0]));    relay_conn far_2_2143_2_b(.in(far_2_2143_1[1]), .out(far_2_2143_2[1]));
    assign layer_2[103] = ~far_2_2143_2[0]; 
    wire [1:0] far_2_2144_0;    relay_conn far_2_2144_0_a(.in(layer_1[341]), .out(far_2_2144_0[0]));    relay_conn far_2_2144_0_b(.in(layer_1[288]), .out(far_2_2144_0[1]));
    assign layer_2[104] = ~far_2_2144_0[1] | (far_2_2144_0[0] & far_2_2144_0[1]); 
    wire [1:0] far_2_2145_0;    relay_conn far_2_2145_0_a(.in(layer_1[724]), .out(far_2_2145_0[0]));    relay_conn far_2_2145_0_b(.in(layer_1[656]), .out(far_2_2145_0[1]));
    wire [1:0] far_2_2145_1;    relay_conn far_2_2145_1_a(.in(far_2_2145_0[0]), .out(far_2_2145_1[0]));    relay_conn far_2_2145_1_b(.in(far_2_2145_0[1]), .out(far_2_2145_1[1]));
    assign layer_2[105] = ~far_2_2145_1[0] | (far_2_2145_1[0] & far_2_2145_1[1]); 
    wire [1:0] far_2_2146_0;    relay_conn far_2_2146_0_a(.in(layer_1[784]), .out(far_2_2146_0[0]));    relay_conn far_2_2146_0_b(.in(layer_1[671]), .out(far_2_2146_0[1]));
    wire [1:0] far_2_2146_1;    relay_conn far_2_2146_1_a(.in(far_2_2146_0[0]), .out(far_2_2146_1[0]));    relay_conn far_2_2146_1_b(.in(far_2_2146_0[1]), .out(far_2_2146_1[1]));
    wire [1:0] far_2_2146_2;    relay_conn far_2_2146_2_a(.in(far_2_2146_1[0]), .out(far_2_2146_2[0]));    relay_conn far_2_2146_2_b(.in(far_2_2146_1[1]), .out(far_2_2146_2[1]));
    assign layer_2[106] = far_2_2146_2[0] | far_2_2146_2[1]; 
    wire [1:0] far_2_2147_0;    relay_conn far_2_2147_0_a(.in(layer_1[1000]), .out(far_2_2147_0[0]));    relay_conn far_2_2147_0_b(.in(layer_1[896]), .out(far_2_2147_0[1]));
    wire [1:0] far_2_2147_1;    relay_conn far_2_2147_1_a(.in(far_2_2147_0[0]), .out(far_2_2147_1[0]));    relay_conn far_2_2147_1_b(.in(far_2_2147_0[1]), .out(far_2_2147_1[1]));
    wire [1:0] far_2_2147_2;    relay_conn far_2_2147_2_a(.in(far_2_2147_1[0]), .out(far_2_2147_2[0]));    relay_conn far_2_2147_2_b(.in(far_2_2147_1[1]), .out(far_2_2147_2[1]));
    assign layer_2[107] = far_2_2147_2[1] & ~far_2_2147_2[0]; 
    wire [1:0] far_2_2148_0;    relay_conn far_2_2148_0_a(.in(layer_1[308]), .out(far_2_2148_0[0]));    relay_conn far_2_2148_0_b(.in(layer_1[429]), .out(far_2_2148_0[1]));
    wire [1:0] far_2_2148_1;    relay_conn far_2_2148_1_a(.in(far_2_2148_0[0]), .out(far_2_2148_1[0]));    relay_conn far_2_2148_1_b(.in(far_2_2148_0[1]), .out(far_2_2148_1[1]));
    wire [1:0] far_2_2148_2;    relay_conn far_2_2148_2_a(.in(far_2_2148_1[0]), .out(far_2_2148_2[0]));    relay_conn far_2_2148_2_b(.in(far_2_2148_1[1]), .out(far_2_2148_2[1]));
    assign layer_2[108] = far_2_2148_2[0] & ~far_2_2148_2[1]; 
    wire [1:0] far_2_2149_0;    relay_conn far_2_2149_0_a(.in(layer_1[796]), .out(far_2_2149_0[0]));    relay_conn far_2_2149_0_b(.in(layer_1[734]), .out(far_2_2149_0[1]));
    assign layer_2[109] = far_2_2149_0[1] & ~far_2_2149_0[0]; 
    assign layer_2[110] = ~layer_1[169] | (layer_1[171] & layer_1[169]); 
    wire [1:0] far_2_2151_0;    relay_conn far_2_2151_0_a(.in(layer_1[776]), .out(far_2_2151_0[0]));    relay_conn far_2_2151_0_b(.in(layer_1[732]), .out(far_2_2151_0[1]));
    assign layer_2[111] = far_2_2151_0[1] & ~far_2_2151_0[0]; 
    wire [1:0] far_2_2152_0;    relay_conn far_2_2152_0_a(.in(layer_1[707]), .out(far_2_2152_0[0]));    relay_conn far_2_2152_0_b(.in(layer_1[657]), .out(far_2_2152_0[1]));
    assign layer_2[112] = ~far_2_2152_0[0] | (far_2_2152_0[0] & far_2_2152_0[1]); 
    assign layer_2[113] = ~(layer_1[920] | layer_1[919]); 
    wire [1:0] far_2_2154_0;    relay_conn far_2_2154_0_a(.in(layer_1[363]), .out(far_2_2154_0[0]));    relay_conn far_2_2154_0_b(.in(layer_1[239]), .out(far_2_2154_0[1]));
    wire [1:0] far_2_2154_1;    relay_conn far_2_2154_1_a(.in(far_2_2154_0[0]), .out(far_2_2154_1[0]));    relay_conn far_2_2154_1_b(.in(far_2_2154_0[1]), .out(far_2_2154_1[1]));
    wire [1:0] far_2_2154_2;    relay_conn far_2_2154_2_a(.in(far_2_2154_1[0]), .out(far_2_2154_2[0]));    relay_conn far_2_2154_2_b(.in(far_2_2154_1[1]), .out(far_2_2154_2[1]));
    assign layer_2[114] = far_2_2154_2[0]; 
    assign layer_2[115] = layer_1[208] & ~layer_1[204]; 
    wire [1:0] far_2_2156_0;    relay_conn far_2_2156_0_a(.in(layer_1[502]), .out(far_2_2156_0[0]));    relay_conn far_2_2156_0_b(.in(layer_1[453]), .out(far_2_2156_0[1]));
    assign layer_2[116] = ~far_2_2156_0[1]; 
    wire [1:0] far_2_2157_0;    relay_conn far_2_2157_0_a(.in(layer_1[409]), .out(far_2_2157_0[0]));    relay_conn far_2_2157_0_b(.in(layer_1[329]), .out(far_2_2157_0[1]));
    wire [1:0] far_2_2157_1;    relay_conn far_2_2157_1_a(.in(far_2_2157_0[0]), .out(far_2_2157_1[0]));    relay_conn far_2_2157_1_b(.in(far_2_2157_0[1]), .out(far_2_2157_1[1]));
    assign layer_2[117] = far_2_2157_1[0] | far_2_2157_1[1]; 
    wire [1:0] far_2_2158_0;    relay_conn far_2_2158_0_a(.in(layer_1[572]), .out(far_2_2158_0[0]));    relay_conn far_2_2158_0_b(.in(layer_1[530]), .out(far_2_2158_0[1]));
    assign layer_2[118] = far_2_2158_0[1] & ~far_2_2158_0[0]; 
    wire [1:0] far_2_2159_0;    relay_conn far_2_2159_0_a(.in(layer_1[312]), .out(far_2_2159_0[0]));    relay_conn far_2_2159_0_b(.in(layer_1[213]), .out(far_2_2159_0[1]));
    wire [1:0] far_2_2159_1;    relay_conn far_2_2159_1_a(.in(far_2_2159_0[0]), .out(far_2_2159_1[0]));    relay_conn far_2_2159_1_b(.in(far_2_2159_0[1]), .out(far_2_2159_1[1]));
    wire [1:0] far_2_2159_2;    relay_conn far_2_2159_2_a(.in(far_2_2159_1[0]), .out(far_2_2159_2[0]));    relay_conn far_2_2159_2_b(.in(far_2_2159_1[1]), .out(far_2_2159_2[1]));
    assign layer_2[119] = far_2_2159_2[0] & far_2_2159_2[1]; 
    wire [1:0] far_2_2160_0;    relay_conn far_2_2160_0_a(.in(layer_1[772]), .out(far_2_2160_0[0]));    relay_conn far_2_2160_0_b(.in(layer_1[652]), .out(far_2_2160_0[1]));
    wire [1:0] far_2_2160_1;    relay_conn far_2_2160_1_a(.in(far_2_2160_0[0]), .out(far_2_2160_1[0]));    relay_conn far_2_2160_1_b(.in(far_2_2160_0[1]), .out(far_2_2160_1[1]));
    wire [1:0] far_2_2160_2;    relay_conn far_2_2160_2_a(.in(far_2_2160_1[0]), .out(far_2_2160_2[0]));    relay_conn far_2_2160_2_b(.in(far_2_2160_1[1]), .out(far_2_2160_2[1]));
    assign layer_2[120] = ~(far_2_2160_2[0] & far_2_2160_2[1]); 
    wire [1:0] far_2_2161_0;    relay_conn far_2_2161_0_a(.in(layer_1[152]), .out(far_2_2161_0[0]));    relay_conn far_2_2161_0_b(.in(layer_1[95]), .out(far_2_2161_0[1]));
    assign layer_2[121] = ~far_2_2161_0[1] | (far_2_2161_0[0] & far_2_2161_0[1]); 
    wire [1:0] far_2_2162_0;    relay_conn far_2_2162_0_a(.in(layer_1[516]), .out(far_2_2162_0[0]));    relay_conn far_2_2162_0_b(.in(layer_1[453]), .out(far_2_2162_0[1]));
    assign layer_2[122] = far_2_2162_0[0] ^ far_2_2162_0[1]; 
    wire [1:0] far_2_2163_0;    relay_conn far_2_2163_0_a(.in(layer_1[682]), .out(far_2_2163_0[0]));    relay_conn far_2_2163_0_b(.in(layer_1[763]), .out(far_2_2163_0[1]));
    wire [1:0] far_2_2163_1;    relay_conn far_2_2163_1_a(.in(far_2_2163_0[0]), .out(far_2_2163_1[0]));    relay_conn far_2_2163_1_b(.in(far_2_2163_0[1]), .out(far_2_2163_1[1]));
    assign layer_2[123] = ~far_2_2163_1[1]; 
    assign layer_2[124] = ~layer_1[160] | (layer_1[160] & layer_1[190]); 
    wire [1:0] far_2_2165_0;    relay_conn far_2_2165_0_a(.in(layer_1[779]), .out(far_2_2165_0[0]));    relay_conn far_2_2165_0_b(.in(layer_1[689]), .out(far_2_2165_0[1]));
    wire [1:0] far_2_2165_1;    relay_conn far_2_2165_1_a(.in(far_2_2165_0[0]), .out(far_2_2165_1[0]));    relay_conn far_2_2165_1_b(.in(far_2_2165_0[1]), .out(far_2_2165_1[1]));
    assign layer_2[125] = far_2_2165_1[0] | far_2_2165_1[1]; 
    assign layer_2[126] = layer_1[888] & ~layer_1[909]; 
    assign layer_2[127] = layer_1[440]; 
    assign layer_2[128] = ~layer_1[954] | (layer_1[954] & layer_1[967]); 
    wire [1:0] far_2_2169_0;    relay_conn far_2_2169_0_a(.in(layer_1[799]), .out(far_2_2169_0[0]));    relay_conn far_2_2169_0_b(.in(layer_1[701]), .out(far_2_2169_0[1]));
    wire [1:0] far_2_2169_1;    relay_conn far_2_2169_1_a(.in(far_2_2169_0[0]), .out(far_2_2169_1[0]));    relay_conn far_2_2169_1_b(.in(far_2_2169_0[1]), .out(far_2_2169_1[1]));
    wire [1:0] far_2_2169_2;    relay_conn far_2_2169_2_a(.in(far_2_2169_1[0]), .out(far_2_2169_2[0]));    relay_conn far_2_2169_2_b(.in(far_2_2169_1[1]), .out(far_2_2169_2[1]));
    assign layer_2[129] = ~far_2_2169_2[1]; 
    wire [1:0] far_2_2170_0;    relay_conn far_2_2170_0_a(.in(layer_1[12]), .out(far_2_2170_0[0]));    relay_conn far_2_2170_0_b(.in(layer_1[55]), .out(far_2_2170_0[1]));
    assign layer_2[130] = far_2_2170_0[0]; 
    wire [1:0] far_2_2171_0;    relay_conn far_2_2171_0_a(.in(layer_1[932]), .out(far_2_2171_0[0]));    relay_conn far_2_2171_0_b(.in(layer_1[1018]), .out(far_2_2171_0[1]));
    wire [1:0] far_2_2171_1;    relay_conn far_2_2171_1_a(.in(far_2_2171_0[0]), .out(far_2_2171_1[0]));    relay_conn far_2_2171_1_b(.in(far_2_2171_0[1]), .out(far_2_2171_1[1]));
    assign layer_2[131] = far_2_2171_1[1]; 
    wire [1:0] far_2_2172_0;    relay_conn far_2_2172_0_a(.in(layer_1[348]), .out(far_2_2172_0[0]));    relay_conn far_2_2172_0_b(.in(layer_1[262]), .out(far_2_2172_0[1]));
    wire [1:0] far_2_2172_1;    relay_conn far_2_2172_1_a(.in(far_2_2172_0[0]), .out(far_2_2172_1[0]));    relay_conn far_2_2172_1_b(.in(far_2_2172_0[1]), .out(far_2_2172_1[1]));
    assign layer_2[132] = far_2_2172_1[1]; 
    wire [1:0] far_2_2173_0;    relay_conn far_2_2173_0_a(.in(layer_1[664]), .out(far_2_2173_0[0]));    relay_conn far_2_2173_0_b(.in(layer_1[724]), .out(far_2_2173_0[1]));
    assign layer_2[133] = far_2_2173_0[0] & far_2_2173_0[1]; 
    assign layer_2[134] = layer_1[419] & layer_1[391]; 
    wire [1:0] far_2_2175_0;    relay_conn far_2_2175_0_a(.in(layer_1[149]), .out(far_2_2175_0[0]));    relay_conn far_2_2175_0_b(.in(layer_1[207]), .out(far_2_2175_0[1]));
    assign layer_2[135] = ~far_2_2175_0[1]; 
    wire [1:0] far_2_2176_0;    relay_conn far_2_2176_0_a(.in(layer_1[596]), .out(far_2_2176_0[0]));    relay_conn far_2_2176_0_b(.in(layer_1[634]), .out(far_2_2176_0[1]));
    assign layer_2[136] = ~(far_2_2176_0[0] & far_2_2176_0[1]); 
    wire [1:0] far_2_2177_0;    relay_conn far_2_2177_0_a(.in(layer_1[543]), .out(far_2_2177_0[0]));    relay_conn far_2_2177_0_b(.in(layer_1[442]), .out(far_2_2177_0[1]));
    wire [1:0] far_2_2177_1;    relay_conn far_2_2177_1_a(.in(far_2_2177_0[0]), .out(far_2_2177_1[0]));    relay_conn far_2_2177_1_b(.in(far_2_2177_0[1]), .out(far_2_2177_1[1]));
    wire [1:0] far_2_2177_2;    relay_conn far_2_2177_2_a(.in(far_2_2177_1[0]), .out(far_2_2177_2[0]));    relay_conn far_2_2177_2_b(.in(far_2_2177_1[1]), .out(far_2_2177_2[1]));
    assign layer_2[137] = ~(far_2_2177_2[0] & far_2_2177_2[1]); 
    wire [1:0] far_2_2178_0;    relay_conn far_2_2178_0_a(.in(layer_1[452]), .out(far_2_2178_0[0]));    relay_conn far_2_2178_0_b(.in(layer_1[334]), .out(far_2_2178_0[1]));
    wire [1:0] far_2_2178_1;    relay_conn far_2_2178_1_a(.in(far_2_2178_0[0]), .out(far_2_2178_1[0]));    relay_conn far_2_2178_1_b(.in(far_2_2178_0[1]), .out(far_2_2178_1[1]));
    wire [1:0] far_2_2178_2;    relay_conn far_2_2178_2_a(.in(far_2_2178_1[0]), .out(far_2_2178_2[0]));    relay_conn far_2_2178_2_b(.in(far_2_2178_1[1]), .out(far_2_2178_2[1]));
    assign layer_2[138] = far_2_2178_2[0] & far_2_2178_2[1]; 
    wire [1:0] far_2_2179_0;    relay_conn far_2_2179_0_a(.in(layer_1[12]), .out(far_2_2179_0[0]));    relay_conn far_2_2179_0_b(.in(layer_1[78]), .out(far_2_2179_0[1]));
    wire [1:0] far_2_2179_1;    relay_conn far_2_2179_1_a(.in(far_2_2179_0[0]), .out(far_2_2179_1[0]));    relay_conn far_2_2179_1_b(.in(far_2_2179_0[1]), .out(far_2_2179_1[1]));
    assign layer_2[139] = ~far_2_2179_1[0] | (far_2_2179_1[0] & far_2_2179_1[1]); 
    wire [1:0] far_2_2180_0;    relay_conn far_2_2180_0_a(.in(layer_1[58]), .out(far_2_2180_0[0]));    relay_conn far_2_2180_0_b(.in(layer_1[159]), .out(far_2_2180_0[1]));
    wire [1:0] far_2_2180_1;    relay_conn far_2_2180_1_a(.in(far_2_2180_0[0]), .out(far_2_2180_1[0]));    relay_conn far_2_2180_1_b(.in(far_2_2180_0[1]), .out(far_2_2180_1[1]));
    wire [1:0] far_2_2180_2;    relay_conn far_2_2180_2_a(.in(far_2_2180_1[0]), .out(far_2_2180_2[0]));    relay_conn far_2_2180_2_b(.in(far_2_2180_1[1]), .out(far_2_2180_2[1]));
    assign layer_2[140] = ~(far_2_2180_2[0] | far_2_2180_2[1]); 
    wire [1:0] far_2_2181_0;    relay_conn far_2_2181_0_a(.in(layer_1[417]), .out(far_2_2181_0[0]));    relay_conn far_2_2181_0_b(.in(layer_1[492]), .out(far_2_2181_0[1]));
    wire [1:0] far_2_2181_1;    relay_conn far_2_2181_1_a(.in(far_2_2181_0[0]), .out(far_2_2181_1[0]));    relay_conn far_2_2181_1_b(.in(far_2_2181_0[1]), .out(far_2_2181_1[1]));
    assign layer_2[141] = ~(far_2_2181_1[0] | far_2_2181_1[1]); 
    assign layer_2[142] = layer_1[885] | layer_1[909]; 
    wire [1:0] far_2_2183_0;    relay_conn far_2_2183_0_a(.in(layer_1[543]), .out(far_2_2183_0[0]));    relay_conn far_2_2183_0_b(.in(layer_1[577]), .out(far_2_2183_0[1]));
    assign layer_2[143] = far_2_2183_0[0] & ~far_2_2183_0[1]; 
    assign layer_2[144] = layer_1[248]; 
    wire [1:0] far_2_2185_0;    relay_conn far_2_2185_0_a(.in(layer_1[533]), .out(far_2_2185_0[0]));    relay_conn far_2_2185_0_b(.in(layer_1[417]), .out(far_2_2185_0[1]));
    wire [1:0] far_2_2185_1;    relay_conn far_2_2185_1_a(.in(far_2_2185_0[0]), .out(far_2_2185_1[0]));    relay_conn far_2_2185_1_b(.in(far_2_2185_0[1]), .out(far_2_2185_1[1]));
    wire [1:0] far_2_2185_2;    relay_conn far_2_2185_2_a(.in(far_2_2185_1[0]), .out(far_2_2185_2[0]));    relay_conn far_2_2185_2_b(.in(far_2_2185_1[1]), .out(far_2_2185_2[1]));
    assign layer_2[145] = ~(far_2_2185_2[0] & far_2_2185_2[1]); 
    wire [1:0] far_2_2186_0;    relay_conn far_2_2186_0_a(.in(layer_1[183]), .out(far_2_2186_0[0]));    relay_conn far_2_2186_0_b(.in(layer_1[62]), .out(far_2_2186_0[1]));
    wire [1:0] far_2_2186_1;    relay_conn far_2_2186_1_a(.in(far_2_2186_0[0]), .out(far_2_2186_1[0]));    relay_conn far_2_2186_1_b(.in(far_2_2186_0[1]), .out(far_2_2186_1[1]));
    wire [1:0] far_2_2186_2;    relay_conn far_2_2186_2_a(.in(far_2_2186_1[0]), .out(far_2_2186_2[0]));    relay_conn far_2_2186_2_b(.in(far_2_2186_1[1]), .out(far_2_2186_2[1]));
    assign layer_2[146] = far_2_2186_2[0] | far_2_2186_2[1]; 
    assign layer_2[147] = layer_1[898] | layer_1[910]; 
    wire [1:0] far_2_2188_0;    relay_conn far_2_2188_0_a(.in(layer_1[249]), .out(far_2_2188_0[0]));    relay_conn far_2_2188_0_b(.in(layer_1[177]), .out(far_2_2188_0[1]));
    wire [1:0] far_2_2188_1;    relay_conn far_2_2188_1_a(.in(far_2_2188_0[0]), .out(far_2_2188_1[0]));    relay_conn far_2_2188_1_b(.in(far_2_2188_0[1]), .out(far_2_2188_1[1]));
    assign layer_2[148] = ~(far_2_2188_1[0] | far_2_2188_1[1]); 
    assign layer_2[149] = layer_1[248] ^ layer_1[230]; 
    assign layer_2[150] = ~layer_1[309]; 
    wire [1:0] far_2_2191_0;    relay_conn far_2_2191_0_a(.in(layer_1[323]), .out(far_2_2191_0[0]));    relay_conn far_2_2191_0_b(.in(layer_1[416]), .out(far_2_2191_0[1]));
    wire [1:0] far_2_2191_1;    relay_conn far_2_2191_1_a(.in(far_2_2191_0[0]), .out(far_2_2191_1[0]));    relay_conn far_2_2191_1_b(.in(far_2_2191_0[1]), .out(far_2_2191_1[1]));
    assign layer_2[151] = far_2_2191_1[0] & ~far_2_2191_1[1]; 
    assign layer_2[152] = layer_1[368] | layer_1[364]; 
    wire [1:0] far_2_2193_0;    relay_conn far_2_2193_0_a(.in(layer_1[619]), .out(far_2_2193_0[0]));    relay_conn far_2_2193_0_b(.in(layer_1[546]), .out(far_2_2193_0[1]));
    wire [1:0] far_2_2193_1;    relay_conn far_2_2193_1_a(.in(far_2_2193_0[0]), .out(far_2_2193_1[0]));    relay_conn far_2_2193_1_b(.in(far_2_2193_0[1]), .out(far_2_2193_1[1]));
    assign layer_2[153] = ~far_2_2193_1[1]; 
    wire [1:0] far_2_2194_0;    relay_conn far_2_2194_0_a(.in(layer_1[270]), .out(far_2_2194_0[0]));    relay_conn far_2_2194_0_b(.in(layer_1[218]), .out(far_2_2194_0[1]));
    assign layer_2[154] = far_2_2194_0[0] & ~far_2_2194_0[1]; 
    wire [1:0] far_2_2195_0;    relay_conn far_2_2195_0_a(.in(layer_1[772]), .out(far_2_2195_0[0]));    relay_conn far_2_2195_0_b(.in(layer_1[685]), .out(far_2_2195_0[1]));
    wire [1:0] far_2_2195_1;    relay_conn far_2_2195_1_a(.in(far_2_2195_0[0]), .out(far_2_2195_1[0]));    relay_conn far_2_2195_1_b(.in(far_2_2195_0[1]), .out(far_2_2195_1[1]));
    assign layer_2[155] = ~(far_2_2195_1[0] & far_2_2195_1[1]); 
    wire [1:0] far_2_2196_0;    relay_conn far_2_2196_0_a(.in(layer_1[784]), .out(far_2_2196_0[0]));    relay_conn far_2_2196_0_b(.in(layer_1[715]), .out(far_2_2196_0[1]));
    wire [1:0] far_2_2196_1;    relay_conn far_2_2196_1_a(.in(far_2_2196_0[0]), .out(far_2_2196_1[0]));    relay_conn far_2_2196_1_b(.in(far_2_2196_0[1]), .out(far_2_2196_1[1]));
    assign layer_2[156] = ~(far_2_2196_1[0] & far_2_2196_1[1]); 
    wire [1:0] far_2_2197_0;    relay_conn far_2_2197_0_a(.in(layer_1[918]), .out(far_2_2197_0[0]));    relay_conn far_2_2197_0_b(.in(layer_1[995]), .out(far_2_2197_0[1]));
    wire [1:0] far_2_2197_1;    relay_conn far_2_2197_1_a(.in(far_2_2197_0[0]), .out(far_2_2197_1[0]));    relay_conn far_2_2197_1_b(.in(far_2_2197_0[1]), .out(far_2_2197_1[1]));
    assign layer_2[157] = ~(far_2_2197_1[0] | far_2_2197_1[1]); 
    wire [1:0] far_2_2198_0;    relay_conn far_2_2198_0_a(.in(layer_1[643]), .out(far_2_2198_0[0]));    relay_conn far_2_2198_0_b(.in(layer_1[520]), .out(far_2_2198_0[1]));
    wire [1:0] far_2_2198_1;    relay_conn far_2_2198_1_a(.in(far_2_2198_0[0]), .out(far_2_2198_1[0]));    relay_conn far_2_2198_1_b(.in(far_2_2198_0[1]), .out(far_2_2198_1[1]));
    wire [1:0] far_2_2198_2;    relay_conn far_2_2198_2_a(.in(far_2_2198_1[0]), .out(far_2_2198_2[0]));    relay_conn far_2_2198_2_b(.in(far_2_2198_1[1]), .out(far_2_2198_2[1]));
    assign layer_2[158] = far_2_2198_2[0] & far_2_2198_2[1]; 
    wire [1:0] far_2_2199_0;    relay_conn far_2_2199_0_a(.in(layer_1[932]), .out(far_2_2199_0[0]));    relay_conn far_2_2199_0_b(.in(layer_1[820]), .out(far_2_2199_0[1]));
    wire [1:0] far_2_2199_1;    relay_conn far_2_2199_1_a(.in(far_2_2199_0[0]), .out(far_2_2199_1[0]));    relay_conn far_2_2199_1_b(.in(far_2_2199_0[1]), .out(far_2_2199_1[1]));
    wire [1:0] far_2_2199_2;    relay_conn far_2_2199_2_a(.in(far_2_2199_1[0]), .out(far_2_2199_2[0]));    relay_conn far_2_2199_2_b(.in(far_2_2199_1[1]), .out(far_2_2199_2[1]));
    assign layer_2[159] = far_2_2199_2[0] & far_2_2199_2[1]; 
    wire [1:0] far_2_2200_0;    relay_conn far_2_2200_0_a(.in(layer_1[855]), .out(far_2_2200_0[0]));    relay_conn far_2_2200_0_b(.in(layer_1[888]), .out(far_2_2200_0[1]));
    assign layer_2[160] = far_2_2200_0[1]; 
    wire [1:0] far_2_2201_0;    relay_conn far_2_2201_0_a(.in(layer_1[962]), .out(far_2_2201_0[0]));    relay_conn far_2_2201_0_b(.in(layer_1[1018]), .out(far_2_2201_0[1]));
    assign layer_2[161] = ~(far_2_2201_0[0] & far_2_2201_0[1]); 
    wire [1:0] far_2_2202_0;    relay_conn far_2_2202_0_a(.in(layer_1[829]), .out(far_2_2202_0[0]));    relay_conn far_2_2202_0_b(.in(layer_1[898]), .out(far_2_2202_0[1]));
    wire [1:0] far_2_2202_1;    relay_conn far_2_2202_1_a(.in(far_2_2202_0[0]), .out(far_2_2202_1[0]));    relay_conn far_2_2202_1_b(.in(far_2_2202_0[1]), .out(far_2_2202_1[1]));
    assign layer_2[162] = far_2_2202_1[1] & ~far_2_2202_1[0]; 
    assign layer_2[163] = ~layer_1[328] | (layer_1[321] & layer_1[328]); 
    wire [1:0] far_2_2204_0;    relay_conn far_2_2204_0_a(.in(layer_1[569]), .out(far_2_2204_0[0]));    relay_conn far_2_2204_0_b(.in(layer_1[533]), .out(far_2_2204_0[1]));
    assign layer_2[164] = far_2_2204_0[1] & ~far_2_2204_0[0]; 
    wire [1:0] far_2_2205_0;    relay_conn far_2_2205_0_a(.in(layer_1[622]), .out(far_2_2205_0[0]));    relay_conn far_2_2205_0_b(.in(layer_1[687]), .out(far_2_2205_0[1]));
    wire [1:0] far_2_2205_1;    relay_conn far_2_2205_1_a(.in(far_2_2205_0[0]), .out(far_2_2205_1[0]));    relay_conn far_2_2205_1_b(.in(far_2_2205_0[1]), .out(far_2_2205_1[1]));
    assign layer_2[165] = far_2_2205_1[0] & far_2_2205_1[1]; 
    wire [1:0] far_2_2206_0;    relay_conn far_2_2206_0_a(.in(layer_1[444]), .out(far_2_2206_0[0]));    relay_conn far_2_2206_0_b(.in(layer_1[364]), .out(far_2_2206_0[1]));
    wire [1:0] far_2_2206_1;    relay_conn far_2_2206_1_a(.in(far_2_2206_0[0]), .out(far_2_2206_1[0]));    relay_conn far_2_2206_1_b(.in(far_2_2206_0[1]), .out(far_2_2206_1[1]));
    assign layer_2[166] = ~(far_2_2206_1[0] | far_2_2206_1[1]); 
    assign layer_2[167] = layer_1[623]; 
    wire [1:0] far_2_2208_0;    relay_conn far_2_2208_0_a(.in(layer_1[795]), .out(far_2_2208_0[0]));    relay_conn far_2_2208_0_b(.in(layer_1[837]), .out(far_2_2208_0[1]));
    assign layer_2[168] = ~far_2_2208_0[0] | (far_2_2208_0[0] & far_2_2208_0[1]); 
    wire [1:0] far_2_2209_0;    relay_conn far_2_2209_0_a(.in(layer_1[891]), .out(far_2_2209_0[0]));    relay_conn far_2_2209_0_b(.in(layer_1[776]), .out(far_2_2209_0[1]));
    wire [1:0] far_2_2209_1;    relay_conn far_2_2209_1_a(.in(far_2_2209_0[0]), .out(far_2_2209_1[0]));    relay_conn far_2_2209_1_b(.in(far_2_2209_0[1]), .out(far_2_2209_1[1]));
    wire [1:0] far_2_2209_2;    relay_conn far_2_2209_2_a(.in(far_2_2209_1[0]), .out(far_2_2209_2[0]));    relay_conn far_2_2209_2_b(.in(far_2_2209_1[1]), .out(far_2_2209_2[1]));
    assign layer_2[169] = far_2_2209_2[0] & ~far_2_2209_2[1]; 
    wire [1:0] far_2_2210_0;    relay_conn far_2_2210_0_a(.in(layer_1[837]), .out(far_2_2210_0[0]));    relay_conn far_2_2210_0_b(.in(layer_1[955]), .out(far_2_2210_0[1]));
    wire [1:0] far_2_2210_1;    relay_conn far_2_2210_1_a(.in(far_2_2210_0[0]), .out(far_2_2210_1[0]));    relay_conn far_2_2210_1_b(.in(far_2_2210_0[1]), .out(far_2_2210_1[1]));
    wire [1:0] far_2_2210_2;    relay_conn far_2_2210_2_a(.in(far_2_2210_1[0]), .out(far_2_2210_2[0]));    relay_conn far_2_2210_2_b(.in(far_2_2210_1[1]), .out(far_2_2210_2[1]));
    assign layer_2[170] = far_2_2210_2[1] & ~far_2_2210_2[0]; 
    wire [1:0] far_2_2211_0;    relay_conn far_2_2211_0_a(.in(layer_1[692]), .out(far_2_2211_0[0]));    relay_conn far_2_2211_0_b(.in(layer_1[575]), .out(far_2_2211_0[1]));
    wire [1:0] far_2_2211_1;    relay_conn far_2_2211_1_a(.in(far_2_2211_0[0]), .out(far_2_2211_1[0]));    relay_conn far_2_2211_1_b(.in(far_2_2211_0[1]), .out(far_2_2211_1[1]));
    wire [1:0] far_2_2211_2;    relay_conn far_2_2211_2_a(.in(far_2_2211_1[0]), .out(far_2_2211_2[0]));    relay_conn far_2_2211_2_b(.in(far_2_2211_1[1]), .out(far_2_2211_2[1]));
    assign layer_2[171] = ~far_2_2211_2[0]; 
    wire [1:0] far_2_2212_0;    relay_conn far_2_2212_0_a(.in(layer_1[507]), .out(far_2_2212_0[0]));    relay_conn far_2_2212_0_b(.in(layer_1[457]), .out(far_2_2212_0[1]));
    assign layer_2[172] = far_2_2212_0[0] & ~far_2_2212_0[1]; 
    wire [1:0] far_2_2213_0;    relay_conn far_2_2213_0_a(.in(layer_1[875]), .out(far_2_2213_0[0]));    relay_conn far_2_2213_0_b(.in(layer_1[768]), .out(far_2_2213_0[1]));
    wire [1:0] far_2_2213_1;    relay_conn far_2_2213_1_a(.in(far_2_2213_0[0]), .out(far_2_2213_1[0]));    relay_conn far_2_2213_1_b(.in(far_2_2213_0[1]), .out(far_2_2213_1[1]));
    wire [1:0] far_2_2213_2;    relay_conn far_2_2213_2_a(.in(far_2_2213_1[0]), .out(far_2_2213_2[0]));    relay_conn far_2_2213_2_b(.in(far_2_2213_1[1]), .out(far_2_2213_2[1]));
    assign layer_2[173] = ~(far_2_2213_2[0] | far_2_2213_2[1]); 
    wire [1:0] far_2_2214_0;    relay_conn far_2_2214_0_a(.in(layer_1[12]), .out(far_2_2214_0[0]));    relay_conn far_2_2214_0_b(.in(layer_1[82]), .out(far_2_2214_0[1]));
    wire [1:0] far_2_2214_1;    relay_conn far_2_2214_1_a(.in(far_2_2214_0[0]), .out(far_2_2214_1[0]));    relay_conn far_2_2214_1_b(.in(far_2_2214_0[1]), .out(far_2_2214_1[1]));
    assign layer_2[174] = ~(far_2_2214_1[0] & far_2_2214_1[1]); 
    assign layer_2[175] = layer_1[50] & ~layer_1[53]; 
    wire [1:0] far_2_2216_0;    relay_conn far_2_2216_0_a(.in(layer_1[239]), .out(far_2_2216_0[0]));    relay_conn far_2_2216_0_b(.in(layer_1[349]), .out(far_2_2216_0[1]));
    wire [1:0] far_2_2216_1;    relay_conn far_2_2216_1_a(.in(far_2_2216_0[0]), .out(far_2_2216_1[0]));    relay_conn far_2_2216_1_b(.in(far_2_2216_0[1]), .out(far_2_2216_1[1]));
    wire [1:0] far_2_2216_2;    relay_conn far_2_2216_2_a(.in(far_2_2216_1[0]), .out(far_2_2216_2[0]));    relay_conn far_2_2216_2_b(.in(far_2_2216_1[1]), .out(far_2_2216_2[1]));
    assign layer_2[176] = far_2_2216_2[1]; 
    wire [1:0] far_2_2217_0;    relay_conn far_2_2217_0_a(.in(layer_1[796]), .out(far_2_2217_0[0]));    relay_conn far_2_2217_0_b(.in(layer_1[867]), .out(far_2_2217_0[1]));
    wire [1:0] far_2_2217_1;    relay_conn far_2_2217_1_a(.in(far_2_2217_0[0]), .out(far_2_2217_1[0]));    relay_conn far_2_2217_1_b(.in(far_2_2217_0[1]), .out(far_2_2217_1[1]));
    assign layer_2[177] = ~far_2_2217_1[1]; 
    wire [1:0] far_2_2218_0;    relay_conn far_2_2218_0_a(.in(layer_1[569]), .out(far_2_2218_0[0]));    relay_conn far_2_2218_0_b(.in(layer_1[688]), .out(far_2_2218_0[1]));
    wire [1:0] far_2_2218_1;    relay_conn far_2_2218_1_a(.in(far_2_2218_0[0]), .out(far_2_2218_1[0]));    relay_conn far_2_2218_1_b(.in(far_2_2218_0[1]), .out(far_2_2218_1[1]));
    wire [1:0] far_2_2218_2;    relay_conn far_2_2218_2_a(.in(far_2_2218_1[0]), .out(far_2_2218_2[0]));    relay_conn far_2_2218_2_b(.in(far_2_2218_1[1]), .out(far_2_2218_2[1]));
    assign layer_2[178] = ~far_2_2218_2[0]; 
    wire [1:0] far_2_2219_0;    relay_conn far_2_2219_0_a(.in(layer_1[18]), .out(far_2_2219_0[0]));    relay_conn far_2_2219_0_b(.in(layer_1[118]), .out(far_2_2219_0[1]));
    wire [1:0] far_2_2219_1;    relay_conn far_2_2219_1_a(.in(far_2_2219_0[0]), .out(far_2_2219_1[0]));    relay_conn far_2_2219_1_b(.in(far_2_2219_0[1]), .out(far_2_2219_1[1]));
    wire [1:0] far_2_2219_2;    relay_conn far_2_2219_2_a(.in(far_2_2219_1[0]), .out(far_2_2219_2[0]));    relay_conn far_2_2219_2_b(.in(far_2_2219_1[1]), .out(far_2_2219_2[1]));
    assign layer_2[179] = ~far_2_2219_2[1] | (far_2_2219_2[0] & far_2_2219_2[1]); 
    wire [1:0] far_2_2220_0;    relay_conn far_2_2220_0_a(.in(layer_1[987]), .out(far_2_2220_0[0]));    relay_conn far_2_2220_0_b(.in(layer_1[955]), .out(far_2_2220_0[1]));
    assign layer_2[180] = ~far_2_2220_0[1] | (far_2_2220_0[0] & far_2_2220_0[1]); 
    wire [1:0] far_2_2221_0;    relay_conn far_2_2221_0_a(.in(layer_1[732]), .out(far_2_2221_0[0]));    relay_conn far_2_2221_0_b(.in(layer_1[653]), .out(far_2_2221_0[1]));
    wire [1:0] far_2_2221_1;    relay_conn far_2_2221_1_a(.in(far_2_2221_0[0]), .out(far_2_2221_1[0]));    relay_conn far_2_2221_1_b(.in(far_2_2221_0[1]), .out(far_2_2221_1[1]));
    assign layer_2[181] = ~(far_2_2221_1[0] | far_2_2221_1[1]); 
    assign layer_2[182] = ~(layer_1[319] & layer_1[315]); 
    wire [1:0] far_2_2223_0;    relay_conn far_2_2223_0_a(.in(layer_1[50]), .out(far_2_2223_0[0]));    relay_conn far_2_2223_0_b(.in(layer_1[82]), .out(far_2_2223_0[1]));
    assign layer_2[183] = far_2_2223_0[0] | far_2_2223_0[1]; 
    wire [1:0] far_2_2224_0;    relay_conn far_2_2224_0_a(.in(layer_1[1007]), .out(far_2_2224_0[0]));    relay_conn far_2_2224_0_b(.in(layer_1[918]), .out(far_2_2224_0[1]));
    wire [1:0] far_2_2224_1;    relay_conn far_2_2224_1_a(.in(far_2_2224_0[0]), .out(far_2_2224_1[0]));    relay_conn far_2_2224_1_b(.in(far_2_2224_0[1]), .out(far_2_2224_1[1]));
    assign layer_2[184] = ~far_2_2224_1[1]; 
    wire [1:0] far_2_2225_0;    relay_conn far_2_2225_0_a(.in(layer_1[918]), .out(far_2_2225_0[0]));    relay_conn far_2_2225_0_b(.in(layer_1[997]), .out(far_2_2225_0[1]));
    wire [1:0] far_2_2225_1;    relay_conn far_2_2225_1_a(.in(far_2_2225_0[0]), .out(far_2_2225_1[0]));    relay_conn far_2_2225_1_b(.in(far_2_2225_0[1]), .out(far_2_2225_1[1]));
    assign layer_2[185] = far_2_2225_1[1] & ~far_2_2225_1[0]; 
    wire [1:0] far_2_2226_0;    relay_conn far_2_2226_0_a(.in(layer_1[759]), .out(far_2_2226_0[0]));    relay_conn far_2_2226_0_b(.in(layer_1[867]), .out(far_2_2226_0[1]));
    wire [1:0] far_2_2226_1;    relay_conn far_2_2226_1_a(.in(far_2_2226_0[0]), .out(far_2_2226_1[0]));    relay_conn far_2_2226_1_b(.in(far_2_2226_0[1]), .out(far_2_2226_1[1]));
    wire [1:0] far_2_2226_2;    relay_conn far_2_2226_2_a(.in(far_2_2226_1[0]), .out(far_2_2226_2[0]));    relay_conn far_2_2226_2_b(.in(far_2_2226_1[1]), .out(far_2_2226_2[1]));
    assign layer_2[186] = far_2_2226_2[0] ^ far_2_2226_2[1]; 
    wire [1:0] far_2_2227_0;    relay_conn far_2_2227_0_a(.in(layer_1[471]), .out(far_2_2227_0[0]));    relay_conn far_2_2227_0_b(.in(layer_1[537]), .out(far_2_2227_0[1]));
    wire [1:0] far_2_2227_1;    relay_conn far_2_2227_1_a(.in(far_2_2227_0[0]), .out(far_2_2227_1[0]));    relay_conn far_2_2227_1_b(.in(far_2_2227_0[1]), .out(far_2_2227_1[1]));
    assign layer_2[187] = ~far_2_2227_1[0] | (far_2_2227_1[0] & far_2_2227_1[1]); 
    wire [1:0] far_2_2228_0;    relay_conn far_2_2228_0_a(.in(layer_1[169]), .out(far_2_2228_0[0]));    relay_conn far_2_2228_0_b(.in(layer_1[119]), .out(far_2_2228_0[1]));
    assign layer_2[188] = ~far_2_2228_0[0]; 
    wire [1:0] far_2_2229_0;    relay_conn far_2_2229_0_a(.in(layer_1[188]), .out(far_2_2229_0[0]));    relay_conn far_2_2229_0_b(.in(layer_1[88]), .out(far_2_2229_0[1]));
    wire [1:0] far_2_2229_1;    relay_conn far_2_2229_1_a(.in(far_2_2229_0[0]), .out(far_2_2229_1[0]));    relay_conn far_2_2229_1_b(.in(far_2_2229_0[1]), .out(far_2_2229_1[1]));
    wire [1:0] far_2_2229_2;    relay_conn far_2_2229_2_a(.in(far_2_2229_1[0]), .out(far_2_2229_2[0]));    relay_conn far_2_2229_2_b(.in(far_2_2229_1[1]), .out(far_2_2229_2[1]));
    assign layer_2[189] = ~far_2_2229_2[0]; 
    wire [1:0] far_2_2230_0;    relay_conn far_2_2230_0_a(.in(layer_1[345]), .out(far_2_2230_0[0]));    relay_conn far_2_2230_0_b(.in(layer_1[469]), .out(far_2_2230_0[1]));
    wire [1:0] far_2_2230_1;    relay_conn far_2_2230_1_a(.in(far_2_2230_0[0]), .out(far_2_2230_1[0]));    relay_conn far_2_2230_1_b(.in(far_2_2230_0[1]), .out(far_2_2230_1[1]));
    wire [1:0] far_2_2230_2;    relay_conn far_2_2230_2_a(.in(far_2_2230_1[0]), .out(far_2_2230_2[0]));    relay_conn far_2_2230_2_b(.in(far_2_2230_1[1]), .out(far_2_2230_2[1]));
    assign layer_2[190] = far_2_2230_2[0] ^ far_2_2230_2[1]; 
    wire [1:0] far_2_2231_0;    relay_conn far_2_2231_0_a(.in(layer_1[972]), .out(far_2_2231_0[0]));    relay_conn far_2_2231_0_b(.in(layer_1[881]), .out(far_2_2231_0[1]));
    wire [1:0] far_2_2231_1;    relay_conn far_2_2231_1_a(.in(far_2_2231_0[0]), .out(far_2_2231_1[0]));    relay_conn far_2_2231_1_b(.in(far_2_2231_0[1]), .out(far_2_2231_1[1]));
    assign layer_2[191] = far_2_2231_1[1] & ~far_2_2231_1[0]; 
    wire [1:0] far_2_2232_0;    relay_conn far_2_2232_0_a(.in(layer_1[155]), .out(far_2_2232_0[0]));    relay_conn far_2_2232_0_b(.in(layer_1[63]), .out(far_2_2232_0[1]));
    wire [1:0] far_2_2232_1;    relay_conn far_2_2232_1_a(.in(far_2_2232_0[0]), .out(far_2_2232_1[0]));    relay_conn far_2_2232_1_b(.in(far_2_2232_0[1]), .out(far_2_2232_1[1]));
    assign layer_2[192] = far_2_2232_1[0] & far_2_2232_1[1]; 
    wire [1:0] far_2_2233_0;    relay_conn far_2_2233_0_a(.in(layer_1[352]), .out(far_2_2233_0[0]));    relay_conn far_2_2233_0_b(.in(layer_1[272]), .out(far_2_2233_0[1]));
    wire [1:0] far_2_2233_1;    relay_conn far_2_2233_1_a(.in(far_2_2233_0[0]), .out(far_2_2233_1[0]));    relay_conn far_2_2233_1_b(.in(far_2_2233_0[1]), .out(far_2_2233_1[1]));
    assign layer_2[193] = ~(far_2_2233_1[0] | far_2_2233_1[1]); 
    assign layer_2[194] = ~(layer_1[446] | layer_1[430]); 
    wire [1:0] far_2_2235_0;    relay_conn far_2_2235_0_a(.in(layer_1[102]), .out(far_2_2235_0[0]));    relay_conn far_2_2235_0_b(.in(layer_1[39]), .out(far_2_2235_0[1]));
    assign layer_2[195] = ~far_2_2235_0[1] | (far_2_2235_0[0] & far_2_2235_0[1]); 
    wire [1:0] far_2_2236_0;    relay_conn far_2_2236_0_a(.in(layer_1[329]), .out(far_2_2236_0[0]));    relay_conn far_2_2236_0_b(.in(layer_1[238]), .out(far_2_2236_0[1]));
    wire [1:0] far_2_2236_1;    relay_conn far_2_2236_1_a(.in(far_2_2236_0[0]), .out(far_2_2236_1[0]));    relay_conn far_2_2236_1_b(.in(far_2_2236_0[1]), .out(far_2_2236_1[1]));
    assign layer_2[196] = far_2_2236_1[0] & far_2_2236_1[1]; 
    wire [1:0] far_2_2237_0;    relay_conn far_2_2237_0_a(.in(layer_1[41]), .out(far_2_2237_0[0]));    relay_conn far_2_2237_0_b(.in(layer_1[133]), .out(far_2_2237_0[1]));
    wire [1:0] far_2_2237_1;    relay_conn far_2_2237_1_a(.in(far_2_2237_0[0]), .out(far_2_2237_1[0]));    relay_conn far_2_2237_1_b(.in(far_2_2237_0[1]), .out(far_2_2237_1[1]));
    assign layer_2[197] = far_2_2237_1[0] | far_2_2237_1[1]; 
    wire [1:0] far_2_2238_0;    relay_conn far_2_2238_0_a(.in(layer_1[498]), .out(far_2_2238_0[0]));    relay_conn far_2_2238_0_b(.in(layer_1[419]), .out(far_2_2238_0[1]));
    wire [1:0] far_2_2238_1;    relay_conn far_2_2238_1_a(.in(far_2_2238_0[0]), .out(far_2_2238_1[0]));    relay_conn far_2_2238_1_b(.in(far_2_2238_0[1]), .out(far_2_2238_1[1]));
    assign layer_2[198] = far_2_2238_1[0] & far_2_2238_1[1]; 
    wire [1:0] far_2_2239_0;    relay_conn far_2_2239_0_a(.in(layer_1[642]), .out(far_2_2239_0[0]));    relay_conn far_2_2239_0_b(.in(layer_1[555]), .out(far_2_2239_0[1]));
    wire [1:0] far_2_2239_1;    relay_conn far_2_2239_1_a(.in(far_2_2239_0[0]), .out(far_2_2239_1[0]));    relay_conn far_2_2239_1_b(.in(far_2_2239_0[1]), .out(far_2_2239_1[1]));
    assign layer_2[199] = ~far_2_2239_1[1]; 
    wire [1:0] far_2_2240_0;    relay_conn far_2_2240_0_a(.in(layer_1[733]), .out(far_2_2240_0[0]));    relay_conn far_2_2240_0_b(.in(layer_1[846]), .out(far_2_2240_0[1]));
    wire [1:0] far_2_2240_1;    relay_conn far_2_2240_1_a(.in(far_2_2240_0[0]), .out(far_2_2240_1[0]));    relay_conn far_2_2240_1_b(.in(far_2_2240_0[1]), .out(far_2_2240_1[1]));
    wire [1:0] far_2_2240_2;    relay_conn far_2_2240_2_a(.in(far_2_2240_1[0]), .out(far_2_2240_2[0]));    relay_conn far_2_2240_2_b(.in(far_2_2240_1[1]), .out(far_2_2240_2[1]));
    assign layer_2[200] = ~far_2_2240_2[0] | (far_2_2240_2[0] & far_2_2240_2[1]); 
    wire [1:0] far_2_2241_0;    relay_conn far_2_2241_0_a(.in(layer_1[946]), .out(far_2_2241_0[0]));    relay_conn far_2_2241_0_b(.in(layer_1[836]), .out(far_2_2241_0[1]));
    wire [1:0] far_2_2241_1;    relay_conn far_2_2241_1_a(.in(far_2_2241_0[0]), .out(far_2_2241_1[0]));    relay_conn far_2_2241_1_b(.in(far_2_2241_0[1]), .out(far_2_2241_1[1]));
    wire [1:0] far_2_2241_2;    relay_conn far_2_2241_2_a(.in(far_2_2241_1[0]), .out(far_2_2241_2[0]));    relay_conn far_2_2241_2_b(.in(far_2_2241_1[1]), .out(far_2_2241_2[1]));
    assign layer_2[201] = ~far_2_2241_2[0]; 
    wire [1:0] far_2_2242_0;    relay_conn far_2_2242_0_a(.in(layer_1[206]), .out(far_2_2242_0[0]));    relay_conn far_2_2242_0_b(.in(layer_1[319]), .out(far_2_2242_0[1]));
    wire [1:0] far_2_2242_1;    relay_conn far_2_2242_1_a(.in(far_2_2242_0[0]), .out(far_2_2242_1[0]));    relay_conn far_2_2242_1_b(.in(far_2_2242_0[1]), .out(far_2_2242_1[1]));
    wire [1:0] far_2_2242_2;    relay_conn far_2_2242_2_a(.in(far_2_2242_1[0]), .out(far_2_2242_2[0]));    relay_conn far_2_2242_2_b(.in(far_2_2242_1[1]), .out(far_2_2242_2[1]));
    assign layer_2[202] = ~far_2_2242_2[1] | (far_2_2242_2[0] & far_2_2242_2[1]); 
    wire [1:0] far_2_2243_0;    relay_conn far_2_2243_0_a(.in(layer_1[688]), .out(far_2_2243_0[0]));    relay_conn far_2_2243_0_b(.in(layer_1[573]), .out(far_2_2243_0[1]));
    wire [1:0] far_2_2243_1;    relay_conn far_2_2243_1_a(.in(far_2_2243_0[0]), .out(far_2_2243_1[0]));    relay_conn far_2_2243_1_b(.in(far_2_2243_0[1]), .out(far_2_2243_1[1]));
    wire [1:0] far_2_2243_2;    relay_conn far_2_2243_2_a(.in(far_2_2243_1[0]), .out(far_2_2243_2[0]));    relay_conn far_2_2243_2_b(.in(far_2_2243_1[1]), .out(far_2_2243_2[1]));
    assign layer_2[203] = ~(far_2_2243_2[0] | far_2_2243_2[1]); 
    wire [1:0] far_2_2244_0;    relay_conn far_2_2244_0_a(.in(layer_1[733]), .out(far_2_2244_0[0]));    relay_conn far_2_2244_0_b(.in(layer_1[772]), .out(far_2_2244_0[1]));
    assign layer_2[204] = far_2_2244_0[1]; 
    wire [1:0] far_2_2245_0;    relay_conn far_2_2245_0_a(.in(layer_1[895]), .out(far_2_2245_0[0]));    relay_conn far_2_2245_0_b(.in(layer_1[844]), .out(far_2_2245_0[1]));
    assign layer_2[205] = ~far_2_2245_0[1] | (far_2_2245_0[0] & far_2_2245_0[1]); 
    wire [1:0] far_2_2246_0;    relay_conn far_2_2246_0_a(.in(layer_1[707]), .out(far_2_2246_0[0]));    relay_conn far_2_2246_0_b(.in(layer_1[749]), .out(far_2_2246_0[1]));
    assign layer_2[206] = far_2_2246_0[1]; 
    assign layer_2[207] = ~(layer_1[37] | layer_1[67]); 
    assign layer_2[208] = layer_1[333] | layer_1[312]; 
    wire [1:0] far_2_2249_0;    relay_conn far_2_2249_0_a(.in(layer_1[193]), .out(far_2_2249_0[0]));    relay_conn far_2_2249_0_b(.in(layer_1[139]), .out(far_2_2249_0[1]));
    assign layer_2[209] = far_2_2249_0[0]; 
    wire [1:0] far_2_2250_0;    relay_conn far_2_2250_0_a(.in(layer_1[795]), .out(far_2_2250_0[0]));    relay_conn far_2_2250_0_b(.in(layer_1[701]), .out(far_2_2250_0[1]));
    wire [1:0] far_2_2250_1;    relay_conn far_2_2250_1_a(.in(far_2_2250_0[0]), .out(far_2_2250_1[0]));    relay_conn far_2_2250_1_b(.in(far_2_2250_0[1]), .out(far_2_2250_1[1]));
    assign layer_2[210] = ~(far_2_2250_1[0] ^ far_2_2250_1[1]); 
    wire [1:0] far_2_2251_0;    relay_conn far_2_2251_0_a(.in(layer_1[84]), .out(far_2_2251_0[0]));    relay_conn far_2_2251_0_b(.in(layer_1[121]), .out(far_2_2251_0[1]));
    assign layer_2[211] = ~far_2_2251_0[0]; 
    wire [1:0] far_2_2252_0;    relay_conn far_2_2252_0_a(.in(layer_1[561]), .out(far_2_2252_0[0]));    relay_conn far_2_2252_0_b(.in(layer_1[459]), .out(far_2_2252_0[1]));
    wire [1:0] far_2_2252_1;    relay_conn far_2_2252_1_a(.in(far_2_2252_0[0]), .out(far_2_2252_1[0]));    relay_conn far_2_2252_1_b(.in(far_2_2252_0[1]), .out(far_2_2252_1[1]));
    wire [1:0] far_2_2252_2;    relay_conn far_2_2252_2_a(.in(far_2_2252_1[0]), .out(far_2_2252_2[0]));    relay_conn far_2_2252_2_b(.in(far_2_2252_1[1]), .out(far_2_2252_2[1]));
    assign layer_2[212] = ~far_2_2252_2[1] | (far_2_2252_2[0] & far_2_2252_2[1]); 
    wire [1:0] far_2_2253_0;    relay_conn far_2_2253_0_a(.in(layer_1[784]), .out(far_2_2253_0[0]));    relay_conn far_2_2253_0_b(.in(layer_1[720]), .out(far_2_2253_0[1]));
    wire [1:0] far_2_2253_1;    relay_conn far_2_2253_1_a(.in(far_2_2253_0[0]), .out(far_2_2253_1[0]));    relay_conn far_2_2253_1_b(.in(far_2_2253_0[1]), .out(far_2_2253_1[1]));
    assign layer_2[213] = ~(far_2_2253_1[0] | far_2_2253_1[1]); 
    assign layer_2[214] = ~layer_1[695]; 
    assign layer_2[215] = layer_1[983] & ~layer_1[972]; 
    assign layer_2[216] = ~(layer_1[814] ^ layer_1[796]); 
    wire [1:0] far_2_2257_0;    relay_conn far_2_2257_0_a(.in(layer_1[765]), .out(far_2_2257_0[0]));    relay_conn far_2_2257_0_b(.in(layer_1[659]), .out(far_2_2257_0[1]));
    wire [1:0] far_2_2257_1;    relay_conn far_2_2257_1_a(.in(far_2_2257_0[0]), .out(far_2_2257_1[0]));    relay_conn far_2_2257_1_b(.in(far_2_2257_0[1]), .out(far_2_2257_1[1]));
    wire [1:0] far_2_2257_2;    relay_conn far_2_2257_2_a(.in(far_2_2257_1[0]), .out(far_2_2257_2[0]));    relay_conn far_2_2257_2_b(.in(far_2_2257_1[1]), .out(far_2_2257_2[1]));
    assign layer_2[217] = far_2_2257_2[1] & ~far_2_2257_2[0]; 
    wire [1:0] far_2_2258_0;    relay_conn far_2_2258_0_a(.in(layer_1[446]), .out(far_2_2258_0[0]));    relay_conn far_2_2258_0_b(.in(layer_1[561]), .out(far_2_2258_0[1]));
    wire [1:0] far_2_2258_1;    relay_conn far_2_2258_1_a(.in(far_2_2258_0[0]), .out(far_2_2258_1[0]));    relay_conn far_2_2258_1_b(.in(far_2_2258_0[1]), .out(far_2_2258_1[1]));
    wire [1:0] far_2_2258_2;    relay_conn far_2_2258_2_a(.in(far_2_2258_1[0]), .out(far_2_2258_2[0]));    relay_conn far_2_2258_2_b(.in(far_2_2258_1[1]), .out(far_2_2258_2[1]));
    assign layer_2[218] = ~far_2_2258_2[1]; 
    wire [1:0] far_2_2259_0;    relay_conn far_2_2259_0_a(.in(layer_1[400]), .out(far_2_2259_0[0]));    relay_conn far_2_2259_0_b(.in(layer_1[522]), .out(far_2_2259_0[1]));
    wire [1:0] far_2_2259_1;    relay_conn far_2_2259_1_a(.in(far_2_2259_0[0]), .out(far_2_2259_1[0]));    relay_conn far_2_2259_1_b(.in(far_2_2259_0[1]), .out(far_2_2259_1[1]));
    wire [1:0] far_2_2259_2;    relay_conn far_2_2259_2_a(.in(far_2_2259_1[0]), .out(far_2_2259_2[0]));    relay_conn far_2_2259_2_b(.in(far_2_2259_1[1]), .out(far_2_2259_2[1]));
    assign layer_2[219] = far_2_2259_2[1]; 
    wire [1:0] far_2_2260_0;    relay_conn far_2_2260_0_a(.in(layer_1[87]), .out(far_2_2260_0[0]));    relay_conn far_2_2260_0_b(.in(layer_1[161]), .out(far_2_2260_0[1]));
    wire [1:0] far_2_2260_1;    relay_conn far_2_2260_1_a(.in(far_2_2260_0[0]), .out(far_2_2260_1[0]));    relay_conn far_2_2260_1_b(.in(far_2_2260_0[1]), .out(far_2_2260_1[1]));
    assign layer_2[220] = far_2_2260_1[0]; 
    assign layer_2[221] = layer_1[795]; 
    wire [1:0] far_2_2262_0;    relay_conn far_2_2262_0_a(.in(layer_1[646]), .out(far_2_2262_0[0]));    relay_conn far_2_2262_0_b(.in(layer_1[771]), .out(far_2_2262_0[1]));
    wire [1:0] far_2_2262_1;    relay_conn far_2_2262_1_a(.in(far_2_2262_0[0]), .out(far_2_2262_1[0]));    relay_conn far_2_2262_1_b(.in(far_2_2262_0[1]), .out(far_2_2262_1[1]));
    wire [1:0] far_2_2262_2;    relay_conn far_2_2262_2_a(.in(far_2_2262_1[0]), .out(far_2_2262_2[0]));    relay_conn far_2_2262_2_b(.in(far_2_2262_1[1]), .out(far_2_2262_2[1]));
    assign layer_2[222] = far_2_2262_2[0] ^ far_2_2262_2[1]; 
    wire [1:0] far_2_2263_0;    relay_conn far_2_2263_0_a(.in(layer_1[102]), .out(far_2_2263_0[0]));    relay_conn far_2_2263_0_b(.in(layer_1[169]), .out(far_2_2263_0[1]));
    wire [1:0] far_2_2263_1;    relay_conn far_2_2263_1_a(.in(far_2_2263_0[0]), .out(far_2_2263_1[0]));    relay_conn far_2_2263_1_b(.in(far_2_2263_0[1]), .out(far_2_2263_1[1]));
    assign layer_2[223] = far_2_2263_1[0] | far_2_2263_1[1]; 
    wire [1:0] far_2_2264_0;    relay_conn far_2_2264_0_a(.in(layer_1[353]), .out(far_2_2264_0[0]));    relay_conn far_2_2264_0_b(.in(layer_1[257]), .out(far_2_2264_0[1]));
    wire [1:0] far_2_2264_1;    relay_conn far_2_2264_1_a(.in(far_2_2264_0[0]), .out(far_2_2264_1[0]));    relay_conn far_2_2264_1_b(.in(far_2_2264_0[1]), .out(far_2_2264_1[1]));
    wire [1:0] far_2_2264_2;    relay_conn far_2_2264_2_a(.in(far_2_2264_1[0]), .out(far_2_2264_2[0]));    relay_conn far_2_2264_2_b(.in(far_2_2264_1[1]), .out(far_2_2264_2[1]));
    assign layer_2[224] = far_2_2264_2[0] ^ far_2_2264_2[1]; 
    wire [1:0] far_2_2265_0;    relay_conn far_2_2265_0_a(.in(layer_1[875]), .out(far_2_2265_0[0]));    relay_conn far_2_2265_0_b(.in(layer_1[757]), .out(far_2_2265_0[1]));
    wire [1:0] far_2_2265_1;    relay_conn far_2_2265_1_a(.in(far_2_2265_0[0]), .out(far_2_2265_1[0]));    relay_conn far_2_2265_1_b(.in(far_2_2265_0[1]), .out(far_2_2265_1[1]));
    wire [1:0] far_2_2265_2;    relay_conn far_2_2265_2_a(.in(far_2_2265_1[0]), .out(far_2_2265_2[0]));    relay_conn far_2_2265_2_b(.in(far_2_2265_1[1]), .out(far_2_2265_2[1]));
    assign layer_2[225] = far_2_2265_2[1]; 
    wire [1:0] far_2_2266_0;    relay_conn far_2_2266_0_a(.in(layer_1[93]), .out(far_2_2266_0[0]));    relay_conn far_2_2266_0_b(.in(layer_1[45]), .out(far_2_2266_0[1]));
    assign layer_2[226] = far_2_2266_0[0]; 
    wire [1:0] far_2_2267_0;    relay_conn far_2_2267_0_a(.in(layer_1[255]), .out(far_2_2267_0[0]));    relay_conn far_2_2267_0_b(.in(layer_1[131]), .out(far_2_2267_0[1]));
    wire [1:0] far_2_2267_1;    relay_conn far_2_2267_1_a(.in(far_2_2267_0[0]), .out(far_2_2267_1[0]));    relay_conn far_2_2267_1_b(.in(far_2_2267_0[1]), .out(far_2_2267_1[1]));
    wire [1:0] far_2_2267_2;    relay_conn far_2_2267_2_a(.in(far_2_2267_1[0]), .out(far_2_2267_2[0]));    relay_conn far_2_2267_2_b(.in(far_2_2267_1[1]), .out(far_2_2267_2[1]));
    assign layer_2[227] = far_2_2267_2[1]; 
    assign layer_2[228] = ~layer_1[867]; 
    wire [1:0] far_2_2269_0;    relay_conn far_2_2269_0_a(.in(layer_1[303]), .out(far_2_2269_0[0]));    relay_conn far_2_2269_0_b(.in(layer_1[239]), .out(far_2_2269_0[1]));
    wire [1:0] far_2_2269_1;    relay_conn far_2_2269_1_a(.in(far_2_2269_0[0]), .out(far_2_2269_1[0]));    relay_conn far_2_2269_1_b(.in(far_2_2269_0[1]), .out(far_2_2269_1[1]));
    assign layer_2[229] = ~(far_2_2269_1[0] | far_2_2269_1[1]); 
    wire [1:0] far_2_2270_0;    relay_conn far_2_2270_0_a(.in(layer_1[965]), .out(far_2_2270_0[0]));    relay_conn far_2_2270_0_b(.in(layer_1[918]), .out(far_2_2270_0[1]));
    assign layer_2[230] = far_2_2270_0[0]; 
    assign layer_2[231] = ~layer_1[810] | (layer_1[810] & layer_1[834]); 
    wire [1:0] far_2_2272_0;    relay_conn far_2_2272_0_a(.in(layer_1[677]), .out(far_2_2272_0[0]));    relay_conn far_2_2272_0_b(.in(layer_1[571]), .out(far_2_2272_0[1]));
    wire [1:0] far_2_2272_1;    relay_conn far_2_2272_1_a(.in(far_2_2272_0[0]), .out(far_2_2272_1[0]));    relay_conn far_2_2272_1_b(.in(far_2_2272_0[1]), .out(far_2_2272_1[1]));
    wire [1:0] far_2_2272_2;    relay_conn far_2_2272_2_a(.in(far_2_2272_1[0]), .out(far_2_2272_2[0]));    relay_conn far_2_2272_2_b(.in(far_2_2272_1[1]), .out(far_2_2272_2[1]));
    assign layer_2[232] = ~far_2_2272_2[1] | (far_2_2272_2[0] & far_2_2272_2[1]); 
    wire [1:0] far_2_2273_0;    relay_conn far_2_2273_0_a(.in(layer_1[27]), .out(far_2_2273_0[0]));    relay_conn far_2_2273_0_b(.in(layer_1[64]), .out(far_2_2273_0[1]));
    assign layer_2[233] = far_2_2273_0[0]; 
    wire [1:0] far_2_2274_0;    relay_conn far_2_2274_0_a(.in(layer_1[685]), .out(far_2_2274_0[0]));    relay_conn far_2_2274_0_b(.in(layer_1[574]), .out(far_2_2274_0[1]));
    wire [1:0] far_2_2274_1;    relay_conn far_2_2274_1_a(.in(far_2_2274_0[0]), .out(far_2_2274_1[0]));    relay_conn far_2_2274_1_b(.in(far_2_2274_0[1]), .out(far_2_2274_1[1]));
    wire [1:0] far_2_2274_2;    relay_conn far_2_2274_2_a(.in(far_2_2274_1[0]), .out(far_2_2274_2[0]));    relay_conn far_2_2274_2_b(.in(far_2_2274_1[1]), .out(far_2_2274_2[1]));
    assign layer_2[234] = far_2_2274_2[1] & ~far_2_2274_2[0]; 
    wire [1:0] far_2_2275_0;    relay_conn far_2_2275_0_a(.in(layer_1[242]), .out(far_2_2275_0[0]));    relay_conn far_2_2275_0_b(.in(layer_1[329]), .out(far_2_2275_0[1]));
    wire [1:0] far_2_2275_1;    relay_conn far_2_2275_1_a(.in(far_2_2275_0[0]), .out(far_2_2275_1[0]));    relay_conn far_2_2275_1_b(.in(far_2_2275_0[1]), .out(far_2_2275_1[1]));
    assign layer_2[235] = far_2_2275_1[0] | far_2_2275_1[1]; 
    wire [1:0] far_2_2276_0;    relay_conn far_2_2276_0_a(.in(layer_1[419]), .out(far_2_2276_0[0]));    relay_conn far_2_2276_0_b(.in(layer_1[482]), .out(far_2_2276_0[1]));
    assign layer_2[236] = far_2_2276_0[1] & ~far_2_2276_0[0]; 
    wire [1:0] far_2_2277_0;    relay_conn far_2_2277_0_a(.in(layer_1[481]), .out(far_2_2277_0[0]));    relay_conn far_2_2277_0_b(.in(layer_1[428]), .out(far_2_2277_0[1]));
    assign layer_2[237] = ~far_2_2277_0[0]; 
    wire [1:0] far_2_2278_0;    relay_conn far_2_2278_0_a(.in(layer_1[795]), .out(far_2_2278_0[0]));    relay_conn far_2_2278_0_b(.in(layer_1[688]), .out(far_2_2278_0[1]));
    wire [1:0] far_2_2278_1;    relay_conn far_2_2278_1_a(.in(far_2_2278_0[0]), .out(far_2_2278_1[0]));    relay_conn far_2_2278_1_b(.in(far_2_2278_0[1]), .out(far_2_2278_1[1]));
    wire [1:0] far_2_2278_2;    relay_conn far_2_2278_2_a(.in(far_2_2278_1[0]), .out(far_2_2278_2[0]));    relay_conn far_2_2278_2_b(.in(far_2_2278_1[1]), .out(far_2_2278_2[1]));
    assign layer_2[238] = far_2_2278_2[1] & ~far_2_2278_2[0]; 
    wire [1:0] far_2_2279_0;    relay_conn far_2_2279_0_a(.in(layer_1[810]), .out(far_2_2279_0[0]));    relay_conn far_2_2279_0_b(.in(layer_1[862]), .out(far_2_2279_0[1]));
    assign layer_2[239] = far_2_2279_0[1]; 
    wire [1:0] far_2_2280_0;    relay_conn far_2_2280_0_a(.in(layer_1[781]), .out(far_2_2280_0[0]));    relay_conn far_2_2280_0_b(.in(layer_1[894]), .out(far_2_2280_0[1]));
    wire [1:0] far_2_2280_1;    relay_conn far_2_2280_1_a(.in(far_2_2280_0[0]), .out(far_2_2280_1[0]));    relay_conn far_2_2280_1_b(.in(far_2_2280_0[1]), .out(far_2_2280_1[1]));
    wire [1:0] far_2_2280_2;    relay_conn far_2_2280_2_a(.in(far_2_2280_1[0]), .out(far_2_2280_2[0]));    relay_conn far_2_2280_2_b(.in(far_2_2280_1[1]), .out(far_2_2280_2[1]));
    assign layer_2[240] = far_2_2280_2[0] & far_2_2280_2[1]; 
    wire [1:0] far_2_2281_0;    relay_conn far_2_2281_0_a(.in(layer_1[162]), .out(far_2_2281_0[0]));    relay_conn far_2_2281_0_b(.in(layer_1[270]), .out(far_2_2281_0[1]));
    wire [1:0] far_2_2281_1;    relay_conn far_2_2281_1_a(.in(far_2_2281_0[0]), .out(far_2_2281_1[0]));    relay_conn far_2_2281_1_b(.in(far_2_2281_0[1]), .out(far_2_2281_1[1]));
    wire [1:0] far_2_2281_2;    relay_conn far_2_2281_2_a(.in(far_2_2281_1[0]), .out(far_2_2281_2[0]));    relay_conn far_2_2281_2_b(.in(far_2_2281_1[1]), .out(far_2_2281_2[1]));
    assign layer_2[241] = ~far_2_2281_2[0]; 
    wire [1:0] far_2_2282_0;    relay_conn far_2_2282_0_a(.in(layer_1[721]), .out(far_2_2282_0[0]));    relay_conn far_2_2282_0_b(.in(layer_1[764]), .out(far_2_2282_0[1]));
    assign layer_2[242] = ~far_2_2282_0[1]; 
    assign layer_2[243] = layer_1[25]; 
    wire [1:0] far_2_2284_0;    relay_conn far_2_2284_0_a(.in(layer_1[1007]), .out(far_2_2284_0[0]));    relay_conn far_2_2284_0_b(.in(layer_1[910]), .out(far_2_2284_0[1]));
    wire [1:0] far_2_2284_1;    relay_conn far_2_2284_1_a(.in(far_2_2284_0[0]), .out(far_2_2284_1[0]));    relay_conn far_2_2284_1_b(.in(far_2_2284_0[1]), .out(far_2_2284_1[1]));
    wire [1:0] far_2_2284_2;    relay_conn far_2_2284_2_a(.in(far_2_2284_1[0]), .out(far_2_2284_2[0]));    relay_conn far_2_2284_2_b(.in(far_2_2284_1[1]), .out(far_2_2284_2[1]));
    assign layer_2[244] = far_2_2284_2[1] & ~far_2_2284_2[0]; 
    wire [1:0] far_2_2285_0;    relay_conn far_2_2285_0_a(.in(layer_1[0]), .out(far_2_2285_0[0]));    relay_conn far_2_2285_0_b(.in(layer_1[107]), .out(far_2_2285_0[1]));
    wire [1:0] far_2_2285_1;    relay_conn far_2_2285_1_a(.in(far_2_2285_0[0]), .out(far_2_2285_1[0]));    relay_conn far_2_2285_1_b(.in(far_2_2285_0[1]), .out(far_2_2285_1[1]));
    wire [1:0] far_2_2285_2;    relay_conn far_2_2285_2_a(.in(far_2_2285_1[0]), .out(far_2_2285_2[0]));    relay_conn far_2_2285_2_b(.in(far_2_2285_1[1]), .out(far_2_2285_2[1]));
    assign layer_2[245] = far_2_2285_2[0]; 
    wire [1:0] far_2_2286_0;    relay_conn far_2_2286_0_a(.in(layer_1[856]), .out(far_2_2286_0[0]));    relay_conn far_2_2286_0_b(.in(layer_1[782]), .out(far_2_2286_0[1]));
    wire [1:0] far_2_2286_1;    relay_conn far_2_2286_1_a(.in(far_2_2286_0[0]), .out(far_2_2286_1[0]));    relay_conn far_2_2286_1_b(.in(far_2_2286_0[1]), .out(far_2_2286_1[1]));
    assign layer_2[246] = ~far_2_2286_1[1]; 
    wire [1:0] far_2_2287_0;    relay_conn far_2_2287_0_a(.in(layer_1[603]), .out(far_2_2287_0[0]));    relay_conn far_2_2287_0_b(.in(layer_1[561]), .out(far_2_2287_0[1]));
    assign layer_2[247] = far_2_2287_0[1] & ~far_2_2287_0[0]; 
    wire [1:0] far_2_2288_0;    relay_conn far_2_2288_0_a(.in(layer_1[558]), .out(far_2_2288_0[0]));    relay_conn far_2_2288_0_b(.in(layer_1[447]), .out(far_2_2288_0[1]));
    wire [1:0] far_2_2288_1;    relay_conn far_2_2288_1_a(.in(far_2_2288_0[0]), .out(far_2_2288_1[0]));    relay_conn far_2_2288_1_b(.in(far_2_2288_0[1]), .out(far_2_2288_1[1]));
    wire [1:0] far_2_2288_2;    relay_conn far_2_2288_2_a(.in(far_2_2288_1[0]), .out(far_2_2288_2[0]));    relay_conn far_2_2288_2_b(.in(far_2_2288_1[1]), .out(far_2_2288_2[1]));
    assign layer_2[248] = ~far_2_2288_2[0] | (far_2_2288_2[0] & far_2_2288_2[1]); 
    assign layer_2[249] = ~(layer_1[813] & layer_1[797]); 
    wire [1:0] far_2_2290_0;    relay_conn far_2_2290_0_a(.in(layer_1[369]), .out(far_2_2290_0[0]));    relay_conn far_2_2290_0_b(.in(layer_1[281]), .out(far_2_2290_0[1]));
    wire [1:0] far_2_2290_1;    relay_conn far_2_2290_1_a(.in(far_2_2290_0[0]), .out(far_2_2290_1[0]));    relay_conn far_2_2290_1_b(.in(far_2_2290_0[1]), .out(far_2_2290_1[1]));
    assign layer_2[250] = ~far_2_2290_1[1] | (far_2_2290_1[0] & far_2_2290_1[1]); 
    assign layer_2[251] = layer_1[724] & ~layer_1[699]; 
    assign layer_2[252] = layer_1[757] & ~layer_1[767]; 
    assign layer_2[253] = ~layer_1[923] | (layer_1[947] & layer_1[923]); 
    wire [1:0] far_2_2294_0;    relay_conn far_2_2294_0_a(.in(layer_1[272]), .out(far_2_2294_0[0]));    relay_conn far_2_2294_0_b(.in(layer_1[371]), .out(far_2_2294_0[1]));
    wire [1:0] far_2_2294_1;    relay_conn far_2_2294_1_a(.in(far_2_2294_0[0]), .out(far_2_2294_1[0]));    relay_conn far_2_2294_1_b(.in(far_2_2294_0[1]), .out(far_2_2294_1[1]));
    wire [1:0] far_2_2294_2;    relay_conn far_2_2294_2_a(.in(far_2_2294_1[0]), .out(far_2_2294_2[0]));    relay_conn far_2_2294_2_b(.in(far_2_2294_1[1]), .out(far_2_2294_2[1]));
    assign layer_2[254] = far_2_2294_2[0] & ~far_2_2294_2[1]; 
    wire [1:0] far_2_2295_0;    relay_conn far_2_2295_0_a(.in(layer_1[665]), .out(far_2_2295_0[0]));    relay_conn far_2_2295_0_b(.in(layer_1[571]), .out(far_2_2295_0[1]));
    wire [1:0] far_2_2295_1;    relay_conn far_2_2295_1_a(.in(far_2_2295_0[0]), .out(far_2_2295_1[0]));    relay_conn far_2_2295_1_b(.in(far_2_2295_0[1]), .out(far_2_2295_1[1]));
    assign layer_2[255] = ~far_2_2295_1[0] | (far_2_2295_1[0] & far_2_2295_1[1]); 
    wire [1:0] far_2_2296_0;    relay_conn far_2_2296_0_a(.in(layer_1[377]), .out(far_2_2296_0[0]));    relay_conn far_2_2296_0_b(.in(layer_1[462]), .out(far_2_2296_0[1]));
    wire [1:0] far_2_2296_1;    relay_conn far_2_2296_1_a(.in(far_2_2296_0[0]), .out(far_2_2296_1[0]));    relay_conn far_2_2296_1_b(.in(far_2_2296_0[1]), .out(far_2_2296_1[1]));
    assign layer_2[256] = far_2_2296_1[1]; 
    assign layer_2[257] = layer_1[854] ^ layer_1[864]; 
    wire [1:0] far_2_2298_0;    relay_conn far_2_2298_0_a(.in(layer_1[180]), .out(far_2_2298_0[0]));    relay_conn far_2_2298_0_b(.in(layer_1[98]), .out(far_2_2298_0[1]));
    wire [1:0] far_2_2298_1;    relay_conn far_2_2298_1_a(.in(far_2_2298_0[0]), .out(far_2_2298_1[0]));    relay_conn far_2_2298_1_b(.in(far_2_2298_0[1]), .out(far_2_2298_1[1]));
    assign layer_2[258] = far_2_2298_1[1] & ~far_2_2298_1[0]; 
    wire [1:0] far_2_2299_0;    relay_conn far_2_2299_0_a(.in(layer_1[854]), .out(far_2_2299_0[0]));    relay_conn far_2_2299_0_b(.in(layer_1[918]), .out(far_2_2299_0[1]));
    wire [1:0] far_2_2299_1;    relay_conn far_2_2299_1_a(.in(far_2_2299_0[0]), .out(far_2_2299_1[0]));    relay_conn far_2_2299_1_b(.in(far_2_2299_0[1]), .out(far_2_2299_1[1]));
    assign layer_2[259] = far_2_2299_1[1]; 
    wire [1:0] far_2_2300_0;    relay_conn far_2_2300_0_a(.in(layer_1[99]), .out(far_2_2300_0[0]));    relay_conn far_2_2300_0_b(.in(layer_1[47]), .out(far_2_2300_0[1]));
    assign layer_2[260] = ~far_2_2300_0[1]; 
    assign layer_2[261] = ~layer_1[212]; 
    assign layer_2[262] = ~(layer_1[913] & layer_1[897]); 
    wire [1:0] far_2_2303_0;    relay_conn far_2_2303_0_a(.in(layer_1[783]), .out(far_2_2303_0[0]));    relay_conn far_2_2303_0_b(.in(layer_1[846]), .out(far_2_2303_0[1]));
    assign layer_2[263] = ~(far_2_2303_0[0] | far_2_2303_0[1]); 
    wire [1:0] far_2_2304_0;    relay_conn far_2_2304_0_a(.in(layer_1[125]), .out(far_2_2304_0[0]));    relay_conn far_2_2304_0_b(.in(layer_1[57]), .out(far_2_2304_0[1]));
    wire [1:0] far_2_2304_1;    relay_conn far_2_2304_1_a(.in(far_2_2304_0[0]), .out(far_2_2304_1[0]));    relay_conn far_2_2304_1_b(.in(far_2_2304_0[1]), .out(far_2_2304_1[1]));
    assign layer_2[264] = far_2_2304_1[0]; 
    wire [1:0] far_2_2305_0;    relay_conn far_2_2305_0_a(.in(layer_1[966]), .out(far_2_2305_0[0]));    relay_conn far_2_2305_0_b(.in(layer_1[846]), .out(far_2_2305_0[1]));
    wire [1:0] far_2_2305_1;    relay_conn far_2_2305_1_a(.in(far_2_2305_0[0]), .out(far_2_2305_1[0]));    relay_conn far_2_2305_1_b(.in(far_2_2305_0[1]), .out(far_2_2305_1[1]));
    wire [1:0] far_2_2305_2;    relay_conn far_2_2305_2_a(.in(far_2_2305_1[0]), .out(far_2_2305_2[0]));    relay_conn far_2_2305_2_b(.in(far_2_2305_1[1]), .out(far_2_2305_2[1]));
    assign layer_2[265] = ~far_2_2305_2[1]; 
    wire [1:0] far_2_2306_0;    relay_conn far_2_2306_0_a(.in(layer_1[858]), .out(far_2_2306_0[0]));    relay_conn far_2_2306_0_b(.in(layer_1[749]), .out(far_2_2306_0[1]));
    wire [1:0] far_2_2306_1;    relay_conn far_2_2306_1_a(.in(far_2_2306_0[0]), .out(far_2_2306_1[0]));    relay_conn far_2_2306_1_b(.in(far_2_2306_0[1]), .out(far_2_2306_1[1]));
    wire [1:0] far_2_2306_2;    relay_conn far_2_2306_2_a(.in(far_2_2306_1[0]), .out(far_2_2306_2[0]));    relay_conn far_2_2306_2_b(.in(far_2_2306_1[1]), .out(far_2_2306_2[1]));
    assign layer_2[266] = ~far_2_2306_2[1]; 
    wire [1:0] far_2_2307_0;    relay_conn far_2_2307_0_a(.in(layer_1[455]), .out(far_2_2307_0[0]));    relay_conn far_2_2307_0_b(.in(layer_1[410]), .out(far_2_2307_0[1]));
    assign layer_2[267] = far_2_2307_0[0] & ~far_2_2307_0[1]; 
    wire [1:0] far_2_2308_0;    relay_conn far_2_2308_0_a(.in(layer_1[169]), .out(far_2_2308_0[0]));    relay_conn far_2_2308_0_b(.in(layer_1[87]), .out(far_2_2308_0[1]));
    wire [1:0] far_2_2308_1;    relay_conn far_2_2308_1_a(.in(far_2_2308_0[0]), .out(far_2_2308_1[0]));    relay_conn far_2_2308_1_b(.in(far_2_2308_0[1]), .out(far_2_2308_1[1]));
    assign layer_2[268] = far_2_2308_1[1] & ~far_2_2308_1[0]; 
    wire [1:0] far_2_2309_0;    relay_conn far_2_2309_0_a(.in(layer_1[932]), .out(far_2_2309_0[0]));    relay_conn far_2_2309_0_b(.in(layer_1[810]), .out(far_2_2309_0[1]));
    wire [1:0] far_2_2309_1;    relay_conn far_2_2309_1_a(.in(far_2_2309_0[0]), .out(far_2_2309_1[0]));    relay_conn far_2_2309_1_b(.in(far_2_2309_0[1]), .out(far_2_2309_1[1]));
    wire [1:0] far_2_2309_2;    relay_conn far_2_2309_2_a(.in(far_2_2309_1[0]), .out(far_2_2309_2[0]));    relay_conn far_2_2309_2_b(.in(far_2_2309_1[1]), .out(far_2_2309_2[1]));
    assign layer_2[269] = far_2_2309_2[0] | far_2_2309_2[1]; 
    wire [1:0] far_2_2310_0;    relay_conn far_2_2310_0_a(.in(layer_1[643]), .out(far_2_2310_0[0]));    relay_conn far_2_2310_0_b(.in(layer_1[559]), .out(far_2_2310_0[1]));
    wire [1:0] far_2_2310_1;    relay_conn far_2_2310_1_a(.in(far_2_2310_0[0]), .out(far_2_2310_1[0]));    relay_conn far_2_2310_1_b(.in(far_2_2310_0[1]), .out(far_2_2310_1[1]));
    assign layer_2[270] = far_2_2310_1[0] | far_2_2310_1[1]; 
    wire [1:0] far_2_2311_0;    relay_conn far_2_2311_0_a(.in(layer_1[743]), .out(far_2_2311_0[0]));    relay_conn far_2_2311_0_b(.in(layer_1[795]), .out(far_2_2311_0[1]));
    assign layer_2[271] = ~(far_2_2311_0[0] & far_2_2311_0[1]); 
    wire [1:0] far_2_2312_0;    relay_conn far_2_2312_0_a(.in(layer_1[991]), .out(far_2_2312_0[0]));    relay_conn far_2_2312_0_b(.in(layer_1[864]), .out(far_2_2312_0[1]));
    wire [1:0] far_2_2312_1;    relay_conn far_2_2312_1_a(.in(far_2_2312_0[0]), .out(far_2_2312_1[0]));    relay_conn far_2_2312_1_b(.in(far_2_2312_0[1]), .out(far_2_2312_1[1]));
    wire [1:0] far_2_2312_2;    relay_conn far_2_2312_2_a(.in(far_2_2312_1[0]), .out(far_2_2312_2[0]));    relay_conn far_2_2312_2_b(.in(far_2_2312_1[1]), .out(far_2_2312_2[1]));
    assign layer_2[272] = ~(far_2_2312_2[0] ^ far_2_2312_2[1]); 
    wire [1:0] far_2_2313_0;    relay_conn far_2_2313_0_a(.in(layer_1[962]), .out(far_2_2313_0[0]));    relay_conn far_2_2313_0_b(.in(layer_1[927]), .out(far_2_2313_0[1]));
    assign layer_2[273] = ~far_2_2313_0[1] | (far_2_2313_0[0] & far_2_2313_0[1]); 
    assign layer_2[274] = ~(layer_1[934] ^ layer_1[924]); 
    wire [1:0] far_2_2315_0;    relay_conn far_2_2315_0_a(.in(layer_1[814]), .out(far_2_2315_0[0]));    relay_conn far_2_2315_0_b(.in(layer_1[772]), .out(far_2_2315_0[1]));
    assign layer_2[275] = far_2_2315_0[0] | far_2_2315_0[1]; 
    assign layer_2[276] = layer_1[919] | layer_1[897]; 
    wire [1:0] far_2_2317_0;    relay_conn far_2_2317_0_a(.in(layer_1[158]), .out(far_2_2317_0[0]));    relay_conn far_2_2317_0_b(.in(layer_1[95]), .out(far_2_2317_0[1]));
    assign layer_2[277] = ~far_2_2317_0[0]; 
    assign layer_2[278] = layer_1[932]; 
    wire [1:0] far_2_2319_0;    relay_conn far_2_2319_0_a(.in(layer_1[169]), .out(far_2_2319_0[0]));    relay_conn far_2_2319_0_b(.in(layer_1[204]), .out(far_2_2319_0[1]));
    assign layer_2[279] = far_2_2319_0[0] & far_2_2319_0[1]; 
    assign layer_2[280] = ~(layer_1[109] & layer_1[84]); 
    wire [1:0] far_2_2321_0;    relay_conn far_2_2321_0_a(.in(layer_1[595]), .out(far_2_2321_0[0]));    relay_conn far_2_2321_0_b(.in(layer_1[690]), .out(far_2_2321_0[1]));
    wire [1:0] far_2_2321_1;    relay_conn far_2_2321_1_a(.in(far_2_2321_0[0]), .out(far_2_2321_1[0]));    relay_conn far_2_2321_1_b(.in(far_2_2321_0[1]), .out(far_2_2321_1[1]));
    assign layer_2[281] = ~(far_2_2321_1[0] ^ far_2_2321_1[1]); 
    wire [1:0] far_2_2322_0;    relay_conn far_2_2322_0_a(.in(layer_1[854]), .out(far_2_2322_0[0]));    relay_conn far_2_2322_0_b(.in(layer_1[777]), .out(far_2_2322_0[1]));
    wire [1:0] far_2_2322_1;    relay_conn far_2_2322_1_a(.in(far_2_2322_0[0]), .out(far_2_2322_1[0]));    relay_conn far_2_2322_1_b(.in(far_2_2322_0[1]), .out(far_2_2322_1[1]));
    assign layer_2[282] = ~(far_2_2322_1[0] | far_2_2322_1[1]); 
    wire [1:0] far_2_2323_0;    relay_conn far_2_2323_0_a(.in(layer_1[876]), .out(far_2_2323_0[0]));    relay_conn far_2_2323_0_b(.in(layer_1[811]), .out(far_2_2323_0[1]));
    wire [1:0] far_2_2323_1;    relay_conn far_2_2323_1_a(.in(far_2_2323_0[0]), .out(far_2_2323_1[0]));    relay_conn far_2_2323_1_b(.in(far_2_2323_0[1]), .out(far_2_2323_1[1]));
    assign layer_2[283] = far_2_2323_1[0]; 
    wire [1:0] far_2_2324_0;    relay_conn far_2_2324_0_a(.in(layer_1[866]), .out(far_2_2324_0[0]));    relay_conn far_2_2324_0_b(.in(layer_1[946]), .out(far_2_2324_0[1]));
    wire [1:0] far_2_2324_1;    relay_conn far_2_2324_1_a(.in(far_2_2324_0[0]), .out(far_2_2324_1[0]));    relay_conn far_2_2324_1_b(.in(far_2_2324_0[1]), .out(far_2_2324_1[1]));
    assign layer_2[284] = ~far_2_2324_1[1]; 
    wire [1:0] far_2_2325_0;    relay_conn far_2_2325_0_a(.in(layer_1[980]), .out(far_2_2325_0[0]));    relay_conn far_2_2325_0_b(.in(layer_1[864]), .out(far_2_2325_0[1]));
    wire [1:0] far_2_2325_1;    relay_conn far_2_2325_1_a(.in(far_2_2325_0[0]), .out(far_2_2325_1[0]));    relay_conn far_2_2325_1_b(.in(far_2_2325_0[1]), .out(far_2_2325_1[1]));
    wire [1:0] far_2_2325_2;    relay_conn far_2_2325_2_a(.in(far_2_2325_1[0]), .out(far_2_2325_2[0]));    relay_conn far_2_2325_2_b(.in(far_2_2325_1[1]), .out(far_2_2325_2[1]));
    assign layer_2[285] = ~far_2_2325_2[1]; 
    wire [1:0] far_2_2326_0;    relay_conn far_2_2326_0_a(.in(layer_1[353]), .out(far_2_2326_0[0]));    relay_conn far_2_2326_0_b(.in(layer_1[280]), .out(far_2_2326_0[1]));
    wire [1:0] far_2_2326_1;    relay_conn far_2_2326_1_a(.in(far_2_2326_0[0]), .out(far_2_2326_1[0]));    relay_conn far_2_2326_1_b(.in(far_2_2326_0[1]), .out(far_2_2326_1[1]));
    assign layer_2[286] = ~(far_2_2326_1[0] & far_2_2326_1[1]); 
    wire [1:0] far_2_2327_0;    relay_conn far_2_2327_0_a(.in(layer_1[359]), .out(far_2_2327_0[0]));    relay_conn far_2_2327_0_b(.in(layer_1[284]), .out(far_2_2327_0[1]));
    wire [1:0] far_2_2327_1;    relay_conn far_2_2327_1_a(.in(far_2_2327_0[0]), .out(far_2_2327_1[0]));    relay_conn far_2_2327_1_b(.in(far_2_2327_0[1]), .out(far_2_2327_1[1]));
    assign layer_2[287] = ~far_2_2327_1[1]; 
    wire [1:0] far_2_2328_0;    relay_conn far_2_2328_0_a(.in(layer_1[692]), .out(far_2_2328_0[0]));    relay_conn far_2_2328_0_b(.in(layer_1[757]), .out(far_2_2328_0[1]));
    wire [1:0] far_2_2328_1;    relay_conn far_2_2328_1_a(.in(far_2_2328_0[0]), .out(far_2_2328_1[0]));    relay_conn far_2_2328_1_b(.in(far_2_2328_0[1]), .out(far_2_2328_1[1]));
    assign layer_2[288] = ~(far_2_2328_1[0] | far_2_2328_1[1]); 
    wire [1:0] far_2_2329_0;    relay_conn far_2_2329_0_a(.in(layer_1[340]), .out(far_2_2329_0[0]));    relay_conn far_2_2329_0_b(.in(layer_1[456]), .out(far_2_2329_0[1]));
    wire [1:0] far_2_2329_1;    relay_conn far_2_2329_1_a(.in(far_2_2329_0[0]), .out(far_2_2329_1[0]));    relay_conn far_2_2329_1_b(.in(far_2_2329_0[1]), .out(far_2_2329_1[1]));
    wire [1:0] far_2_2329_2;    relay_conn far_2_2329_2_a(.in(far_2_2329_1[0]), .out(far_2_2329_2[0]));    relay_conn far_2_2329_2_b(.in(far_2_2329_1[1]), .out(far_2_2329_2[1]));
    assign layer_2[289] = ~(far_2_2329_2[0] & far_2_2329_2[1]); 
    assign layer_2[290] = layer_1[292] & ~layer_1[309]; 
    wire [1:0] far_2_2331_0;    relay_conn far_2_2331_0_a(.in(layer_1[967]), .out(far_2_2331_0[0]));    relay_conn far_2_2331_0_b(.in(layer_1[864]), .out(far_2_2331_0[1]));
    wire [1:0] far_2_2331_1;    relay_conn far_2_2331_1_a(.in(far_2_2331_0[0]), .out(far_2_2331_1[0]));    relay_conn far_2_2331_1_b(.in(far_2_2331_0[1]), .out(far_2_2331_1[1]));
    wire [1:0] far_2_2331_2;    relay_conn far_2_2331_2_a(.in(far_2_2331_1[0]), .out(far_2_2331_2[0]));    relay_conn far_2_2331_2_b(.in(far_2_2331_1[1]), .out(far_2_2331_2[1]));
    assign layer_2[291] = far_2_2331_2[0] ^ far_2_2331_2[1]; 
    wire [1:0] far_2_2332_0;    relay_conn far_2_2332_0_a(.in(layer_1[358]), .out(far_2_2332_0[0]));    relay_conn far_2_2332_0_b(.in(layer_1[303]), .out(far_2_2332_0[1]));
    assign layer_2[292] = ~(far_2_2332_0[0] | far_2_2332_0[1]); 
    wire [1:0] far_2_2333_0;    relay_conn far_2_2333_0_a(.in(layer_1[477]), .out(far_2_2333_0[0]));    relay_conn far_2_2333_0_b(.in(layer_1[537]), .out(far_2_2333_0[1]));
    assign layer_2[293] = far_2_2333_0[0] | far_2_2333_0[1]; 
    wire [1:0] far_2_2334_0;    relay_conn far_2_2334_0_a(.in(layer_1[1008]), .out(far_2_2334_0[0]));    relay_conn far_2_2334_0_b(.in(layer_1[966]), .out(far_2_2334_0[1]));
    assign layer_2[294] = ~(far_2_2334_0[0] | far_2_2334_0[1]); 
    wire [1:0] far_2_2335_0;    relay_conn far_2_2335_0_a(.in(layer_1[965]), .out(far_2_2335_0[0]));    relay_conn far_2_2335_0_b(.in(layer_1[932]), .out(far_2_2335_0[1]));
    assign layer_2[295] = ~(far_2_2335_0[0] | far_2_2335_0[1]); 
    wire [1:0] far_2_2336_0;    relay_conn far_2_2336_0_a(.in(layer_1[796]), .out(far_2_2336_0[0]));    relay_conn far_2_2336_0_b(.in(layer_1[902]), .out(far_2_2336_0[1]));
    wire [1:0] far_2_2336_1;    relay_conn far_2_2336_1_a(.in(far_2_2336_0[0]), .out(far_2_2336_1[0]));    relay_conn far_2_2336_1_b(.in(far_2_2336_0[1]), .out(far_2_2336_1[1]));
    wire [1:0] far_2_2336_2;    relay_conn far_2_2336_2_a(.in(far_2_2336_1[0]), .out(far_2_2336_2[0]));    relay_conn far_2_2336_2_b(.in(far_2_2336_1[1]), .out(far_2_2336_2[1]));
    assign layer_2[296] = ~far_2_2336_2[1]; 
    assign layer_2[297] = ~(layer_1[241] | layer_1[215]); 
    wire [1:0] far_2_2338_0;    relay_conn far_2_2338_0_a(.in(layer_1[338]), .out(far_2_2338_0[0]));    relay_conn far_2_2338_0_b(.in(layer_1[458]), .out(far_2_2338_0[1]));
    wire [1:0] far_2_2338_1;    relay_conn far_2_2338_1_a(.in(far_2_2338_0[0]), .out(far_2_2338_1[0]));    relay_conn far_2_2338_1_b(.in(far_2_2338_0[1]), .out(far_2_2338_1[1]));
    wire [1:0] far_2_2338_2;    relay_conn far_2_2338_2_a(.in(far_2_2338_1[0]), .out(far_2_2338_2[0]));    relay_conn far_2_2338_2_b(.in(far_2_2338_1[1]), .out(far_2_2338_2[1]));
    assign layer_2[298] = far_2_2338_2[0] | far_2_2338_2[1]; 
    wire [1:0] far_2_2339_0;    relay_conn far_2_2339_0_a(.in(layer_1[244]), .out(far_2_2339_0[0]));    relay_conn far_2_2339_0_b(.in(layer_1[196]), .out(far_2_2339_0[1]));
    assign layer_2[299] = ~(far_2_2339_0[0] | far_2_2339_0[1]); 
    assign layer_2[300] = layer_1[555] & layer_1[578]; 
    wire [1:0] far_2_2341_0;    relay_conn far_2_2341_0_a(.in(layer_1[215]), .out(far_2_2341_0[0]));    relay_conn far_2_2341_0_b(.in(layer_1[291]), .out(far_2_2341_0[1]));
    wire [1:0] far_2_2341_1;    relay_conn far_2_2341_1_a(.in(far_2_2341_0[0]), .out(far_2_2341_1[0]));    relay_conn far_2_2341_1_b(.in(far_2_2341_0[1]), .out(far_2_2341_1[1]));
    assign layer_2[301] = ~(far_2_2341_1[0] ^ far_2_2341_1[1]); 
    wire [1:0] far_2_2342_0;    relay_conn far_2_2342_0_a(.in(layer_1[745]), .out(far_2_2342_0[0]));    relay_conn far_2_2342_0_b(.in(layer_1[784]), .out(far_2_2342_0[1]));
    assign layer_2[302] = far_2_2342_0[0] & far_2_2342_0[1]; 
    assign layer_2[303] = layer_1[118] & layer_1[103]; 
    assign layer_2[304] = ~layer_1[991] | (layer_1[991] & layer_1[987]); 
    wire [1:0] far_2_2345_0;    relay_conn far_2_2345_0_a(.in(layer_1[186]), .out(far_2_2345_0[0]));    relay_conn far_2_2345_0_b(.in(layer_1[303]), .out(far_2_2345_0[1]));
    wire [1:0] far_2_2345_1;    relay_conn far_2_2345_1_a(.in(far_2_2345_0[0]), .out(far_2_2345_1[0]));    relay_conn far_2_2345_1_b(.in(far_2_2345_0[1]), .out(far_2_2345_1[1]));
    wire [1:0] far_2_2345_2;    relay_conn far_2_2345_2_a(.in(far_2_2345_1[0]), .out(far_2_2345_2[0]));    relay_conn far_2_2345_2_b(.in(far_2_2345_1[1]), .out(far_2_2345_2[1]));
    assign layer_2[305] = far_2_2345_2[0] & far_2_2345_2[1]; 
    wire [1:0] far_2_2346_0;    relay_conn far_2_2346_0_a(.in(layer_1[542]), .out(far_2_2346_0[0]));    relay_conn far_2_2346_0_b(.in(layer_1[654]), .out(far_2_2346_0[1]));
    wire [1:0] far_2_2346_1;    relay_conn far_2_2346_1_a(.in(far_2_2346_0[0]), .out(far_2_2346_1[0]));    relay_conn far_2_2346_1_b(.in(far_2_2346_0[1]), .out(far_2_2346_1[1]));
    wire [1:0] far_2_2346_2;    relay_conn far_2_2346_2_a(.in(far_2_2346_1[0]), .out(far_2_2346_2[0]));    relay_conn far_2_2346_2_b(.in(far_2_2346_1[1]), .out(far_2_2346_2[1]));
    assign layer_2[306] = far_2_2346_2[0]; 
    wire [1:0] far_2_2347_0;    relay_conn far_2_2347_0_a(.in(layer_1[855]), .out(far_2_2347_0[0]));    relay_conn far_2_2347_0_b(.in(layer_1[935]), .out(far_2_2347_0[1]));
    wire [1:0] far_2_2347_1;    relay_conn far_2_2347_1_a(.in(far_2_2347_0[0]), .out(far_2_2347_1[0]));    relay_conn far_2_2347_1_b(.in(far_2_2347_0[1]), .out(far_2_2347_1[1]));
    assign layer_2[307] = far_2_2347_1[0] | far_2_2347_1[1]; 
    assign layer_2[308] = layer_1[746] & ~layer_1[717]; 
    wire [1:0] far_2_2349_0;    relay_conn far_2_2349_0_a(.in(layer_1[87]), .out(far_2_2349_0[0]));    relay_conn far_2_2349_0_b(.in(layer_1[11]), .out(far_2_2349_0[1]));
    wire [1:0] far_2_2349_1;    relay_conn far_2_2349_1_a(.in(far_2_2349_0[0]), .out(far_2_2349_1[0]));    relay_conn far_2_2349_1_b(.in(far_2_2349_0[1]), .out(far_2_2349_1[1]));
    assign layer_2[309] = far_2_2349_1[0] & far_2_2349_1[1]; 
    wire [1:0] far_2_2350_0;    relay_conn far_2_2350_0_a(.in(layer_1[671]), .out(far_2_2350_0[0]));    relay_conn far_2_2350_0_b(.in(layer_1[569]), .out(far_2_2350_0[1]));
    wire [1:0] far_2_2350_1;    relay_conn far_2_2350_1_a(.in(far_2_2350_0[0]), .out(far_2_2350_1[0]));    relay_conn far_2_2350_1_b(.in(far_2_2350_0[1]), .out(far_2_2350_1[1]));
    wire [1:0] far_2_2350_2;    relay_conn far_2_2350_2_a(.in(far_2_2350_1[0]), .out(far_2_2350_2[0]));    relay_conn far_2_2350_2_b(.in(far_2_2350_1[1]), .out(far_2_2350_2[1]));
    assign layer_2[310] = far_2_2350_2[0] & far_2_2350_2[1]; 
    wire [1:0] far_2_2351_0;    relay_conn far_2_2351_0_a(.in(layer_1[836]), .out(far_2_2351_0[0]));    relay_conn far_2_2351_0_b(.in(layer_1[743]), .out(far_2_2351_0[1]));
    wire [1:0] far_2_2351_1;    relay_conn far_2_2351_1_a(.in(far_2_2351_0[0]), .out(far_2_2351_1[0]));    relay_conn far_2_2351_1_b(.in(far_2_2351_0[1]), .out(far_2_2351_1[1]));
    assign layer_2[311] = far_2_2351_1[0] & far_2_2351_1[1]; 
    wire [1:0] far_2_2352_0;    relay_conn far_2_2352_0_a(.in(layer_1[190]), .out(far_2_2352_0[0]));    relay_conn far_2_2352_0_b(.in(layer_1[280]), .out(far_2_2352_0[1]));
    wire [1:0] far_2_2352_1;    relay_conn far_2_2352_1_a(.in(far_2_2352_0[0]), .out(far_2_2352_1[0]));    relay_conn far_2_2352_1_b(.in(far_2_2352_0[1]), .out(far_2_2352_1[1]));
    assign layer_2[312] = ~far_2_2352_1[1] | (far_2_2352_1[0] & far_2_2352_1[1]); 
    wire [1:0] far_2_2353_0;    relay_conn far_2_2353_0_a(.in(layer_1[705]), .out(far_2_2353_0[0]));    relay_conn far_2_2353_0_b(.in(layer_1[795]), .out(far_2_2353_0[1]));
    wire [1:0] far_2_2353_1;    relay_conn far_2_2353_1_a(.in(far_2_2353_0[0]), .out(far_2_2353_1[0]));    relay_conn far_2_2353_1_b(.in(far_2_2353_0[1]), .out(far_2_2353_1[1]));
    assign layer_2[313] = ~far_2_2353_1[0] | (far_2_2353_1[0] & far_2_2353_1[1]); 
    assign layer_2[314] = layer_1[393] & layer_1[404]; 
    assign layer_2[315] = ~layer_1[32]; 
    wire [1:0] far_2_2356_0;    relay_conn far_2_2356_0_a(.in(layer_1[596]), .out(far_2_2356_0[0]));    relay_conn far_2_2356_0_b(.in(layer_1[671]), .out(far_2_2356_0[1]));
    wire [1:0] far_2_2356_1;    relay_conn far_2_2356_1_a(.in(far_2_2356_0[0]), .out(far_2_2356_1[0]));    relay_conn far_2_2356_1_b(.in(far_2_2356_0[1]), .out(far_2_2356_1[1]));
    assign layer_2[316] = ~(far_2_2356_1[0] ^ far_2_2356_1[1]); 
    assign layer_2[317] = ~layer_1[492] | (layer_1[467] & layer_1[492]); 
    wire [1:0] far_2_2358_0;    relay_conn far_2_2358_0_a(.in(layer_1[167]), .out(far_2_2358_0[0]));    relay_conn far_2_2358_0_b(.in(layer_1[86]), .out(far_2_2358_0[1]));
    wire [1:0] far_2_2358_1;    relay_conn far_2_2358_1_a(.in(far_2_2358_0[0]), .out(far_2_2358_1[0]));    relay_conn far_2_2358_1_b(.in(far_2_2358_0[1]), .out(far_2_2358_1[1]));
    assign layer_2[318] = ~(far_2_2358_1[0] & far_2_2358_1[1]); 
    wire [1:0] far_2_2359_0;    relay_conn far_2_2359_0_a(.in(layer_1[637]), .out(far_2_2359_0[0]));    relay_conn far_2_2359_0_b(.in(layer_1[746]), .out(far_2_2359_0[1]));
    wire [1:0] far_2_2359_1;    relay_conn far_2_2359_1_a(.in(far_2_2359_0[0]), .out(far_2_2359_1[0]));    relay_conn far_2_2359_1_b(.in(far_2_2359_0[1]), .out(far_2_2359_1[1]));
    wire [1:0] far_2_2359_2;    relay_conn far_2_2359_2_a(.in(far_2_2359_1[0]), .out(far_2_2359_2[0]));    relay_conn far_2_2359_2_b(.in(far_2_2359_1[1]), .out(far_2_2359_2[1]));
    assign layer_2[319] = far_2_2359_2[0]; 
    assign layer_2[320] = ~layer_1[622] | (layer_1[622] & layer_1[620]); 
    wire [1:0] far_2_2361_0;    relay_conn far_2_2361_0_a(.in(layer_1[66]), .out(far_2_2361_0[0]));    relay_conn far_2_2361_0_b(.in(layer_1[2]), .out(far_2_2361_0[1]));
    wire [1:0] far_2_2361_1;    relay_conn far_2_2361_1_a(.in(far_2_2361_0[0]), .out(far_2_2361_1[0]));    relay_conn far_2_2361_1_b(.in(far_2_2361_0[1]), .out(far_2_2361_1[1]));
    assign layer_2[321] = ~far_2_2361_1[0]; 
    wire [1:0] far_2_2362_0;    relay_conn far_2_2362_0_a(.in(layer_1[763]), .out(far_2_2362_0[0]));    relay_conn far_2_2362_0_b(.in(layer_1[846]), .out(far_2_2362_0[1]));
    wire [1:0] far_2_2362_1;    relay_conn far_2_2362_1_a(.in(far_2_2362_0[0]), .out(far_2_2362_1[0]));    relay_conn far_2_2362_1_b(.in(far_2_2362_0[1]), .out(far_2_2362_1[1]));
    assign layer_2[322] = far_2_2362_1[0] | far_2_2362_1[1]; 
    wire [1:0] far_2_2363_0;    relay_conn far_2_2363_0_a(.in(layer_1[1012]), .out(far_2_2363_0[0]));    relay_conn far_2_2363_0_b(.in(layer_1[966]), .out(far_2_2363_0[1]));
    assign layer_2[323] = far_2_2363_0[1]; 
    wire [1:0] far_2_2364_0;    relay_conn far_2_2364_0_a(.in(layer_1[780]), .out(far_2_2364_0[0]));    relay_conn far_2_2364_0_b(.in(layer_1[695]), .out(far_2_2364_0[1]));
    wire [1:0] far_2_2364_1;    relay_conn far_2_2364_1_a(.in(far_2_2364_0[0]), .out(far_2_2364_1[0]));    relay_conn far_2_2364_1_b(.in(far_2_2364_0[1]), .out(far_2_2364_1[1]));
    assign layer_2[324] = far_2_2364_1[0]; 
    wire [1:0] far_2_2365_0;    relay_conn far_2_2365_0_a(.in(layer_1[561]), .out(far_2_2365_0[0]));    relay_conn far_2_2365_0_b(.in(layer_1[505]), .out(far_2_2365_0[1]));
    assign layer_2[325] = far_2_2365_0[0] & far_2_2365_0[1]; 
    wire [1:0] far_2_2366_0;    relay_conn far_2_2366_0_a(.in(layer_1[405]), .out(far_2_2366_0[0]));    relay_conn far_2_2366_0_b(.in(layer_1[329]), .out(far_2_2366_0[1]));
    wire [1:0] far_2_2366_1;    relay_conn far_2_2366_1_a(.in(far_2_2366_0[0]), .out(far_2_2366_1[0]));    relay_conn far_2_2366_1_b(.in(far_2_2366_0[1]), .out(far_2_2366_1[1]));
    assign layer_2[326] = far_2_2366_1[0] | far_2_2366_1[1]; 
    assign layer_2[327] = ~layer_1[908] | (layer_1[927] & layer_1[908]); 
    wire [1:0] far_2_2368_0;    relay_conn far_2_2368_0_a(.in(layer_1[796]), .out(far_2_2368_0[0]));    relay_conn far_2_2368_0_b(.in(layer_1[711]), .out(far_2_2368_0[1]));
    wire [1:0] far_2_2368_1;    relay_conn far_2_2368_1_a(.in(far_2_2368_0[0]), .out(far_2_2368_1[0]));    relay_conn far_2_2368_1_b(.in(far_2_2368_0[1]), .out(far_2_2368_1[1]));
    assign layer_2[328] = ~(far_2_2368_1[0] | far_2_2368_1[1]); 
    wire [1:0] far_2_2369_0;    relay_conn far_2_2369_0_a(.in(layer_1[93]), .out(far_2_2369_0[0]));    relay_conn far_2_2369_0_b(.in(layer_1[9]), .out(far_2_2369_0[1]));
    wire [1:0] far_2_2369_1;    relay_conn far_2_2369_1_a(.in(far_2_2369_0[0]), .out(far_2_2369_1[0]));    relay_conn far_2_2369_1_b(.in(far_2_2369_0[1]), .out(far_2_2369_1[1]));
    assign layer_2[329] = ~far_2_2369_1[1] | (far_2_2369_1[0] & far_2_2369_1[1]); 
    assign layer_2[330] = layer_1[7] & layer_1[34]; 
    wire [1:0] far_2_2371_0;    relay_conn far_2_2371_0_a(.in(layer_1[303]), .out(far_2_2371_0[0]));    relay_conn far_2_2371_0_b(.in(layer_1[253]), .out(far_2_2371_0[1]));
    assign layer_2[331] = ~(far_2_2371_0[0] ^ far_2_2371_0[1]); 
    wire [1:0] far_2_2372_0;    relay_conn far_2_2372_0_a(.in(layer_1[784]), .out(far_2_2372_0[0]));    relay_conn far_2_2372_0_b(.in(layer_1[866]), .out(far_2_2372_0[1]));
    wire [1:0] far_2_2372_1;    relay_conn far_2_2372_1_a(.in(far_2_2372_0[0]), .out(far_2_2372_1[0]));    relay_conn far_2_2372_1_b(.in(far_2_2372_0[1]), .out(far_2_2372_1[1]));
    assign layer_2[332] = ~far_2_2372_1[0] | (far_2_2372_1[0] & far_2_2372_1[1]); 
    assign layer_2[333] = ~layer_1[46] | (layer_1[47] & layer_1[46]); 
    wire [1:0] far_2_2374_0;    relay_conn far_2_2374_0_a(.in(layer_1[749]), .out(far_2_2374_0[0]));    relay_conn far_2_2374_0_b(.in(layer_1[663]), .out(far_2_2374_0[1]));
    wire [1:0] far_2_2374_1;    relay_conn far_2_2374_1_a(.in(far_2_2374_0[0]), .out(far_2_2374_1[0]));    relay_conn far_2_2374_1_b(.in(far_2_2374_0[1]), .out(far_2_2374_1[1]));
    assign layer_2[334] = far_2_2374_1[0] & far_2_2374_1[1]; 
    wire [1:0] far_2_2375_0;    relay_conn far_2_2375_0_a(.in(layer_1[955]), .out(far_2_2375_0[0]));    relay_conn far_2_2375_0_b(.in(layer_1[832]), .out(far_2_2375_0[1]));
    wire [1:0] far_2_2375_1;    relay_conn far_2_2375_1_a(.in(far_2_2375_0[0]), .out(far_2_2375_1[0]));    relay_conn far_2_2375_1_b(.in(far_2_2375_0[1]), .out(far_2_2375_1[1]));
    wire [1:0] far_2_2375_2;    relay_conn far_2_2375_2_a(.in(far_2_2375_1[0]), .out(far_2_2375_2[0]));    relay_conn far_2_2375_2_b(.in(far_2_2375_1[1]), .out(far_2_2375_2[1]));
    assign layer_2[335] = far_2_2375_2[0] & ~far_2_2375_2[1]; 
    assign layer_2[336] = ~layer_1[639] | (layer_1[619] & layer_1[639]); 
    wire [1:0] far_2_2377_0;    relay_conn far_2_2377_0_a(.in(layer_1[317]), .out(far_2_2377_0[0]));    relay_conn far_2_2377_0_b(.in(layer_1[248]), .out(far_2_2377_0[1]));
    wire [1:0] far_2_2377_1;    relay_conn far_2_2377_1_a(.in(far_2_2377_0[0]), .out(far_2_2377_1[0]));    relay_conn far_2_2377_1_b(.in(far_2_2377_0[1]), .out(far_2_2377_1[1]));
    assign layer_2[337] = far_2_2377_1[0] ^ far_2_2377_1[1]; 
    wire [1:0] far_2_2378_0;    relay_conn far_2_2378_0_a(.in(layer_1[424]), .out(far_2_2378_0[0]));    relay_conn far_2_2378_0_b(.in(layer_1[469]), .out(far_2_2378_0[1]));
    assign layer_2[338] = ~far_2_2378_0[0] | (far_2_2378_0[0] & far_2_2378_0[1]); 
    assign layer_2[339] = layer_1[16] | layer_1[4]; 
    wire [1:0] far_2_2380_0;    relay_conn far_2_2380_0_a(.in(layer_1[404]), .out(far_2_2380_0[0]));    relay_conn far_2_2380_0_b(.in(layer_1[444]), .out(far_2_2380_0[1]));
    assign layer_2[340] = ~far_2_2380_0[1] | (far_2_2380_0[0] & far_2_2380_0[1]); 
    wire [1:0] far_2_2381_0;    relay_conn far_2_2381_0_a(.in(layer_1[558]), .out(far_2_2381_0[0]));    relay_conn far_2_2381_0_b(.in(layer_1[674]), .out(far_2_2381_0[1]));
    wire [1:0] far_2_2381_1;    relay_conn far_2_2381_1_a(.in(far_2_2381_0[0]), .out(far_2_2381_1[0]));    relay_conn far_2_2381_1_b(.in(far_2_2381_0[1]), .out(far_2_2381_1[1]));
    wire [1:0] far_2_2381_2;    relay_conn far_2_2381_2_a(.in(far_2_2381_1[0]), .out(far_2_2381_2[0]));    relay_conn far_2_2381_2_b(.in(far_2_2381_1[1]), .out(far_2_2381_2[1]));
    assign layer_2[341] = far_2_2381_2[0] & far_2_2381_2[1]; 
    assign layer_2[342] = ~layer_1[248] | (layer_1[248] & layer_1[250]); 
    wire [1:0] far_2_2383_0;    relay_conn far_2_2383_0_a(.in(layer_1[577]), .out(far_2_2383_0[0]));    relay_conn far_2_2383_0_b(.in(layer_1[537]), .out(far_2_2383_0[1]));
    assign layer_2[343] = ~(far_2_2383_0[0] & far_2_2383_0[1]); 
    wire [1:0] far_2_2384_0;    relay_conn far_2_2384_0_a(.in(layer_1[45]), .out(far_2_2384_0[0]));    relay_conn far_2_2384_0_b(.in(layer_1[130]), .out(far_2_2384_0[1]));
    wire [1:0] far_2_2384_1;    relay_conn far_2_2384_1_a(.in(far_2_2384_0[0]), .out(far_2_2384_1[0]));    relay_conn far_2_2384_1_b(.in(far_2_2384_0[1]), .out(far_2_2384_1[1]));
    assign layer_2[344] = ~(far_2_2384_1[0] ^ far_2_2384_1[1]); 
    wire [1:0] far_2_2385_0;    relay_conn far_2_2385_0_a(.in(layer_1[768]), .out(far_2_2385_0[0]));    relay_conn far_2_2385_0_b(.in(layer_1[876]), .out(far_2_2385_0[1]));
    wire [1:0] far_2_2385_1;    relay_conn far_2_2385_1_a(.in(far_2_2385_0[0]), .out(far_2_2385_1[0]));    relay_conn far_2_2385_1_b(.in(far_2_2385_0[1]), .out(far_2_2385_1[1]));
    wire [1:0] far_2_2385_2;    relay_conn far_2_2385_2_a(.in(far_2_2385_1[0]), .out(far_2_2385_2[0]));    relay_conn far_2_2385_2_b(.in(far_2_2385_1[1]), .out(far_2_2385_2[1]));
    assign layer_2[345] = far_2_2385_2[1]; 
    wire [1:0] far_2_2386_0;    relay_conn far_2_2386_0_a(.in(layer_1[432]), .out(far_2_2386_0[0]));    relay_conn far_2_2386_0_b(.in(layer_1[558]), .out(far_2_2386_0[1]));
    wire [1:0] far_2_2386_1;    relay_conn far_2_2386_1_a(.in(far_2_2386_0[0]), .out(far_2_2386_1[0]));    relay_conn far_2_2386_1_b(.in(far_2_2386_0[1]), .out(far_2_2386_1[1]));
    wire [1:0] far_2_2386_2;    relay_conn far_2_2386_2_a(.in(far_2_2386_1[0]), .out(far_2_2386_2[0]));    relay_conn far_2_2386_2_b(.in(far_2_2386_1[1]), .out(far_2_2386_2[1]));
    assign layer_2[346] = far_2_2386_2[0] & far_2_2386_2[1]; 
    assign layer_2[347] = layer_1[50]; 
    wire [1:0] far_2_2388_0;    relay_conn far_2_2388_0_a(.in(layer_1[894]), .out(far_2_2388_0[0]));    relay_conn far_2_2388_0_b(.in(layer_1[962]), .out(far_2_2388_0[1]));
    wire [1:0] far_2_2388_1;    relay_conn far_2_2388_1_a(.in(far_2_2388_0[0]), .out(far_2_2388_1[0]));    relay_conn far_2_2388_1_b(.in(far_2_2388_0[1]), .out(far_2_2388_1[1]));
    assign layer_2[348] = ~far_2_2388_1[1] | (far_2_2388_1[0] & far_2_2388_1[1]); 
    wire [1:0] far_2_2389_0;    relay_conn far_2_2389_0_a(.in(layer_1[88]), .out(far_2_2389_0[0]));    relay_conn far_2_2389_0_b(.in(layer_1[9]), .out(far_2_2389_0[1]));
    wire [1:0] far_2_2389_1;    relay_conn far_2_2389_1_a(.in(far_2_2389_0[0]), .out(far_2_2389_1[0]));    relay_conn far_2_2389_1_b(.in(far_2_2389_0[1]), .out(far_2_2389_1[1]));
    assign layer_2[349] = ~(far_2_2389_1[0] ^ far_2_2389_1[1]); 
    wire [1:0] far_2_2390_0;    relay_conn far_2_2390_0_a(.in(layer_1[347]), .out(far_2_2390_0[0]));    relay_conn far_2_2390_0_b(.in(layer_1[428]), .out(far_2_2390_0[1]));
    wire [1:0] far_2_2390_1;    relay_conn far_2_2390_1_a(.in(far_2_2390_0[0]), .out(far_2_2390_1[0]));    relay_conn far_2_2390_1_b(.in(far_2_2390_0[1]), .out(far_2_2390_1[1]));
    assign layer_2[350] = ~far_2_2390_1[1]; 
    wire [1:0] far_2_2391_0;    relay_conn far_2_2391_0_a(.in(layer_1[203]), .out(far_2_2391_0[0]));    relay_conn far_2_2391_0_b(.in(layer_1[162]), .out(far_2_2391_0[1]));
    assign layer_2[351] = ~(far_2_2391_0[0] | far_2_2391_0[1]); 
    wire [1:0] far_2_2392_0;    relay_conn far_2_2392_0_a(.in(layer_1[885]), .out(far_2_2392_0[0]));    relay_conn far_2_2392_0_b(.in(layer_1[935]), .out(far_2_2392_0[1]));
    assign layer_2[352] = far_2_2392_0[0] & ~far_2_2392_0[1]; 
    wire [1:0] far_2_2393_0;    relay_conn far_2_2393_0_a(.in(layer_1[0]), .out(far_2_2393_0[0]));    relay_conn far_2_2393_0_b(.in(layer_1[64]), .out(far_2_2393_0[1]));
    wire [1:0] far_2_2393_1;    relay_conn far_2_2393_1_a(.in(far_2_2393_0[0]), .out(far_2_2393_1[0]));    relay_conn far_2_2393_1_b(.in(far_2_2393_0[1]), .out(far_2_2393_1[1]));
    assign layer_2[353] = far_2_2393_1[0] ^ far_2_2393_1[1]; 
    wire [1:0] far_2_2394_0;    relay_conn far_2_2394_0_a(.in(layer_1[105]), .out(far_2_2394_0[0]));    relay_conn far_2_2394_0_b(.in(layer_1[28]), .out(far_2_2394_0[1]));
    wire [1:0] far_2_2394_1;    relay_conn far_2_2394_1_a(.in(far_2_2394_0[0]), .out(far_2_2394_1[0]));    relay_conn far_2_2394_1_b(.in(far_2_2394_0[1]), .out(far_2_2394_1[1]));
    assign layer_2[354] = ~far_2_2394_1[1] | (far_2_2394_1[0] & far_2_2394_1[1]); 
    wire [1:0] far_2_2395_0;    relay_conn far_2_2395_0_a(.in(layer_1[664]), .out(far_2_2395_0[0]));    relay_conn far_2_2395_0_b(.in(layer_1[732]), .out(far_2_2395_0[1]));
    wire [1:0] far_2_2395_1;    relay_conn far_2_2395_1_a(.in(far_2_2395_0[0]), .out(far_2_2395_1[0]));    relay_conn far_2_2395_1_b(.in(far_2_2395_0[1]), .out(far_2_2395_1[1]));
    assign layer_2[355] = ~(far_2_2395_1[0] & far_2_2395_1[1]); 
    wire [1:0] far_2_2396_0;    relay_conn far_2_2396_0_a(.in(layer_1[567]), .out(far_2_2396_0[0]));    relay_conn far_2_2396_0_b(.in(layer_1[617]), .out(far_2_2396_0[1]));
    assign layer_2[356] = ~(far_2_2396_0[0] & far_2_2396_0[1]); 
    wire [1:0] far_2_2397_0;    relay_conn far_2_2397_0_a(.in(layer_1[795]), .out(far_2_2397_0[0]));    relay_conn far_2_2397_0_b(.in(layer_1[676]), .out(far_2_2397_0[1]));
    wire [1:0] far_2_2397_1;    relay_conn far_2_2397_1_a(.in(far_2_2397_0[0]), .out(far_2_2397_1[0]));    relay_conn far_2_2397_1_b(.in(far_2_2397_0[1]), .out(far_2_2397_1[1]));
    wire [1:0] far_2_2397_2;    relay_conn far_2_2397_2_a(.in(far_2_2397_1[0]), .out(far_2_2397_2[0]));    relay_conn far_2_2397_2_b(.in(far_2_2397_1[1]), .out(far_2_2397_2[1]));
    assign layer_2[357] = ~far_2_2397_2[1] | (far_2_2397_2[0] & far_2_2397_2[1]); 
    wire [1:0] far_2_2398_0;    relay_conn far_2_2398_0_a(.in(layer_1[901]), .out(far_2_2398_0[0]));    relay_conn far_2_2398_0_b(.in(layer_1[807]), .out(far_2_2398_0[1]));
    wire [1:0] far_2_2398_1;    relay_conn far_2_2398_1_a(.in(far_2_2398_0[0]), .out(far_2_2398_1[0]));    relay_conn far_2_2398_1_b(.in(far_2_2398_0[1]), .out(far_2_2398_1[1]));
    assign layer_2[358] = ~(far_2_2398_1[0] | far_2_2398_1[1]); 
    wire [1:0] far_2_2399_0;    relay_conn far_2_2399_0_a(.in(layer_1[159]), .out(far_2_2399_0[0]));    relay_conn far_2_2399_0_b(.in(layer_1[248]), .out(far_2_2399_0[1]));
    wire [1:0] far_2_2399_1;    relay_conn far_2_2399_1_a(.in(far_2_2399_0[0]), .out(far_2_2399_1[0]));    relay_conn far_2_2399_1_b(.in(far_2_2399_0[1]), .out(far_2_2399_1[1]));
    assign layer_2[359] = ~(far_2_2399_1[0] & far_2_2399_1[1]); 
    wire [1:0] far_2_2400_0;    relay_conn far_2_2400_0_a(.in(layer_1[184]), .out(far_2_2400_0[0]));    relay_conn far_2_2400_0_b(.in(layer_1[246]), .out(far_2_2400_0[1]));
    assign layer_2[360] = ~far_2_2400_0[1] | (far_2_2400_0[0] & far_2_2400_0[1]); 
    wire [1:0] far_2_2401_0;    relay_conn far_2_2401_0_a(.in(layer_1[615]), .out(far_2_2401_0[0]));    relay_conn far_2_2401_0_b(.in(layer_1[514]), .out(far_2_2401_0[1]));
    wire [1:0] far_2_2401_1;    relay_conn far_2_2401_1_a(.in(far_2_2401_0[0]), .out(far_2_2401_1[0]));    relay_conn far_2_2401_1_b(.in(far_2_2401_0[1]), .out(far_2_2401_1[1]));
    wire [1:0] far_2_2401_2;    relay_conn far_2_2401_2_a(.in(far_2_2401_1[0]), .out(far_2_2401_2[0]));    relay_conn far_2_2401_2_b(.in(far_2_2401_1[1]), .out(far_2_2401_2[1]));
    assign layer_2[361] = ~(far_2_2401_2[0] | far_2_2401_2[1]); 
    wire [1:0] far_2_2402_0;    relay_conn far_2_2402_0_a(.in(layer_1[180]), .out(far_2_2402_0[0]));    relay_conn far_2_2402_0_b(.in(layer_1[213]), .out(far_2_2402_0[1]));
    assign layer_2[362] = ~far_2_2402_0[1] | (far_2_2402_0[0] & far_2_2402_0[1]); 
    wire [1:0] far_2_2403_0;    relay_conn far_2_2403_0_a(.in(layer_1[442]), .out(far_2_2403_0[0]));    relay_conn far_2_2403_0_b(.in(layer_1[559]), .out(far_2_2403_0[1]));
    wire [1:0] far_2_2403_1;    relay_conn far_2_2403_1_a(.in(far_2_2403_0[0]), .out(far_2_2403_1[0]));    relay_conn far_2_2403_1_b(.in(far_2_2403_0[1]), .out(far_2_2403_1[1]));
    wire [1:0] far_2_2403_2;    relay_conn far_2_2403_2_a(.in(far_2_2403_1[0]), .out(far_2_2403_2[0]));    relay_conn far_2_2403_2_b(.in(far_2_2403_1[1]), .out(far_2_2403_2[1]));
    assign layer_2[363] = far_2_2403_2[0] ^ far_2_2403_2[1]; 
    wire [1:0] far_2_2404_0;    relay_conn far_2_2404_0_a(.in(layer_1[184]), .out(far_2_2404_0[0]));    relay_conn far_2_2404_0_b(.in(layer_1[261]), .out(far_2_2404_0[1]));
    wire [1:0] far_2_2404_1;    relay_conn far_2_2404_1_a(.in(far_2_2404_0[0]), .out(far_2_2404_1[0]));    relay_conn far_2_2404_1_b(.in(far_2_2404_0[1]), .out(far_2_2404_1[1]));
    assign layer_2[364] = far_2_2404_1[0] & ~far_2_2404_1[1]; 
    wire [1:0] far_2_2405_0;    relay_conn far_2_2405_0_a(.in(layer_1[796]), .out(far_2_2405_0[0]));    relay_conn far_2_2405_0_b(.in(layer_1[742]), .out(far_2_2405_0[1]));
    assign layer_2[365] = far_2_2405_0[1] & ~far_2_2405_0[0]; 
    wire [1:0] far_2_2406_0;    relay_conn far_2_2406_0_a(.in(layer_1[605]), .out(far_2_2406_0[0]));    relay_conn far_2_2406_0_b(.in(layer_1[477]), .out(far_2_2406_0[1]));
    wire [1:0] far_2_2406_1;    relay_conn far_2_2406_1_a(.in(far_2_2406_0[0]), .out(far_2_2406_1[0]));    relay_conn far_2_2406_1_b(.in(far_2_2406_0[1]), .out(far_2_2406_1[1]));
    wire [1:0] far_2_2406_2;    relay_conn far_2_2406_2_a(.in(far_2_2406_1[0]), .out(far_2_2406_2[0]));    relay_conn far_2_2406_2_b(.in(far_2_2406_1[1]), .out(far_2_2406_2[1]));
    wire [1:0] far_2_2406_3;    relay_conn far_2_2406_3_a(.in(far_2_2406_2[0]), .out(far_2_2406_3[0]));    relay_conn far_2_2406_3_b(.in(far_2_2406_2[1]), .out(far_2_2406_3[1]));
    assign layer_2[366] = far_2_2406_3[0] & far_2_2406_3[1]; 
    assign layer_2[367] = ~(layer_1[55] | layer_1[66]); 
    wire [1:0] far_2_2408_0;    relay_conn far_2_2408_0_a(.in(layer_1[212]), .out(far_2_2408_0[0]));    relay_conn far_2_2408_0_b(.in(layer_1[248]), .out(far_2_2408_0[1]));
    assign layer_2[368] = ~far_2_2408_0[1] | (far_2_2408_0[0] & far_2_2408_0[1]); 
    assign layer_2[369] = ~(layer_1[109] | layer_1[99]); 
    wire [1:0] far_2_2410_0;    relay_conn far_2_2410_0_a(.in(layer_1[326]), .out(far_2_2410_0[0]));    relay_conn far_2_2410_0_b(.in(layer_1[294]), .out(far_2_2410_0[1]));
    assign layer_2[370] = far_2_2410_0[1]; 
    wire [1:0] far_2_2411_0;    relay_conn far_2_2411_0_a(.in(layer_1[898]), .out(far_2_2411_0[0]));    relay_conn far_2_2411_0_b(.in(layer_1[965]), .out(far_2_2411_0[1]));
    wire [1:0] far_2_2411_1;    relay_conn far_2_2411_1_a(.in(far_2_2411_0[0]), .out(far_2_2411_1[0]));    relay_conn far_2_2411_1_b(.in(far_2_2411_0[1]), .out(far_2_2411_1[1]));
    assign layer_2[371] = far_2_2411_1[1]; 
    assign layer_2[372] = layer_1[928] ^ layer_1[955]; 
    wire [1:0] far_2_2413_0;    relay_conn far_2_2413_0_a(.in(layer_1[557]), .out(far_2_2413_0[0]));    relay_conn far_2_2413_0_b(.in(layer_1[662]), .out(far_2_2413_0[1]));
    wire [1:0] far_2_2413_1;    relay_conn far_2_2413_1_a(.in(far_2_2413_0[0]), .out(far_2_2413_1[0]));    relay_conn far_2_2413_1_b(.in(far_2_2413_0[1]), .out(far_2_2413_1[1]));
    wire [1:0] far_2_2413_2;    relay_conn far_2_2413_2_a(.in(far_2_2413_1[0]), .out(far_2_2413_2[0]));    relay_conn far_2_2413_2_b(.in(far_2_2413_1[1]), .out(far_2_2413_2[1]));
    assign layer_2[373] = far_2_2413_2[0]; 
    assign layer_2[374] = layer_1[373] & ~layer_1[390]; 
    assign layer_2[375] = ~(layer_1[63] & layer_1[40]); 
    wire [1:0] far_2_2416_0;    relay_conn far_2_2416_0_a(.in(layer_1[390]), .out(far_2_2416_0[0]));    relay_conn far_2_2416_0_b(.in(layer_1[440]), .out(far_2_2416_0[1]));
    assign layer_2[376] = far_2_2416_0[1]; 
    wire [1:0] far_2_2417_0;    relay_conn far_2_2417_0_a(.in(layer_1[422]), .out(far_2_2417_0[0]));    relay_conn far_2_2417_0_b(.in(layer_1[524]), .out(far_2_2417_0[1]));
    wire [1:0] far_2_2417_1;    relay_conn far_2_2417_1_a(.in(far_2_2417_0[0]), .out(far_2_2417_1[0]));    relay_conn far_2_2417_1_b(.in(far_2_2417_0[1]), .out(far_2_2417_1[1]));
    wire [1:0] far_2_2417_2;    relay_conn far_2_2417_2_a(.in(far_2_2417_1[0]), .out(far_2_2417_2[0]));    relay_conn far_2_2417_2_b(.in(far_2_2417_1[1]), .out(far_2_2417_2[1]));
    assign layer_2[377] = far_2_2417_2[1] & ~far_2_2417_2[0]; 
    wire [1:0] far_2_2418_0;    relay_conn far_2_2418_0_a(.in(layer_1[40]), .out(far_2_2418_0[0]));    relay_conn far_2_2418_0_b(.in(layer_1[156]), .out(far_2_2418_0[1]));
    wire [1:0] far_2_2418_1;    relay_conn far_2_2418_1_a(.in(far_2_2418_0[0]), .out(far_2_2418_1[0]));    relay_conn far_2_2418_1_b(.in(far_2_2418_0[1]), .out(far_2_2418_1[1]));
    wire [1:0] far_2_2418_2;    relay_conn far_2_2418_2_a(.in(far_2_2418_1[0]), .out(far_2_2418_2[0]));    relay_conn far_2_2418_2_b(.in(far_2_2418_1[1]), .out(far_2_2418_2[1]));
    assign layer_2[378] = ~far_2_2418_2[0]; 
    wire [1:0] far_2_2419_0;    relay_conn far_2_2419_0_a(.in(layer_1[333]), .out(far_2_2419_0[0]));    relay_conn far_2_2419_0_b(.in(layer_1[222]), .out(far_2_2419_0[1]));
    wire [1:0] far_2_2419_1;    relay_conn far_2_2419_1_a(.in(far_2_2419_0[0]), .out(far_2_2419_1[0]));    relay_conn far_2_2419_1_b(.in(far_2_2419_0[1]), .out(far_2_2419_1[1]));
    wire [1:0] far_2_2419_2;    relay_conn far_2_2419_2_a(.in(far_2_2419_1[0]), .out(far_2_2419_2[0]));    relay_conn far_2_2419_2_b(.in(far_2_2419_1[1]), .out(far_2_2419_2[1]));
    assign layer_2[379] = far_2_2419_2[1]; 
    wire [1:0] far_2_2420_0;    relay_conn far_2_2420_0_a(.in(layer_1[533]), .out(far_2_2420_0[0]));    relay_conn far_2_2420_0_b(.in(layer_1[626]), .out(far_2_2420_0[1]));
    wire [1:0] far_2_2420_1;    relay_conn far_2_2420_1_a(.in(far_2_2420_0[0]), .out(far_2_2420_1[0]));    relay_conn far_2_2420_1_b(.in(far_2_2420_0[1]), .out(far_2_2420_1[1]));
    assign layer_2[380] = far_2_2420_1[0] & far_2_2420_1[1]; 
    assign layer_2[381] = layer_1[471] & ~layer_1[442]; 
    wire [1:0] far_2_2422_0;    relay_conn far_2_2422_0_a(.in(layer_1[361]), .out(far_2_2422_0[0]));    relay_conn far_2_2422_0_b(.in(layer_1[400]), .out(far_2_2422_0[1]));
    assign layer_2[382] = ~(far_2_2422_0[0] & far_2_2422_0[1]); 
    assign layer_2[383] = layer_1[437]; 
    wire [1:0] far_2_2424_0;    relay_conn far_2_2424_0_a(.in(layer_1[846]), .out(far_2_2424_0[0]));    relay_conn far_2_2424_0_b(.in(layer_1[910]), .out(far_2_2424_0[1]));
    wire [1:0] far_2_2424_1;    relay_conn far_2_2424_1_a(.in(far_2_2424_0[0]), .out(far_2_2424_1[0]));    relay_conn far_2_2424_1_b(.in(far_2_2424_0[1]), .out(far_2_2424_1[1]));
    assign layer_2[384] = far_2_2424_1[0] | far_2_2424_1[1]; 
    wire [1:0] far_2_2425_0;    relay_conn far_2_2425_0_a(.in(layer_1[202]), .out(far_2_2425_0[0]));    relay_conn far_2_2425_0_b(.in(layer_1[155]), .out(far_2_2425_0[1]));
    assign layer_2[385] = far_2_2425_0[0] & far_2_2425_0[1]; 
    assign layer_2[386] = ~layer_1[558]; 
    wire [1:0] far_2_2427_0;    relay_conn far_2_2427_0_a(.in(layer_1[144]), .out(far_2_2427_0[0]));    relay_conn far_2_2427_0_b(.in(layer_1[217]), .out(far_2_2427_0[1]));
    wire [1:0] far_2_2427_1;    relay_conn far_2_2427_1_a(.in(far_2_2427_0[0]), .out(far_2_2427_1[0]));    relay_conn far_2_2427_1_b(.in(far_2_2427_0[1]), .out(far_2_2427_1[1]));
    assign layer_2[387] = ~far_2_2427_1[1] | (far_2_2427_1[0] & far_2_2427_1[1]); 
    wire [1:0] far_2_2428_0;    relay_conn far_2_2428_0_a(.in(layer_1[153]), .out(far_2_2428_0[0]));    relay_conn far_2_2428_0_b(.in(layer_1[74]), .out(far_2_2428_0[1]));
    wire [1:0] far_2_2428_1;    relay_conn far_2_2428_1_a(.in(far_2_2428_0[0]), .out(far_2_2428_1[0]));    relay_conn far_2_2428_1_b(.in(far_2_2428_0[1]), .out(far_2_2428_1[1]));
    assign layer_2[388] = ~(far_2_2428_1[0] | far_2_2428_1[1]); 
    wire [1:0] far_2_2429_0;    relay_conn far_2_2429_0_a(.in(layer_1[169]), .out(far_2_2429_0[0]));    relay_conn far_2_2429_0_b(.in(layer_1[223]), .out(far_2_2429_0[1]));
    assign layer_2[389] = ~far_2_2429_0[0]; 
    wire [1:0] far_2_2430_0;    relay_conn far_2_2430_0_a(.in(layer_1[71]), .out(far_2_2430_0[0]));    relay_conn far_2_2430_0_b(.in(layer_1[25]), .out(far_2_2430_0[1]));
    assign layer_2[390] = far_2_2430_0[0] & far_2_2430_0[1]; 
    assign layer_2[391] = layer_1[177] & ~layer_1[202]; 
    wire [1:0] far_2_2432_0;    relay_conn far_2_2432_0_a(.in(layer_1[482]), .out(far_2_2432_0[0]));    relay_conn far_2_2432_0_b(.in(layer_1[557]), .out(far_2_2432_0[1]));
    wire [1:0] far_2_2432_1;    relay_conn far_2_2432_1_a(.in(far_2_2432_0[0]), .out(far_2_2432_1[0]));    relay_conn far_2_2432_1_b(.in(far_2_2432_0[1]), .out(far_2_2432_1[1]));
    assign layer_2[392] = ~(far_2_2432_1[0] | far_2_2432_1[1]); 
    wire [1:0] far_2_2433_0;    relay_conn far_2_2433_0_a(.in(layer_1[296]), .out(far_2_2433_0[0]));    relay_conn far_2_2433_0_b(.in(layer_1[202]), .out(far_2_2433_0[1]));
    wire [1:0] far_2_2433_1;    relay_conn far_2_2433_1_a(.in(far_2_2433_0[0]), .out(far_2_2433_1[0]));    relay_conn far_2_2433_1_b(.in(far_2_2433_0[1]), .out(far_2_2433_1[1]));
    assign layer_2[393] = ~far_2_2433_1[1] | (far_2_2433_1[0] & far_2_2433_1[1]); 
    wire [1:0] far_2_2434_0;    relay_conn far_2_2434_0_a(.in(layer_1[298]), .out(far_2_2434_0[0]));    relay_conn far_2_2434_0_b(.in(layer_1[368]), .out(far_2_2434_0[1]));
    wire [1:0] far_2_2434_1;    relay_conn far_2_2434_1_a(.in(far_2_2434_0[0]), .out(far_2_2434_1[0]));    relay_conn far_2_2434_1_b(.in(far_2_2434_0[1]), .out(far_2_2434_1[1]));
    assign layer_2[394] = ~far_2_2434_1[1] | (far_2_2434_1[0] & far_2_2434_1[1]); 
    wire [1:0] far_2_2435_0;    relay_conn far_2_2435_0_a(.in(layer_1[288]), .out(far_2_2435_0[0]));    relay_conn far_2_2435_0_b(.in(layer_1[327]), .out(far_2_2435_0[1]));
    assign layer_2[395] = ~far_2_2435_0[0]; 
    wire [1:0] far_2_2436_0;    relay_conn far_2_2436_0_a(.in(layer_1[177]), .out(far_2_2436_0[0]));    relay_conn far_2_2436_0_b(.in(layer_1[287]), .out(far_2_2436_0[1]));
    wire [1:0] far_2_2436_1;    relay_conn far_2_2436_1_a(.in(far_2_2436_0[0]), .out(far_2_2436_1[0]));    relay_conn far_2_2436_1_b(.in(far_2_2436_0[1]), .out(far_2_2436_1[1]));
    wire [1:0] far_2_2436_2;    relay_conn far_2_2436_2_a(.in(far_2_2436_1[0]), .out(far_2_2436_2[0]));    relay_conn far_2_2436_2_b(.in(far_2_2436_1[1]), .out(far_2_2436_2[1]));
    assign layer_2[396] = far_2_2436_2[1] & ~far_2_2436_2[0]; 
    wire [1:0] far_2_2437_0;    relay_conn far_2_2437_0_a(.in(layer_1[251]), .out(far_2_2437_0[0]));    relay_conn far_2_2437_0_b(.in(layer_1[190]), .out(far_2_2437_0[1]));
    assign layer_2[397] = far_2_2437_0[0] | far_2_2437_0[1]; 
    wire [1:0] far_2_2438_0;    relay_conn far_2_2438_0_a(.in(layer_1[801]), .out(far_2_2438_0[0]));    relay_conn far_2_2438_0_b(.in(layer_1[917]), .out(far_2_2438_0[1]));
    wire [1:0] far_2_2438_1;    relay_conn far_2_2438_1_a(.in(far_2_2438_0[0]), .out(far_2_2438_1[0]));    relay_conn far_2_2438_1_b(.in(far_2_2438_0[1]), .out(far_2_2438_1[1]));
    wire [1:0] far_2_2438_2;    relay_conn far_2_2438_2_a(.in(far_2_2438_1[0]), .out(far_2_2438_2[0]));    relay_conn far_2_2438_2_b(.in(far_2_2438_1[1]), .out(far_2_2438_2[1]));
    assign layer_2[398] = far_2_2438_2[0] | far_2_2438_2[1]; 
    wire [1:0] far_2_2439_0;    relay_conn far_2_2439_0_a(.in(layer_1[707]), .out(far_2_2439_0[0]));    relay_conn far_2_2439_0_b(.in(layer_1[835]), .out(far_2_2439_0[1]));
    wire [1:0] far_2_2439_1;    relay_conn far_2_2439_1_a(.in(far_2_2439_0[0]), .out(far_2_2439_1[0]));    relay_conn far_2_2439_1_b(.in(far_2_2439_0[1]), .out(far_2_2439_1[1]));
    wire [1:0] far_2_2439_2;    relay_conn far_2_2439_2_a(.in(far_2_2439_1[0]), .out(far_2_2439_2[0]));    relay_conn far_2_2439_2_b(.in(far_2_2439_1[1]), .out(far_2_2439_2[1]));
    wire [1:0] far_2_2439_3;    relay_conn far_2_2439_3_a(.in(far_2_2439_2[0]), .out(far_2_2439_3[0]));    relay_conn far_2_2439_3_b(.in(far_2_2439_2[1]), .out(far_2_2439_3[1]));
    assign layer_2[399] = far_2_2439_3[0] | far_2_2439_3[1]; 
    assign layer_2[400] = ~(layer_1[64] ^ layer_1[38]); 
    wire [1:0] far_2_2441_0;    relay_conn far_2_2441_0_a(.in(layer_1[241]), .out(far_2_2441_0[0]));    relay_conn far_2_2441_0_b(.in(layer_1[317]), .out(far_2_2441_0[1]));
    wire [1:0] far_2_2441_1;    relay_conn far_2_2441_1_a(.in(far_2_2441_0[0]), .out(far_2_2441_1[0]));    relay_conn far_2_2441_1_b(.in(far_2_2441_0[1]), .out(far_2_2441_1[1]));
    assign layer_2[401] = ~(far_2_2441_1[0] | far_2_2441_1[1]); 
    wire [1:0] far_2_2442_0;    relay_conn far_2_2442_0_a(.in(layer_1[204]), .out(far_2_2442_0[0]));    relay_conn far_2_2442_0_b(.in(layer_1[99]), .out(far_2_2442_0[1]));
    wire [1:0] far_2_2442_1;    relay_conn far_2_2442_1_a(.in(far_2_2442_0[0]), .out(far_2_2442_1[0]));    relay_conn far_2_2442_1_b(.in(far_2_2442_0[1]), .out(far_2_2442_1[1]));
    wire [1:0] far_2_2442_2;    relay_conn far_2_2442_2_a(.in(far_2_2442_1[0]), .out(far_2_2442_2[0]));    relay_conn far_2_2442_2_b(.in(far_2_2442_1[1]), .out(far_2_2442_2[1]));
    assign layer_2[402] = ~(far_2_2442_2[0] ^ far_2_2442_2[1]); 
    wire [1:0] far_2_2443_0;    relay_conn far_2_2443_0_a(.in(layer_1[663]), .out(far_2_2443_0[0]));    relay_conn far_2_2443_0_b(.in(layer_1[750]), .out(far_2_2443_0[1]));
    wire [1:0] far_2_2443_1;    relay_conn far_2_2443_1_a(.in(far_2_2443_0[0]), .out(far_2_2443_1[0]));    relay_conn far_2_2443_1_b(.in(far_2_2443_0[1]), .out(far_2_2443_1[1]));
    assign layer_2[403] = far_2_2443_1[0] & ~far_2_2443_1[1]; 
    wire [1:0] far_2_2444_0;    relay_conn far_2_2444_0_a(.in(layer_1[393]), .out(far_2_2444_0[0]));    relay_conn far_2_2444_0_b(.in(layer_1[467]), .out(far_2_2444_0[1]));
    wire [1:0] far_2_2444_1;    relay_conn far_2_2444_1_a(.in(far_2_2444_0[0]), .out(far_2_2444_1[0]));    relay_conn far_2_2444_1_b(.in(far_2_2444_0[1]), .out(far_2_2444_1[1]));
    assign layer_2[404] = far_2_2444_1[0]; 
    wire [1:0] far_2_2445_0;    relay_conn far_2_2445_0_a(.in(layer_1[929]), .out(far_2_2445_0[0]));    relay_conn far_2_2445_0_b(.in(layer_1[987]), .out(far_2_2445_0[1]));
    assign layer_2[405] = far_2_2445_0[0] | far_2_2445_0[1]; 
    wire [1:0] far_2_2446_0;    relay_conn far_2_2446_0_a(.in(layer_1[787]), .out(far_2_2446_0[0]));    relay_conn far_2_2446_0_b(.in(layer_1[884]), .out(far_2_2446_0[1]));
    wire [1:0] far_2_2446_1;    relay_conn far_2_2446_1_a(.in(far_2_2446_0[0]), .out(far_2_2446_1[0]));    relay_conn far_2_2446_1_b(.in(far_2_2446_0[1]), .out(far_2_2446_1[1]));
    wire [1:0] far_2_2446_2;    relay_conn far_2_2446_2_a(.in(far_2_2446_1[0]), .out(far_2_2446_2[0]));    relay_conn far_2_2446_2_b(.in(far_2_2446_1[1]), .out(far_2_2446_2[1]));
    assign layer_2[406] = ~(far_2_2446_2[0] | far_2_2446_2[1]); 
    assign layer_2[407] = ~(layer_1[50] | layer_1[57]); 
    assign layer_2[408] = layer_1[41] & ~layer_1[33]; 
    assign layer_2[409] = layer_1[1] & ~layer_1[21]; 
    wire [1:0] far_2_2450_0;    relay_conn far_2_2450_0_a(.in(layer_1[11]), .out(far_2_2450_0[0]));    relay_conn far_2_2450_0_b(.in(layer_1[87]), .out(far_2_2450_0[1]));
    wire [1:0] far_2_2450_1;    relay_conn far_2_2450_1_a(.in(far_2_2450_0[0]), .out(far_2_2450_1[0]));    relay_conn far_2_2450_1_b(.in(far_2_2450_0[1]), .out(far_2_2450_1[1]));
    assign layer_2[410] = ~(far_2_2450_1[0] | far_2_2450_1[1]); 
    wire [1:0] far_2_2451_0;    relay_conn far_2_2451_0_a(.in(layer_1[338]), .out(far_2_2451_0[0]));    relay_conn far_2_2451_0_b(.in(layer_1[455]), .out(far_2_2451_0[1]));
    wire [1:0] far_2_2451_1;    relay_conn far_2_2451_1_a(.in(far_2_2451_0[0]), .out(far_2_2451_1[0]));    relay_conn far_2_2451_1_b(.in(far_2_2451_0[1]), .out(far_2_2451_1[1]));
    wire [1:0] far_2_2451_2;    relay_conn far_2_2451_2_a(.in(far_2_2451_1[0]), .out(far_2_2451_2[0]));    relay_conn far_2_2451_2_b(.in(far_2_2451_1[1]), .out(far_2_2451_2[1]));
    assign layer_2[411] = ~(far_2_2451_2[0] ^ far_2_2451_2[1]); 
    wire [1:0] far_2_2452_0;    relay_conn far_2_2452_0_a(.in(layer_1[221]), .out(far_2_2452_0[0]));    relay_conn far_2_2452_0_b(.in(layer_1[296]), .out(far_2_2452_0[1]));
    wire [1:0] far_2_2452_1;    relay_conn far_2_2452_1_a(.in(far_2_2452_0[0]), .out(far_2_2452_1[0]));    relay_conn far_2_2452_1_b(.in(far_2_2452_0[1]), .out(far_2_2452_1[1]));
    assign layer_2[412] = ~far_2_2452_1[1] | (far_2_2452_1[0] & far_2_2452_1[1]); 
    wire [1:0] far_2_2453_0;    relay_conn far_2_2453_0_a(.in(layer_1[1006]), .out(far_2_2453_0[0]));    relay_conn far_2_2453_0_b(.in(layer_1[917]), .out(far_2_2453_0[1]));
    wire [1:0] far_2_2453_1;    relay_conn far_2_2453_1_a(.in(far_2_2453_0[0]), .out(far_2_2453_1[0]));    relay_conn far_2_2453_1_b(.in(far_2_2453_0[1]), .out(far_2_2453_1[1]));
    assign layer_2[413] = far_2_2453_1[1]; 
    assign layer_2[414] = ~layer_1[439]; 
    wire [1:0] far_2_2455_0;    relay_conn far_2_2455_0_a(.in(layer_1[583]), .out(far_2_2455_0[0]));    relay_conn far_2_2455_0_b(.in(layer_1[645]), .out(far_2_2455_0[1]));
    assign layer_2[415] = far_2_2455_0[1]; 
    wire [1:0] far_2_2456_0;    relay_conn far_2_2456_0_a(.in(layer_1[854]), .out(far_2_2456_0[0]));    relay_conn far_2_2456_0_b(.in(layer_1[900]), .out(far_2_2456_0[1]));
    assign layer_2[416] = far_2_2456_0[0]; 
    assign layer_2[417] = ~layer_1[184]; 
    assign layer_2[418] = layer_1[692]; 
    wire [1:0] far_2_2459_0;    relay_conn far_2_2459_0_a(.in(layer_1[352]), .out(far_2_2459_0[0]));    relay_conn far_2_2459_0_b(.in(layer_1[435]), .out(far_2_2459_0[1]));
    wire [1:0] far_2_2459_1;    relay_conn far_2_2459_1_a(.in(far_2_2459_0[0]), .out(far_2_2459_1[0]));    relay_conn far_2_2459_1_b(.in(far_2_2459_0[1]), .out(far_2_2459_1[1]));
    assign layer_2[419] = far_2_2459_1[0]; 
    wire [1:0] far_2_2460_0;    relay_conn far_2_2460_0_a(.in(layer_1[110]), .out(far_2_2460_0[0]));    relay_conn far_2_2460_0_b(.in(layer_1[201]), .out(far_2_2460_0[1]));
    wire [1:0] far_2_2460_1;    relay_conn far_2_2460_1_a(.in(far_2_2460_0[0]), .out(far_2_2460_1[0]));    relay_conn far_2_2460_1_b(.in(far_2_2460_0[1]), .out(far_2_2460_1[1]));
    assign layer_2[420] = far_2_2460_1[1]; 
    wire [1:0] far_2_2461_0;    relay_conn far_2_2461_0_a(.in(layer_1[768]), .out(far_2_2461_0[0]));    relay_conn far_2_2461_0_b(.in(layer_1[676]), .out(far_2_2461_0[1]));
    wire [1:0] far_2_2461_1;    relay_conn far_2_2461_1_a(.in(far_2_2461_0[0]), .out(far_2_2461_1[0]));    relay_conn far_2_2461_1_b(.in(far_2_2461_0[1]), .out(far_2_2461_1[1]));
    assign layer_2[421] = far_2_2461_1[0]; 
    wire [1:0] far_2_2462_0;    relay_conn far_2_2462_0_a(.in(layer_1[162]), .out(far_2_2462_0[0]));    relay_conn far_2_2462_0_b(.in(layer_1[212]), .out(far_2_2462_0[1]));
    assign layer_2[422] = far_2_2462_0[1]; 
    wire [1:0] far_2_2463_0;    relay_conn far_2_2463_0_a(.in(layer_1[984]), .out(far_2_2463_0[0]));    relay_conn far_2_2463_0_b(.in(layer_1[885]), .out(far_2_2463_0[1]));
    wire [1:0] far_2_2463_1;    relay_conn far_2_2463_1_a(.in(far_2_2463_0[0]), .out(far_2_2463_1[0]));    relay_conn far_2_2463_1_b(.in(far_2_2463_0[1]), .out(far_2_2463_1[1]));
    wire [1:0] far_2_2463_2;    relay_conn far_2_2463_2_a(.in(far_2_2463_1[0]), .out(far_2_2463_2[0]));    relay_conn far_2_2463_2_b(.in(far_2_2463_1[1]), .out(far_2_2463_2[1]));
    assign layer_2[423] = far_2_2463_2[0] | far_2_2463_2[1]; 
    wire [1:0] far_2_2464_0;    relay_conn far_2_2464_0_a(.in(layer_1[980]), .out(far_2_2464_0[0]));    relay_conn far_2_2464_0_b(.in(layer_1[928]), .out(far_2_2464_0[1]));
    assign layer_2[424] = ~far_2_2464_0[1]; 
    wire [1:0] far_2_2465_0;    relay_conn far_2_2465_0_a(.in(layer_1[9]), .out(far_2_2465_0[0]));    relay_conn far_2_2465_0_b(.in(layer_1[81]), .out(far_2_2465_0[1]));
    wire [1:0] far_2_2465_1;    relay_conn far_2_2465_1_a(.in(far_2_2465_0[0]), .out(far_2_2465_1[0]));    relay_conn far_2_2465_1_b(.in(far_2_2465_0[1]), .out(far_2_2465_1[1]));
    assign layer_2[425] = ~far_2_2465_1[1]; 
    wire [1:0] far_2_2466_0;    relay_conn far_2_2466_0_a(.in(layer_1[746]), .out(far_2_2466_0[0]));    relay_conn far_2_2466_0_b(.in(layer_1[833]), .out(far_2_2466_0[1]));
    wire [1:0] far_2_2466_1;    relay_conn far_2_2466_1_a(.in(far_2_2466_0[0]), .out(far_2_2466_1[0]));    relay_conn far_2_2466_1_b(.in(far_2_2466_0[1]), .out(far_2_2466_1[1]));
    assign layer_2[426] = ~far_2_2466_1[0] | (far_2_2466_1[0] & far_2_2466_1[1]); 
    wire [1:0] far_2_2467_0;    relay_conn far_2_2467_0_a(.in(layer_1[805]), .out(far_2_2467_0[0]));    relay_conn far_2_2467_0_b(.in(layer_1[903]), .out(far_2_2467_0[1]));
    wire [1:0] far_2_2467_1;    relay_conn far_2_2467_1_a(.in(far_2_2467_0[0]), .out(far_2_2467_1[0]));    relay_conn far_2_2467_1_b(.in(far_2_2467_0[1]), .out(far_2_2467_1[1]));
    wire [1:0] far_2_2467_2;    relay_conn far_2_2467_2_a(.in(far_2_2467_1[0]), .out(far_2_2467_2[0]));    relay_conn far_2_2467_2_b(.in(far_2_2467_1[1]), .out(far_2_2467_2[1]));
    assign layer_2[427] = ~far_2_2467_2[1]; 
    assign layer_2[428] = ~(layer_1[31] | layer_1[12]); 
    wire [1:0] far_2_2469_0;    relay_conn far_2_2469_0_a(.in(layer_1[265]), .out(far_2_2469_0[0]));    relay_conn far_2_2469_0_b(.in(layer_1[350]), .out(far_2_2469_0[1]));
    wire [1:0] far_2_2469_1;    relay_conn far_2_2469_1_a(.in(far_2_2469_0[0]), .out(far_2_2469_1[0]));    relay_conn far_2_2469_1_b(.in(far_2_2469_0[1]), .out(far_2_2469_1[1]));
    assign layer_2[429] = ~far_2_2469_1[1] | (far_2_2469_1[0] & far_2_2469_1[1]); 
    wire [1:0] far_2_2470_0;    relay_conn far_2_2470_0_a(.in(layer_1[578]), .out(far_2_2470_0[0]));    relay_conn far_2_2470_0_b(.in(layer_1[699]), .out(far_2_2470_0[1]));
    wire [1:0] far_2_2470_1;    relay_conn far_2_2470_1_a(.in(far_2_2470_0[0]), .out(far_2_2470_1[0]));    relay_conn far_2_2470_1_b(.in(far_2_2470_0[1]), .out(far_2_2470_1[1]));
    wire [1:0] far_2_2470_2;    relay_conn far_2_2470_2_a(.in(far_2_2470_1[0]), .out(far_2_2470_2[0]));    relay_conn far_2_2470_2_b(.in(far_2_2470_1[1]), .out(far_2_2470_2[1]));
    assign layer_2[430] = ~far_2_2470_2[0] | (far_2_2470_2[0] & far_2_2470_2[1]); 
    wire [1:0] far_2_2471_0;    relay_conn far_2_2471_0_a(.in(layer_1[164]), .out(far_2_2471_0[0]));    relay_conn far_2_2471_0_b(.in(layer_1[45]), .out(far_2_2471_0[1]));
    wire [1:0] far_2_2471_1;    relay_conn far_2_2471_1_a(.in(far_2_2471_0[0]), .out(far_2_2471_1[0]));    relay_conn far_2_2471_1_b(.in(far_2_2471_0[1]), .out(far_2_2471_1[1]));
    wire [1:0] far_2_2471_2;    relay_conn far_2_2471_2_a(.in(far_2_2471_1[0]), .out(far_2_2471_2[0]));    relay_conn far_2_2471_2_b(.in(far_2_2471_1[1]), .out(far_2_2471_2[1]));
    assign layer_2[431] = far_2_2471_2[0] | far_2_2471_2[1]; 
    wire [1:0] far_2_2472_0;    relay_conn far_2_2472_0_a(.in(layer_1[807]), .out(far_2_2472_0[0]));    relay_conn far_2_2472_0_b(.in(layer_1[903]), .out(far_2_2472_0[1]));
    wire [1:0] far_2_2472_1;    relay_conn far_2_2472_1_a(.in(far_2_2472_0[0]), .out(far_2_2472_1[0]));    relay_conn far_2_2472_1_b(.in(far_2_2472_0[1]), .out(far_2_2472_1[1]));
    wire [1:0] far_2_2472_2;    relay_conn far_2_2472_2_a(.in(far_2_2472_1[0]), .out(far_2_2472_2[0]));    relay_conn far_2_2472_2_b(.in(far_2_2472_1[1]), .out(far_2_2472_2[1]));
    assign layer_2[432] = ~far_2_2472_2[1] | (far_2_2472_2[0] & far_2_2472_2[1]); 
    assign layer_2[433] = ~layer_1[516] | (layer_1[521] & layer_1[516]); 
    wire [1:0] far_2_2474_0;    relay_conn far_2_2474_0_a(.in(layer_1[439]), .out(far_2_2474_0[0]));    relay_conn far_2_2474_0_b(.in(layer_1[312]), .out(far_2_2474_0[1]));
    wire [1:0] far_2_2474_1;    relay_conn far_2_2474_1_a(.in(far_2_2474_0[0]), .out(far_2_2474_1[0]));    relay_conn far_2_2474_1_b(.in(far_2_2474_0[1]), .out(far_2_2474_1[1]));
    wire [1:0] far_2_2474_2;    relay_conn far_2_2474_2_a(.in(far_2_2474_1[0]), .out(far_2_2474_2[0]));    relay_conn far_2_2474_2_b(.in(far_2_2474_1[1]), .out(far_2_2474_2[1]));
    assign layer_2[434] = ~(far_2_2474_2[0] | far_2_2474_2[1]); 
    wire [1:0] far_2_2475_0;    relay_conn far_2_2475_0_a(.in(layer_1[197]), .out(far_2_2475_0[0]));    relay_conn far_2_2475_0_b(.in(layer_1[85]), .out(far_2_2475_0[1]));
    wire [1:0] far_2_2475_1;    relay_conn far_2_2475_1_a(.in(far_2_2475_0[0]), .out(far_2_2475_1[0]));    relay_conn far_2_2475_1_b(.in(far_2_2475_0[1]), .out(far_2_2475_1[1]));
    wire [1:0] far_2_2475_2;    relay_conn far_2_2475_2_a(.in(far_2_2475_1[0]), .out(far_2_2475_2[0]));    relay_conn far_2_2475_2_b(.in(far_2_2475_1[1]), .out(far_2_2475_2[1]));
    assign layer_2[435] = ~far_2_2475_2[1]; 
    wire [1:0] far_2_2476_0;    relay_conn far_2_2476_0_a(.in(layer_1[416]), .out(far_2_2476_0[0]));    relay_conn far_2_2476_0_b(.in(layer_1[498]), .out(far_2_2476_0[1]));
    wire [1:0] far_2_2476_1;    relay_conn far_2_2476_1_a(.in(far_2_2476_0[0]), .out(far_2_2476_1[0]));    relay_conn far_2_2476_1_b(.in(far_2_2476_0[1]), .out(far_2_2476_1[1]));
    assign layer_2[436] = ~(far_2_2476_1[0] | far_2_2476_1[1]); 
    wire [1:0] far_2_2477_0;    relay_conn far_2_2477_0_a(.in(layer_1[619]), .out(far_2_2477_0[0]));    relay_conn far_2_2477_0_b(.in(layer_1[729]), .out(far_2_2477_0[1]));
    wire [1:0] far_2_2477_1;    relay_conn far_2_2477_1_a(.in(far_2_2477_0[0]), .out(far_2_2477_1[0]));    relay_conn far_2_2477_1_b(.in(far_2_2477_0[1]), .out(far_2_2477_1[1]));
    wire [1:0] far_2_2477_2;    relay_conn far_2_2477_2_a(.in(far_2_2477_1[0]), .out(far_2_2477_2[0]));    relay_conn far_2_2477_2_b(.in(far_2_2477_1[1]), .out(far_2_2477_2[1]));
    assign layer_2[437] = ~(far_2_2477_2[0] & far_2_2477_2[1]); 
    wire [1:0] far_2_2478_0;    relay_conn far_2_2478_0_a(.in(layer_1[433]), .out(far_2_2478_0[0]));    relay_conn far_2_2478_0_b(.in(layer_1[542]), .out(far_2_2478_0[1]));
    wire [1:0] far_2_2478_1;    relay_conn far_2_2478_1_a(.in(far_2_2478_0[0]), .out(far_2_2478_1[0]));    relay_conn far_2_2478_1_b(.in(far_2_2478_0[1]), .out(far_2_2478_1[1]));
    wire [1:0] far_2_2478_2;    relay_conn far_2_2478_2_a(.in(far_2_2478_1[0]), .out(far_2_2478_2[0]));    relay_conn far_2_2478_2_b(.in(far_2_2478_1[1]), .out(far_2_2478_2[1]));
    assign layer_2[438] = ~far_2_2478_2[1] | (far_2_2478_2[0] & far_2_2478_2[1]); 
    wire [1:0] far_2_2479_0;    relay_conn far_2_2479_0_a(.in(layer_1[757]), .out(far_2_2479_0[0]));    relay_conn far_2_2479_0_b(.in(layer_1[816]), .out(far_2_2479_0[1]));
    assign layer_2[439] = ~(far_2_2479_0[0] ^ far_2_2479_0[1]); 
    wire [1:0] far_2_2480_0;    relay_conn far_2_2480_0_a(.in(layer_1[303]), .out(far_2_2480_0[0]));    relay_conn far_2_2480_0_b(.in(layer_1[178]), .out(far_2_2480_0[1]));
    wire [1:0] far_2_2480_1;    relay_conn far_2_2480_1_a(.in(far_2_2480_0[0]), .out(far_2_2480_1[0]));    relay_conn far_2_2480_1_b(.in(far_2_2480_0[1]), .out(far_2_2480_1[1]));
    wire [1:0] far_2_2480_2;    relay_conn far_2_2480_2_a(.in(far_2_2480_1[0]), .out(far_2_2480_2[0]));    relay_conn far_2_2480_2_b(.in(far_2_2480_1[1]), .out(far_2_2480_2[1]));
    assign layer_2[440] = ~far_2_2480_2[1] | (far_2_2480_2[0] & far_2_2480_2[1]); 
    wire [1:0] far_2_2481_0;    relay_conn far_2_2481_0_a(.in(layer_1[240]), .out(far_2_2481_0[0]));    relay_conn far_2_2481_0_b(.in(layer_1[280]), .out(far_2_2481_0[1]));
    assign layer_2[441] = far_2_2481_0[0] ^ far_2_2481_0[1]; 
    wire [1:0] far_2_2482_0;    relay_conn far_2_2482_0_a(.in(layer_1[63]), .out(far_2_2482_0[0]));    relay_conn far_2_2482_0_b(.in(layer_1[139]), .out(far_2_2482_0[1]));
    wire [1:0] far_2_2482_1;    relay_conn far_2_2482_1_a(.in(far_2_2482_0[0]), .out(far_2_2482_1[0]));    relay_conn far_2_2482_1_b(.in(far_2_2482_0[1]), .out(far_2_2482_1[1]));
    assign layer_2[442] = ~far_2_2482_1[1] | (far_2_2482_1[0] & far_2_2482_1[1]); 
    assign layer_2[443] = ~layer_1[288] | (layer_1[316] & layer_1[288]); 
    wire [1:0] far_2_2484_0;    relay_conn far_2_2484_0_a(.in(layer_1[342]), .out(far_2_2484_0[0]));    relay_conn far_2_2484_0_b(.in(layer_1[411]), .out(far_2_2484_0[1]));
    wire [1:0] far_2_2484_1;    relay_conn far_2_2484_1_a(.in(far_2_2484_0[0]), .out(far_2_2484_1[0]));    relay_conn far_2_2484_1_b(.in(far_2_2484_0[1]), .out(far_2_2484_1[1]));
    assign layer_2[444] = far_2_2484_1[0]; 
    assign layer_2[445] = layer_1[57] & ~layer_1[44]; 
    wire [1:0] far_2_2486_0;    relay_conn far_2_2486_0_a(.in(layer_1[854]), .out(far_2_2486_0[0]));    relay_conn far_2_2486_0_b(.in(layer_1[814]), .out(far_2_2486_0[1]));
    assign layer_2[446] = ~far_2_2486_0[0]; 
    wire [1:0] far_2_2487_0;    relay_conn far_2_2487_0_a(.in(layer_1[986]), .out(far_2_2487_0[0]));    relay_conn far_2_2487_0_b(.in(layer_1[875]), .out(far_2_2487_0[1]));
    wire [1:0] far_2_2487_1;    relay_conn far_2_2487_1_a(.in(far_2_2487_0[0]), .out(far_2_2487_1[0]));    relay_conn far_2_2487_1_b(.in(far_2_2487_0[1]), .out(far_2_2487_1[1]));
    wire [1:0] far_2_2487_2;    relay_conn far_2_2487_2_a(.in(far_2_2487_1[0]), .out(far_2_2487_2[0]));    relay_conn far_2_2487_2_b(.in(far_2_2487_1[1]), .out(far_2_2487_2[1]));
    assign layer_2[447] = ~far_2_2487_2[0] | (far_2_2487_2[0] & far_2_2487_2[1]); 
    assign layer_2[448] = layer_1[722] & layer_1[743]; 
    wire [1:0] far_2_2489_0;    relay_conn far_2_2489_0_a(.in(layer_1[288]), .out(far_2_2489_0[0]));    relay_conn far_2_2489_0_b(.in(layer_1[341]), .out(far_2_2489_0[1]));
    assign layer_2[449] = ~far_2_2489_0[1] | (far_2_2489_0[0] & far_2_2489_0[1]); 
    assign layer_2[450] = ~layer_1[855]; 
    wire [1:0] far_2_2491_0;    relay_conn far_2_2491_0_a(.in(layer_1[997]), .out(far_2_2491_0[0]));    relay_conn far_2_2491_0_b(.in(layer_1[878]), .out(far_2_2491_0[1]));
    wire [1:0] far_2_2491_1;    relay_conn far_2_2491_1_a(.in(far_2_2491_0[0]), .out(far_2_2491_1[0]));    relay_conn far_2_2491_1_b(.in(far_2_2491_0[1]), .out(far_2_2491_1[1]));
    wire [1:0] far_2_2491_2;    relay_conn far_2_2491_2_a(.in(far_2_2491_1[0]), .out(far_2_2491_2[0]));    relay_conn far_2_2491_2_b(.in(far_2_2491_1[1]), .out(far_2_2491_2[1]));
    assign layer_2[451] = far_2_2491_2[1]; 
    wire [1:0] far_2_2492_0;    relay_conn far_2_2492_0_a(.in(layer_1[716]), .out(far_2_2492_0[0]));    relay_conn far_2_2492_0_b(.in(layer_1[814]), .out(far_2_2492_0[1]));
    wire [1:0] far_2_2492_1;    relay_conn far_2_2492_1_a(.in(far_2_2492_0[0]), .out(far_2_2492_1[0]));    relay_conn far_2_2492_1_b(.in(far_2_2492_0[1]), .out(far_2_2492_1[1]));
    wire [1:0] far_2_2492_2;    relay_conn far_2_2492_2_a(.in(far_2_2492_1[0]), .out(far_2_2492_2[0]));    relay_conn far_2_2492_2_b(.in(far_2_2492_1[1]), .out(far_2_2492_2[1]));
    assign layer_2[452] = ~(far_2_2492_2[0] & far_2_2492_2[1]); 
    wire [1:0] far_2_2493_0;    relay_conn far_2_2493_0_a(.in(layer_1[288]), .out(far_2_2493_0[0]));    relay_conn far_2_2493_0_b(.in(layer_1[217]), .out(far_2_2493_0[1]));
    wire [1:0] far_2_2493_1;    relay_conn far_2_2493_1_a(.in(far_2_2493_0[0]), .out(far_2_2493_1[0]));    relay_conn far_2_2493_1_b(.in(far_2_2493_0[1]), .out(far_2_2493_1[1]));
    assign layer_2[453] = ~far_2_2493_1[1] | (far_2_2493_1[0] & far_2_2493_1[1]); 
    wire [1:0] far_2_2494_0;    relay_conn far_2_2494_0_a(.in(layer_1[952]), .out(far_2_2494_0[0]));    relay_conn far_2_2494_0_b(.in(layer_1[869]), .out(far_2_2494_0[1]));
    wire [1:0] far_2_2494_1;    relay_conn far_2_2494_1_a(.in(far_2_2494_0[0]), .out(far_2_2494_1[0]));    relay_conn far_2_2494_1_b(.in(far_2_2494_0[1]), .out(far_2_2494_1[1]));
    assign layer_2[454] = ~(far_2_2494_1[0] & far_2_2494_1[1]); 
    assign layer_2[455] = ~(layer_1[752] | layer_1[781]); 
    wire [1:0] far_2_2496_0;    relay_conn far_2_2496_0_a(.in(layer_1[363]), .out(far_2_2496_0[0]));    relay_conn far_2_2496_0_b(.in(layer_1[442]), .out(far_2_2496_0[1]));
    wire [1:0] far_2_2496_1;    relay_conn far_2_2496_1_a(.in(far_2_2496_0[0]), .out(far_2_2496_1[0]));    relay_conn far_2_2496_1_b(.in(far_2_2496_0[1]), .out(far_2_2496_1[1]));
    assign layer_2[456] = ~(far_2_2496_1[0] & far_2_2496_1[1]); 
    assign layer_2[457] = layer_1[162] & ~layer_1[188]; 
    assign layer_2[458] = layer_1[25] ^ layer_1[44]; 
    assign layer_2[459] = ~layer_1[31]; 
    wire [1:0] far_2_2500_0;    relay_conn far_2_2500_0_a(.in(layer_1[453]), .out(far_2_2500_0[0]));    relay_conn far_2_2500_0_b(.in(layer_1[390]), .out(far_2_2500_0[1]));
    assign layer_2[460] = far_2_2500_0[1] & ~far_2_2500_0[0]; 
    wire [1:0] far_2_2501_0;    relay_conn far_2_2501_0_a(.in(layer_1[676]), .out(far_2_2501_0[0]));    relay_conn far_2_2501_0_b(.in(layer_1[710]), .out(far_2_2501_0[1]));
    assign layer_2[461] = ~(far_2_2501_0[0] | far_2_2501_0[1]); 
    wire [1:0] far_2_2502_0;    relay_conn far_2_2502_0_a(.in(layer_1[879]), .out(far_2_2502_0[0]));    relay_conn far_2_2502_0_b(.in(layer_1[798]), .out(far_2_2502_0[1]));
    wire [1:0] far_2_2502_1;    relay_conn far_2_2502_1_a(.in(far_2_2502_0[0]), .out(far_2_2502_1[0]));    relay_conn far_2_2502_1_b(.in(far_2_2502_0[1]), .out(far_2_2502_1[1]));
    assign layer_2[462] = ~far_2_2502_1[0] | (far_2_2502_1[0] & far_2_2502_1[1]); 
    assign layer_2[463] = layer_1[958] & ~layer_1[966]; 
    wire [1:0] far_2_2504_0;    relay_conn far_2_2504_0_a(.in(layer_1[233]), .out(far_2_2504_0[0]));    relay_conn far_2_2504_0_b(.in(layer_1[177]), .out(far_2_2504_0[1]));
    assign layer_2[464] = far_2_2504_0[1]; 
    wire [1:0] far_2_2505_0;    relay_conn far_2_2505_0_a(.in(layer_1[646]), .out(far_2_2505_0[0]));    relay_conn far_2_2505_0_b(.in(layer_1[772]), .out(far_2_2505_0[1]));
    wire [1:0] far_2_2505_1;    relay_conn far_2_2505_1_a(.in(far_2_2505_0[0]), .out(far_2_2505_1[0]));    relay_conn far_2_2505_1_b(.in(far_2_2505_0[1]), .out(far_2_2505_1[1]));
    wire [1:0] far_2_2505_2;    relay_conn far_2_2505_2_a(.in(far_2_2505_1[0]), .out(far_2_2505_2[0]));    relay_conn far_2_2505_2_b(.in(far_2_2505_1[1]), .out(far_2_2505_2[1]));
    assign layer_2[465] = far_2_2505_2[0]; 
    wire [1:0] far_2_2506_0;    relay_conn far_2_2506_0_a(.in(layer_1[360]), .out(far_2_2506_0[0]));    relay_conn far_2_2506_0_b(.in(layer_1[409]), .out(far_2_2506_0[1]));
    assign layer_2[466] = far_2_2506_0[1] & ~far_2_2506_0[0]; 
    wire [1:0] far_2_2507_0;    relay_conn far_2_2507_0_a(.in(layer_1[177]), .out(far_2_2507_0[0]));    relay_conn far_2_2507_0_b(.in(layer_1[223]), .out(far_2_2507_0[1]));
    assign layer_2[467] = ~far_2_2507_0[0] | (far_2_2507_0[0] & far_2_2507_0[1]); 
    assign layer_2[468] = layer_1[875] & layer_1[862]; 
    wire [1:0] far_2_2509_0;    relay_conn far_2_2509_0_a(.in(layer_1[180]), .out(far_2_2509_0[0]));    relay_conn far_2_2509_0_b(.in(layer_1[88]), .out(far_2_2509_0[1]));
    wire [1:0] far_2_2509_1;    relay_conn far_2_2509_1_a(.in(far_2_2509_0[0]), .out(far_2_2509_1[0]));    relay_conn far_2_2509_1_b(.in(far_2_2509_0[1]), .out(far_2_2509_1[1]));
    assign layer_2[469] = far_2_2509_1[1] & ~far_2_2509_1[0]; 
    wire [1:0] far_2_2510_0;    relay_conn far_2_2510_0_a(.in(layer_1[918]), .out(far_2_2510_0[0]));    relay_conn far_2_2510_0_b(.in(layer_1[852]), .out(far_2_2510_0[1]));
    wire [1:0] far_2_2510_1;    relay_conn far_2_2510_1_a(.in(far_2_2510_0[0]), .out(far_2_2510_1[0]));    relay_conn far_2_2510_1_b(.in(far_2_2510_0[1]), .out(far_2_2510_1[1]));
    assign layer_2[470] = ~(far_2_2510_1[0] | far_2_2510_1[1]); 
    wire [1:0] far_2_2511_0;    relay_conn far_2_2511_0_a(.in(layer_1[471]), .out(far_2_2511_0[0]));    relay_conn far_2_2511_0_b(.in(layer_1[532]), .out(far_2_2511_0[1]));
    assign layer_2[471] = ~far_2_2511_0[1]; 
    wire [1:0] far_2_2512_0;    relay_conn far_2_2512_0_a(.in(layer_1[391]), .out(far_2_2512_0[0]));    relay_conn far_2_2512_0_b(.in(layer_1[440]), .out(far_2_2512_0[1]));
    assign layer_2[472] = far_2_2512_0[0] & ~far_2_2512_0[1]; 
    assign layer_2[473] = layer_1[95] & ~layer_1[115]; 
    wire [1:0] far_2_2514_0;    relay_conn far_2_2514_0_a(.in(layer_1[655]), .out(far_2_2514_0[0]));    relay_conn far_2_2514_0_b(.in(layer_1[597]), .out(far_2_2514_0[1]));
    assign layer_2[474] = ~(far_2_2514_0[0] & far_2_2514_0[1]); 
    assign layer_2[475] = layer_1[435] & ~layer_1[424]; 
    wire [1:0] far_2_2516_0;    relay_conn far_2_2516_0_a(.in(layer_1[163]), .out(far_2_2516_0[0]));    relay_conn far_2_2516_0_b(.in(layer_1[248]), .out(far_2_2516_0[1]));
    wire [1:0] far_2_2516_1;    relay_conn far_2_2516_1_a(.in(far_2_2516_0[0]), .out(far_2_2516_1[0]));    relay_conn far_2_2516_1_b(.in(far_2_2516_0[1]), .out(far_2_2516_1[1]));
    assign layer_2[476] = ~far_2_2516_1[0]; 
    wire [1:0] far_2_2517_0;    relay_conn far_2_2517_0_a(.in(layer_1[773]), .out(far_2_2517_0[0]));    relay_conn far_2_2517_0_b(.in(layer_1[724]), .out(far_2_2517_0[1]));
    assign layer_2[477] = far_2_2517_0[1]; 
    wire [1:0] far_2_2518_0;    relay_conn far_2_2518_0_a(.in(layer_1[603]), .out(far_2_2518_0[0]));    relay_conn far_2_2518_0_b(.in(layer_1[731]), .out(far_2_2518_0[1]));
    wire [1:0] far_2_2518_1;    relay_conn far_2_2518_1_a(.in(far_2_2518_0[0]), .out(far_2_2518_1[0]));    relay_conn far_2_2518_1_b(.in(far_2_2518_0[1]), .out(far_2_2518_1[1]));
    wire [1:0] far_2_2518_2;    relay_conn far_2_2518_2_a(.in(far_2_2518_1[0]), .out(far_2_2518_2[0]));    relay_conn far_2_2518_2_b(.in(far_2_2518_1[1]), .out(far_2_2518_2[1]));
    wire [1:0] far_2_2518_3;    relay_conn far_2_2518_3_a(.in(far_2_2518_2[0]), .out(far_2_2518_3[0]));    relay_conn far_2_2518_3_b(.in(far_2_2518_2[1]), .out(far_2_2518_3[1]));
    assign layer_2[478] = far_2_2518_3[0]; 
    wire [1:0] far_2_2519_0;    relay_conn far_2_2519_0_a(.in(layer_1[607]), .out(far_2_2519_0[0]));    relay_conn far_2_2519_0_b(.in(layer_1[695]), .out(far_2_2519_0[1]));
    wire [1:0] far_2_2519_1;    relay_conn far_2_2519_1_a(.in(far_2_2519_0[0]), .out(far_2_2519_1[0]));    relay_conn far_2_2519_1_b(.in(far_2_2519_0[1]), .out(far_2_2519_1[1]));
    assign layer_2[479] = far_2_2519_1[1]; 
    assign layer_2[480] = layer_1[84] | layer_1[86]; 
    wire [1:0] far_2_2521_0;    relay_conn far_2_2521_0_a(.in(layer_1[205]), .out(far_2_2521_0[0]));    relay_conn far_2_2521_0_b(.in(layer_1[166]), .out(far_2_2521_0[1]));
    assign layer_2[481] = ~far_2_2521_0[1] | (far_2_2521_0[0] & far_2_2521_0[1]); 
    assign layer_2[482] = ~(layer_1[71] | layer_1[66]); 
    assign layer_2[483] = layer_1[537] | layer_1[562]; 
    wire [1:0] far_2_2524_0;    relay_conn far_2_2524_0_a(.in(layer_1[949]), .out(far_2_2524_0[0]));    relay_conn far_2_2524_0_b(.in(layer_1[1004]), .out(far_2_2524_0[1]));
    assign layer_2[484] = far_2_2524_0[1] & ~far_2_2524_0[0]; 
    wire [1:0] far_2_2525_0;    relay_conn far_2_2525_0_a(.in(layer_1[743]), .out(far_2_2525_0[0]));    relay_conn far_2_2525_0_b(.in(layer_1[775]), .out(far_2_2525_0[1]));
    assign layer_2[485] = ~(far_2_2525_0[0] & far_2_2525_0[1]); 
    wire [1:0] far_2_2526_0;    relay_conn far_2_2526_0_a(.in(layer_1[932]), .out(far_2_2526_0[0]));    relay_conn far_2_2526_0_b(.in(layer_1[965]), .out(far_2_2526_0[1]));
    assign layer_2[486] = ~far_2_2526_0[1]; 
    wire [1:0] far_2_2527_0;    relay_conn far_2_2527_0_a(.in(layer_1[288]), .out(far_2_2527_0[0]));    relay_conn far_2_2527_0_b(.in(layer_1[248]), .out(far_2_2527_0[1]));
    assign layer_2[487] = far_2_2527_0[1] & ~far_2_2527_0[0]; 
    wire [1:0] far_2_2528_0;    relay_conn far_2_2528_0_a(.in(layer_1[274]), .out(far_2_2528_0[0]));    relay_conn far_2_2528_0_b(.in(layer_1[385]), .out(far_2_2528_0[1]));
    wire [1:0] far_2_2528_1;    relay_conn far_2_2528_1_a(.in(far_2_2528_0[0]), .out(far_2_2528_1[0]));    relay_conn far_2_2528_1_b(.in(far_2_2528_0[1]), .out(far_2_2528_1[1]));
    wire [1:0] far_2_2528_2;    relay_conn far_2_2528_2_a(.in(far_2_2528_1[0]), .out(far_2_2528_2[0]));    relay_conn far_2_2528_2_b(.in(far_2_2528_1[1]), .out(far_2_2528_2[1]));
    assign layer_2[488] = far_2_2528_2[0] & far_2_2528_2[1]; 
    wire [1:0] far_2_2529_0;    relay_conn far_2_2529_0_a(.in(layer_1[617]), .out(far_2_2529_0[0]));    relay_conn far_2_2529_0_b(.in(layer_1[689]), .out(far_2_2529_0[1]));
    wire [1:0] far_2_2529_1;    relay_conn far_2_2529_1_a(.in(far_2_2529_0[0]), .out(far_2_2529_1[0]));    relay_conn far_2_2529_1_b(.in(far_2_2529_0[1]), .out(far_2_2529_1[1]));
    assign layer_2[489] = ~(far_2_2529_1[0] & far_2_2529_1[1]); 
    assign layer_2[490] = ~layer_1[331] | (layer_1[331] & layer_1[344]); 
    assign layer_2[491] = ~layer_1[40] | (layer_1[40] & layer_1[39]); 
    wire [1:0] far_2_2532_0;    relay_conn far_2_2532_0_a(.in(layer_1[534]), .out(far_2_2532_0[0]));    relay_conn far_2_2532_0_b(.in(layer_1[466]), .out(far_2_2532_0[1]));
    wire [1:0] far_2_2532_1;    relay_conn far_2_2532_1_a(.in(far_2_2532_0[0]), .out(far_2_2532_1[0]));    relay_conn far_2_2532_1_b(.in(far_2_2532_0[1]), .out(far_2_2532_1[1]));
    assign layer_2[492] = ~(far_2_2532_1[0] & far_2_2532_1[1]); 
    assign layer_2[493] = layer_1[543]; 
    assign layer_2[494] = layer_1[524] & ~layer_1[532]; 
    wire [1:0] far_2_2535_0;    relay_conn far_2_2535_0_a(.in(layer_1[603]), .out(far_2_2535_0[0]));    relay_conn far_2_2535_0_b(.in(layer_1[672]), .out(far_2_2535_0[1]));
    wire [1:0] far_2_2535_1;    relay_conn far_2_2535_1_a(.in(far_2_2535_0[0]), .out(far_2_2535_1[0]));    relay_conn far_2_2535_1_b(.in(far_2_2535_0[1]), .out(far_2_2535_1[1]));
    assign layer_2[495] = ~far_2_2535_1[0] | (far_2_2535_1[0] & far_2_2535_1[1]); 
    wire [1:0] far_2_2536_0;    relay_conn far_2_2536_0_a(.in(layer_1[949]), .out(far_2_2536_0[0]));    relay_conn far_2_2536_0_b(.in(layer_1[874]), .out(far_2_2536_0[1]));
    wire [1:0] far_2_2536_1;    relay_conn far_2_2536_1_a(.in(far_2_2536_0[0]), .out(far_2_2536_1[0]));    relay_conn far_2_2536_1_b(.in(far_2_2536_0[1]), .out(far_2_2536_1[1]));
    assign layer_2[496] = ~(far_2_2536_1[0] | far_2_2536_1[1]); 
    wire [1:0] far_2_2537_0;    relay_conn far_2_2537_0_a(.in(layer_1[12]), .out(far_2_2537_0[0]));    relay_conn far_2_2537_0_b(.in(layer_1[57]), .out(far_2_2537_0[1]));
    assign layer_2[497] = ~far_2_2537_0[1] | (far_2_2537_0[0] & far_2_2537_0[1]); 
    assign layer_2[498] = ~layer_1[918] | (layer_1[941] & layer_1[918]); 
    wire [1:0] far_2_2539_0;    relay_conn far_2_2539_0_a(.in(layer_1[632]), .out(far_2_2539_0[0]));    relay_conn far_2_2539_0_b(.in(layer_1[704]), .out(far_2_2539_0[1]));
    wire [1:0] far_2_2539_1;    relay_conn far_2_2539_1_a(.in(far_2_2539_0[0]), .out(far_2_2539_1[0]));    relay_conn far_2_2539_1_b(.in(far_2_2539_0[1]), .out(far_2_2539_1[1]));
    assign layer_2[499] = far_2_2539_1[0]; 
    wire [1:0] far_2_2540_0;    relay_conn far_2_2540_0_a(.in(layer_1[756]), .out(far_2_2540_0[0]));    relay_conn far_2_2540_0_b(.in(layer_1[826]), .out(far_2_2540_0[1]));
    wire [1:0] far_2_2540_1;    relay_conn far_2_2540_1_a(.in(far_2_2540_0[0]), .out(far_2_2540_1[0]));    relay_conn far_2_2540_1_b(.in(far_2_2540_0[1]), .out(far_2_2540_1[1]));
    assign layer_2[500] = ~far_2_2540_1[0] | (far_2_2540_1[0] & far_2_2540_1[1]); 
    assign layer_2[501] = ~layer_1[632]; 
    wire [1:0] far_2_2542_0;    relay_conn far_2_2542_0_a(.in(layer_1[232]), .out(far_2_2542_0[0]));    relay_conn far_2_2542_0_b(.in(layer_1[317]), .out(far_2_2542_0[1]));
    wire [1:0] far_2_2542_1;    relay_conn far_2_2542_1_a(.in(far_2_2542_0[0]), .out(far_2_2542_1[0]));    relay_conn far_2_2542_1_b(.in(far_2_2542_0[1]), .out(far_2_2542_1[1]));
    assign layer_2[502] = ~(far_2_2542_1[0] & far_2_2542_1[1]); 
    wire [1:0] far_2_2543_0;    relay_conn far_2_2543_0_a(.in(layer_1[542]), .out(far_2_2543_0[0]));    relay_conn far_2_2543_0_b(.in(layer_1[437]), .out(far_2_2543_0[1]));
    wire [1:0] far_2_2543_1;    relay_conn far_2_2543_1_a(.in(far_2_2543_0[0]), .out(far_2_2543_1[0]));    relay_conn far_2_2543_1_b(.in(far_2_2543_0[1]), .out(far_2_2543_1[1]));
    wire [1:0] far_2_2543_2;    relay_conn far_2_2543_2_a(.in(far_2_2543_1[0]), .out(far_2_2543_2[0]));    relay_conn far_2_2543_2_b(.in(far_2_2543_1[1]), .out(far_2_2543_2[1]));
    assign layer_2[503] = ~far_2_2543_2[1] | (far_2_2543_2[0] & far_2_2543_2[1]); 
    wire [1:0] far_2_2544_0;    relay_conn far_2_2544_0_a(.in(layer_1[106]), .out(far_2_2544_0[0]));    relay_conn far_2_2544_0_b(.in(layer_1[158]), .out(far_2_2544_0[1]));
    assign layer_2[504] = ~far_2_2544_0[1] | (far_2_2544_0[0] & far_2_2544_0[1]); 
    wire [1:0] far_2_2545_0;    relay_conn far_2_2545_0_a(.in(layer_1[795]), .out(far_2_2545_0[0]));    relay_conn far_2_2545_0_b(.in(layer_1[916]), .out(far_2_2545_0[1]));
    wire [1:0] far_2_2545_1;    relay_conn far_2_2545_1_a(.in(far_2_2545_0[0]), .out(far_2_2545_1[0]));    relay_conn far_2_2545_1_b(.in(far_2_2545_0[1]), .out(far_2_2545_1[1]));
    wire [1:0] far_2_2545_2;    relay_conn far_2_2545_2_a(.in(far_2_2545_1[0]), .out(far_2_2545_2[0]));    relay_conn far_2_2545_2_b(.in(far_2_2545_1[1]), .out(far_2_2545_2[1]));
    assign layer_2[505] = far_2_2545_2[1]; 
    assign layer_2[506] = layer_1[558] ^ layer_1[555]; 
    wire [1:0] far_2_2547_0;    relay_conn far_2_2547_0_a(.in(layer_1[213]), .out(far_2_2547_0[0]));    relay_conn far_2_2547_0_b(.in(layer_1[139]), .out(far_2_2547_0[1]));
    wire [1:0] far_2_2547_1;    relay_conn far_2_2547_1_a(.in(far_2_2547_0[0]), .out(far_2_2547_1[0]));    relay_conn far_2_2547_1_b(.in(far_2_2547_0[1]), .out(far_2_2547_1[1]));
    assign layer_2[507] = far_2_2547_1[0] ^ far_2_2547_1[1]; 
    assign layer_2[508] = ~layer_1[619]; 
    wire [1:0] far_2_2549_0;    relay_conn far_2_2549_0_a(.in(layer_1[688]), .out(far_2_2549_0[0]));    relay_conn far_2_2549_0_b(.in(layer_1[780]), .out(far_2_2549_0[1]));
    wire [1:0] far_2_2549_1;    relay_conn far_2_2549_1_a(.in(far_2_2549_0[0]), .out(far_2_2549_1[0]));    relay_conn far_2_2549_1_b(.in(far_2_2549_0[1]), .out(far_2_2549_1[1]));
    assign layer_2[509] = far_2_2549_1[1]; 
    assign layer_2[510] = layer_1[918]; 
    wire [1:0] far_2_2551_0;    relay_conn far_2_2551_0_a(.in(layer_1[248]), .out(far_2_2551_0[0]));    relay_conn far_2_2551_0_b(.in(layer_1[204]), .out(far_2_2551_0[1]));
    assign layer_2[511] = far_2_2551_0[0]; 
    wire [1:0] far_2_2552_0;    relay_conn far_2_2552_0_a(.in(layer_1[285]), .out(far_2_2552_0[0]));    relay_conn far_2_2552_0_b(.in(layer_1[238]), .out(far_2_2552_0[1]));
    assign layer_2[512] = far_2_2552_0[0] & ~far_2_2552_0[1]; 
    wire [1:0] far_2_2553_0;    relay_conn far_2_2553_0_a(.in(layer_1[983]), .out(far_2_2553_0[0]));    relay_conn far_2_2553_0_b(.in(layer_1[932]), .out(far_2_2553_0[1]));
    assign layer_2[513] = far_2_2553_0[0] & far_2_2553_0[1]; 
    assign layer_2[514] = layer_1[767]; 
    wire [1:0] far_2_2555_0;    relay_conn far_2_2555_0_a(.in(layer_1[426]), .out(far_2_2555_0[0]));    relay_conn far_2_2555_0_b(.in(layer_1[316]), .out(far_2_2555_0[1]));
    wire [1:0] far_2_2555_1;    relay_conn far_2_2555_1_a(.in(far_2_2555_0[0]), .out(far_2_2555_1[0]));    relay_conn far_2_2555_1_b(.in(far_2_2555_0[1]), .out(far_2_2555_1[1]));
    wire [1:0] far_2_2555_2;    relay_conn far_2_2555_2_a(.in(far_2_2555_1[0]), .out(far_2_2555_2[0]));    relay_conn far_2_2555_2_b(.in(far_2_2555_1[1]), .out(far_2_2555_2[1]));
    assign layer_2[515] = ~far_2_2555_2[1]; 
    wire [1:0] far_2_2556_0;    relay_conn far_2_2556_0_a(.in(layer_1[596]), .out(far_2_2556_0[0]));    relay_conn far_2_2556_0_b(.in(layer_1[664]), .out(far_2_2556_0[1]));
    wire [1:0] far_2_2556_1;    relay_conn far_2_2556_1_a(.in(far_2_2556_0[0]), .out(far_2_2556_1[0]));    relay_conn far_2_2556_1_b(.in(far_2_2556_0[1]), .out(far_2_2556_1[1]));
    assign layer_2[516] = ~far_2_2556_1[0]; 
    wire [1:0] far_2_2557_0;    relay_conn far_2_2557_0_a(.in(layer_1[192]), .out(far_2_2557_0[0]));    relay_conn far_2_2557_0_b(.in(layer_1[248]), .out(far_2_2557_0[1]));
    assign layer_2[517] = far_2_2557_0[1]; 
    wire [1:0] far_2_2558_0;    relay_conn far_2_2558_0_a(.in(layer_1[349]), .out(far_2_2558_0[0]));    relay_conn far_2_2558_0_b(.in(layer_1[311]), .out(far_2_2558_0[1]));
    assign layer_2[518] = far_2_2558_0[0]; 
    wire [1:0] far_2_2559_0;    relay_conn far_2_2559_0_a(.in(layer_1[125]), .out(far_2_2559_0[0]));    relay_conn far_2_2559_0_b(.in(layer_1[239]), .out(far_2_2559_0[1]));
    wire [1:0] far_2_2559_1;    relay_conn far_2_2559_1_a(.in(far_2_2559_0[0]), .out(far_2_2559_1[0]));    relay_conn far_2_2559_1_b(.in(far_2_2559_0[1]), .out(far_2_2559_1[1]));
    wire [1:0] far_2_2559_2;    relay_conn far_2_2559_2_a(.in(far_2_2559_1[0]), .out(far_2_2559_2[0]));    relay_conn far_2_2559_2_b(.in(far_2_2559_1[1]), .out(far_2_2559_2[1]));
    assign layer_2[519] = ~(far_2_2559_2[0] & far_2_2559_2[1]); 
    assign layer_2[520] = ~layer_1[772] | (layer_1[772] & layer_1[743]); 
    wire [1:0] far_2_2561_0;    relay_conn far_2_2561_0_a(.in(layer_1[910]), .out(far_2_2561_0[0]));    relay_conn far_2_2561_0_b(.in(layer_1[1015]), .out(far_2_2561_0[1]));
    wire [1:0] far_2_2561_1;    relay_conn far_2_2561_1_a(.in(far_2_2561_0[0]), .out(far_2_2561_1[0]));    relay_conn far_2_2561_1_b(.in(far_2_2561_0[1]), .out(far_2_2561_1[1]));
    wire [1:0] far_2_2561_2;    relay_conn far_2_2561_2_a(.in(far_2_2561_1[0]), .out(far_2_2561_2[0]));    relay_conn far_2_2561_2_b(.in(far_2_2561_1[1]), .out(far_2_2561_2[1]));
    assign layer_2[521] = ~far_2_2561_2[0] | (far_2_2561_2[0] & far_2_2561_2[1]); 
    wire [1:0] far_2_2562_0;    relay_conn far_2_2562_0_a(.in(layer_1[728]), .out(far_2_2562_0[0]));    relay_conn far_2_2562_0_b(.in(layer_1[652]), .out(far_2_2562_0[1]));
    wire [1:0] far_2_2562_1;    relay_conn far_2_2562_1_a(.in(far_2_2562_0[0]), .out(far_2_2562_1[0]));    relay_conn far_2_2562_1_b(.in(far_2_2562_0[1]), .out(far_2_2562_1[1]));
    assign layer_2[522] = far_2_2562_1[0] & ~far_2_2562_1[1]; 
    assign layer_2[523] = ~layer_1[409] | (layer_1[409] & layer_1[405]); 
    wire [1:0] far_2_2564_0;    relay_conn far_2_2564_0_a(.in(layer_1[521]), .out(far_2_2564_0[0]));    relay_conn far_2_2564_0_b(.in(layer_1[609]), .out(far_2_2564_0[1]));
    wire [1:0] far_2_2564_1;    relay_conn far_2_2564_1_a(.in(far_2_2564_0[0]), .out(far_2_2564_1[0]));    relay_conn far_2_2564_1_b(.in(far_2_2564_0[1]), .out(far_2_2564_1[1]));
    assign layer_2[524] = far_2_2564_1[1]; 
    wire [1:0] far_2_2565_0;    relay_conn far_2_2565_0_a(.in(layer_1[190]), .out(far_2_2565_0[0]));    relay_conn far_2_2565_0_b(.in(layer_1[262]), .out(far_2_2565_0[1]));
    wire [1:0] far_2_2565_1;    relay_conn far_2_2565_1_a(.in(far_2_2565_0[0]), .out(far_2_2565_1[0]));    relay_conn far_2_2565_1_b(.in(far_2_2565_0[1]), .out(far_2_2565_1[1]));
    assign layer_2[525] = ~(far_2_2565_1[0] & far_2_2565_1[1]); 
    assign layer_2[526] = ~layer_1[333]; 
    wire [1:0] far_2_2567_0;    relay_conn far_2_2567_0_a(.in(layer_1[400]), .out(far_2_2567_0[0]));    relay_conn far_2_2567_0_b(.in(layer_1[446]), .out(far_2_2567_0[1]));
    assign layer_2[527] = ~far_2_2567_0[0] | (far_2_2567_0[0] & far_2_2567_0[1]); 
    assign layer_2[528] = ~(layer_1[64] | layer_1[83]); 
    wire [1:0] far_2_2569_0;    relay_conn far_2_2569_0_a(.in(layer_1[646]), .out(far_2_2569_0[0]));    relay_conn far_2_2569_0_b(.in(layer_1[682]), .out(far_2_2569_0[1]));
    assign layer_2[529] = far_2_2569_0[0] & ~far_2_2569_0[1]; 
    wire [1:0] far_2_2570_0;    relay_conn far_2_2570_0_a(.in(layer_1[682]), .out(far_2_2570_0[0]));    relay_conn far_2_2570_0_b(.in(layer_1[742]), .out(far_2_2570_0[1]));
    assign layer_2[530] = far_2_2570_0[0] ^ far_2_2570_0[1]; 
    wire [1:0] far_2_2571_0;    relay_conn far_2_2571_0_a(.in(layer_1[255]), .out(far_2_2571_0[0]));    relay_conn far_2_2571_0_b(.in(layer_1[336]), .out(far_2_2571_0[1]));
    wire [1:0] far_2_2571_1;    relay_conn far_2_2571_1_a(.in(far_2_2571_0[0]), .out(far_2_2571_1[0]));    relay_conn far_2_2571_1_b(.in(far_2_2571_0[1]), .out(far_2_2571_1[1]));
    assign layer_2[531] = far_2_2571_1[0] & ~far_2_2571_1[1]; 
    wire [1:0] far_2_2572_0;    relay_conn far_2_2572_0_a(.in(layer_1[771]), .out(far_2_2572_0[0]));    relay_conn far_2_2572_0_b(.in(layer_1[715]), .out(far_2_2572_0[1]));
    assign layer_2[532] = far_2_2572_0[1] & ~far_2_2572_0[0]; 
    assign layer_2[533] = ~(layer_1[527] ^ layer_1[498]); 
    wire [1:0] far_2_2574_0;    relay_conn far_2_2574_0_a(.in(layer_1[722]), .out(far_2_2574_0[0]));    relay_conn far_2_2574_0_b(.in(layer_1[816]), .out(far_2_2574_0[1]));
    wire [1:0] far_2_2574_1;    relay_conn far_2_2574_1_a(.in(far_2_2574_0[0]), .out(far_2_2574_1[0]));    relay_conn far_2_2574_1_b(.in(far_2_2574_0[1]), .out(far_2_2574_1[1]));
    assign layer_2[534] = far_2_2574_1[0] & ~far_2_2574_1[1]; 
    wire [1:0] far_2_2575_0;    relay_conn far_2_2575_0_a(.in(layer_1[188]), .out(far_2_2575_0[0]));    relay_conn far_2_2575_0_b(.in(layer_1[265]), .out(far_2_2575_0[1]));
    wire [1:0] far_2_2575_1;    relay_conn far_2_2575_1_a(.in(far_2_2575_0[0]), .out(far_2_2575_1[0]));    relay_conn far_2_2575_1_b(.in(far_2_2575_0[1]), .out(far_2_2575_1[1]));
    assign layer_2[535] = far_2_2575_1[0] & ~far_2_2575_1[1]; 
    wire [1:0] far_2_2576_0;    relay_conn far_2_2576_0_a(.in(layer_1[721]), .out(far_2_2576_0[0]));    relay_conn far_2_2576_0_b(.in(layer_1[594]), .out(far_2_2576_0[1]));
    wire [1:0] far_2_2576_1;    relay_conn far_2_2576_1_a(.in(far_2_2576_0[0]), .out(far_2_2576_1[0]));    relay_conn far_2_2576_1_b(.in(far_2_2576_0[1]), .out(far_2_2576_1[1]));
    wire [1:0] far_2_2576_2;    relay_conn far_2_2576_2_a(.in(far_2_2576_1[0]), .out(far_2_2576_2[0]));    relay_conn far_2_2576_2_b(.in(far_2_2576_1[1]), .out(far_2_2576_2[1]));
    assign layer_2[536] = ~far_2_2576_2[1]; 
    wire [1:0] far_2_2577_0;    relay_conn far_2_2577_0_a(.in(layer_1[115]), .out(far_2_2577_0[0]));    relay_conn far_2_2577_0_b(.in(layer_1[55]), .out(far_2_2577_0[1]));
    assign layer_2[537] = ~(far_2_2577_0[0] ^ far_2_2577_0[1]); 
    wire [1:0] far_2_2578_0;    relay_conn far_2_2578_0_a(.in(layer_1[352]), .out(far_2_2578_0[0]));    relay_conn far_2_2578_0_b(.in(layer_1[303]), .out(far_2_2578_0[1]));
    assign layer_2[538] = far_2_2578_0[0] | far_2_2578_0[1]; 
    wire [1:0] far_2_2579_0;    relay_conn far_2_2579_0_a(.in(layer_1[364]), .out(far_2_2579_0[0]));    relay_conn far_2_2579_0_b(.in(layer_1[409]), .out(far_2_2579_0[1]));
    assign layer_2[539] = ~(far_2_2579_0[0] | far_2_2579_0[1]); 
    wire [1:0] far_2_2580_0;    relay_conn far_2_2580_0_a(.in(layer_1[622]), .out(far_2_2580_0[0]));    relay_conn far_2_2580_0_b(.in(layer_1[724]), .out(far_2_2580_0[1]));
    wire [1:0] far_2_2580_1;    relay_conn far_2_2580_1_a(.in(far_2_2580_0[0]), .out(far_2_2580_1[0]));    relay_conn far_2_2580_1_b(.in(far_2_2580_0[1]), .out(far_2_2580_1[1]));
    wire [1:0] far_2_2580_2;    relay_conn far_2_2580_2_a(.in(far_2_2580_1[0]), .out(far_2_2580_2[0]));    relay_conn far_2_2580_2_b(.in(far_2_2580_1[1]), .out(far_2_2580_2[1]));
    assign layer_2[540] = ~far_2_2580_2[1] | (far_2_2580_2[0] & far_2_2580_2[1]); 
    wire [1:0] far_2_2581_0;    relay_conn far_2_2581_0_a(.in(layer_1[1002]), .out(far_2_2581_0[0]));    relay_conn far_2_2581_0_b(.in(layer_1[960]), .out(far_2_2581_0[1]));
    assign layer_2[541] = ~far_2_2581_0[0] | (far_2_2581_0[0] & far_2_2581_0[1]); 
    wire [1:0] far_2_2582_0;    relay_conn far_2_2582_0_a(.in(layer_1[1000]), .out(far_2_2582_0[0]));    relay_conn far_2_2582_0_b(.in(layer_1[897]), .out(far_2_2582_0[1]));
    wire [1:0] far_2_2582_1;    relay_conn far_2_2582_1_a(.in(far_2_2582_0[0]), .out(far_2_2582_1[0]));    relay_conn far_2_2582_1_b(.in(far_2_2582_0[1]), .out(far_2_2582_1[1]));
    wire [1:0] far_2_2582_2;    relay_conn far_2_2582_2_a(.in(far_2_2582_1[0]), .out(far_2_2582_2[0]));    relay_conn far_2_2582_2_b(.in(far_2_2582_1[1]), .out(far_2_2582_2[1]));
    assign layer_2[542] = far_2_2582_2[0] ^ far_2_2582_2[1]; 
    assign layer_2[543] = layer_1[192] | layer_1[204]; 
    wire [1:0] far_2_2584_0;    relay_conn far_2_2584_0_a(.in(layer_1[133]), .out(far_2_2584_0[0]));    relay_conn far_2_2584_0_b(.in(layer_1[48]), .out(far_2_2584_0[1]));
    wire [1:0] far_2_2584_1;    relay_conn far_2_2584_1_a(.in(far_2_2584_0[0]), .out(far_2_2584_1[0]));    relay_conn far_2_2584_1_b(.in(far_2_2584_0[1]), .out(far_2_2584_1[1]));
    assign layer_2[544] = ~(far_2_2584_1[0] & far_2_2584_1[1]); 
    wire [1:0] far_2_2585_0;    relay_conn far_2_2585_0_a(.in(layer_1[962]), .out(far_2_2585_0[0]));    relay_conn far_2_2585_0_b(.in(layer_1[864]), .out(far_2_2585_0[1]));
    wire [1:0] far_2_2585_1;    relay_conn far_2_2585_1_a(.in(far_2_2585_0[0]), .out(far_2_2585_1[0]));    relay_conn far_2_2585_1_b(.in(far_2_2585_0[1]), .out(far_2_2585_1[1]));
    wire [1:0] far_2_2585_2;    relay_conn far_2_2585_2_a(.in(far_2_2585_1[0]), .out(far_2_2585_2[0]));    relay_conn far_2_2585_2_b(.in(far_2_2585_1[1]), .out(far_2_2585_2[1]));
    assign layer_2[545] = far_2_2585_2[0] | far_2_2585_2[1]; 
    wire [1:0] far_2_2586_0;    relay_conn far_2_2586_0_a(.in(layer_1[532]), .out(far_2_2586_0[0]));    relay_conn far_2_2586_0_b(.in(layer_1[603]), .out(far_2_2586_0[1]));
    wire [1:0] far_2_2586_1;    relay_conn far_2_2586_1_a(.in(far_2_2586_0[0]), .out(far_2_2586_1[0]));    relay_conn far_2_2586_1_b(.in(far_2_2586_0[1]), .out(far_2_2586_1[1]));
    assign layer_2[546] = far_2_2586_1[0] | far_2_2586_1[1]; 
    wire [1:0] far_2_2587_0;    relay_conn far_2_2587_0_a(.in(layer_1[532]), .out(far_2_2587_0[0]));    relay_conn far_2_2587_0_b(.in(layer_1[404]), .out(far_2_2587_0[1]));
    wire [1:0] far_2_2587_1;    relay_conn far_2_2587_1_a(.in(far_2_2587_0[0]), .out(far_2_2587_1[0]));    relay_conn far_2_2587_1_b(.in(far_2_2587_0[1]), .out(far_2_2587_1[1]));
    wire [1:0] far_2_2587_2;    relay_conn far_2_2587_2_a(.in(far_2_2587_1[0]), .out(far_2_2587_2[0]));    relay_conn far_2_2587_2_b(.in(far_2_2587_1[1]), .out(far_2_2587_2[1]));
    wire [1:0] far_2_2587_3;    relay_conn far_2_2587_3_a(.in(far_2_2587_2[0]), .out(far_2_2587_3[0]));    relay_conn far_2_2587_3_b(.in(far_2_2587_2[1]), .out(far_2_2587_3[1]));
    assign layer_2[547] = far_2_2587_3[0]; 
    assign layer_2[548] = ~(layer_1[353] | layer_1[349]); 
    wire [1:0] far_2_2589_0;    relay_conn far_2_2589_0_a(.in(layer_1[5]), .out(far_2_2589_0[0]));    relay_conn far_2_2589_0_b(.in(layer_1[45]), .out(far_2_2589_0[1]));
    assign layer_2[549] = ~(far_2_2589_0[0] | far_2_2589_0[1]); 
    wire [1:0] far_2_2590_0;    relay_conn far_2_2590_0_a(.in(layer_1[710]), .out(far_2_2590_0[0]));    relay_conn far_2_2590_0_b(.in(layer_1[646]), .out(far_2_2590_0[1]));
    wire [1:0] far_2_2590_1;    relay_conn far_2_2590_1_a(.in(far_2_2590_0[0]), .out(far_2_2590_1[0]));    relay_conn far_2_2590_1_b(.in(far_2_2590_0[1]), .out(far_2_2590_1[1]));
    assign layer_2[550] = ~far_2_2590_1[1]; 
    wire [1:0] far_2_2591_0;    relay_conn far_2_2591_0_a(.in(layer_1[280]), .out(far_2_2591_0[0]));    relay_conn far_2_2591_0_b(.in(layer_1[391]), .out(far_2_2591_0[1]));
    wire [1:0] far_2_2591_1;    relay_conn far_2_2591_1_a(.in(far_2_2591_0[0]), .out(far_2_2591_1[0]));    relay_conn far_2_2591_1_b(.in(far_2_2591_0[1]), .out(far_2_2591_1[1]));
    wire [1:0] far_2_2591_2;    relay_conn far_2_2591_2_a(.in(far_2_2591_1[0]), .out(far_2_2591_2[0]));    relay_conn far_2_2591_2_b(.in(far_2_2591_1[1]), .out(far_2_2591_2[1]));
    assign layer_2[551] = far_2_2591_2[1]; 
    wire [1:0] far_2_2592_0;    relay_conn far_2_2592_0_a(.in(layer_1[439]), .out(far_2_2592_0[0]));    relay_conn far_2_2592_0_b(.in(layer_1[350]), .out(far_2_2592_0[1]));
    wire [1:0] far_2_2592_1;    relay_conn far_2_2592_1_a(.in(far_2_2592_0[0]), .out(far_2_2592_1[0]));    relay_conn far_2_2592_1_b(.in(far_2_2592_0[1]), .out(far_2_2592_1[1]));
    assign layer_2[552] = ~far_2_2592_1[0]; 
    wire [1:0] far_2_2593_0;    relay_conn far_2_2593_0_a(.in(layer_1[153]), .out(far_2_2593_0[0]));    relay_conn far_2_2593_0_b(.in(layer_1[281]), .out(far_2_2593_0[1]));
    wire [1:0] far_2_2593_1;    relay_conn far_2_2593_1_a(.in(far_2_2593_0[0]), .out(far_2_2593_1[0]));    relay_conn far_2_2593_1_b(.in(far_2_2593_0[1]), .out(far_2_2593_1[1]));
    wire [1:0] far_2_2593_2;    relay_conn far_2_2593_2_a(.in(far_2_2593_1[0]), .out(far_2_2593_2[0]));    relay_conn far_2_2593_2_b(.in(far_2_2593_1[1]), .out(far_2_2593_2[1]));
    wire [1:0] far_2_2593_3;    relay_conn far_2_2593_3_a(.in(far_2_2593_2[0]), .out(far_2_2593_3[0]));    relay_conn far_2_2593_3_b(.in(far_2_2593_2[1]), .out(far_2_2593_3[1]));
    assign layer_2[553] = far_2_2593_3[1]; 
    assign layer_2[554] = layer_1[427]; 
    wire [1:0] far_2_2595_0;    relay_conn far_2_2595_0_a(.in(layer_1[157]), .out(far_2_2595_0[0]));    relay_conn far_2_2595_0_b(.in(layer_1[203]), .out(far_2_2595_0[1]));
    assign layer_2[555] = ~(far_2_2595_0[0] ^ far_2_2595_0[1]); 
    wire [1:0] far_2_2596_0;    relay_conn far_2_2596_0_a(.in(layer_1[691]), .out(far_2_2596_0[0]));    relay_conn far_2_2596_0_b(.in(layer_1[617]), .out(far_2_2596_0[1]));
    wire [1:0] far_2_2596_1;    relay_conn far_2_2596_1_a(.in(far_2_2596_0[0]), .out(far_2_2596_1[0]));    relay_conn far_2_2596_1_b(.in(far_2_2596_0[1]), .out(far_2_2596_1[1]));
    assign layer_2[556] = far_2_2596_1[1] & ~far_2_2596_1[0]; 
    wire [1:0] far_2_2597_0;    relay_conn far_2_2597_0_a(.in(layer_1[997]), .out(far_2_2597_0[0]));    relay_conn far_2_2597_0_b(.in(layer_1[934]), .out(far_2_2597_0[1]));
    assign layer_2[557] = ~(far_2_2597_0[0] ^ far_2_2597_0[1]); 
    assign layer_2[558] = ~layer_1[874] | (layer_1[854] & layer_1[874]); 
    wire [1:0] far_2_2599_0;    relay_conn far_2_2599_0_a(.in(layer_1[319]), .out(far_2_2599_0[0]));    relay_conn far_2_2599_0_b(.in(layer_1[267]), .out(far_2_2599_0[1]));
    assign layer_2[559] = ~far_2_2599_0[0]; 
    wire [1:0] far_2_2600_0;    relay_conn far_2_2600_0_a(.in(layer_1[177]), .out(far_2_2600_0[0]));    relay_conn far_2_2600_0_b(.in(layer_1[93]), .out(far_2_2600_0[1]));
    wire [1:0] far_2_2600_1;    relay_conn far_2_2600_1_a(.in(far_2_2600_0[0]), .out(far_2_2600_1[0]));    relay_conn far_2_2600_1_b(.in(far_2_2600_0[1]), .out(far_2_2600_1[1]));
    assign layer_2[560] = far_2_2600_1[0]; 
    wire [1:0] far_2_2601_0;    relay_conn far_2_2601_0_a(.in(layer_1[502]), .out(far_2_2601_0[0]));    relay_conn far_2_2601_0_b(.in(layer_1[400]), .out(far_2_2601_0[1]));
    wire [1:0] far_2_2601_1;    relay_conn far_2_2601_1_a(.in(far_2_2601_0[0]), .out(far_2_2601_1[0]));    relay_conn far_2_2601_1_b(.in(far_2_2601_0[1]), .out(far_2_2601_1[1]));
    wire [1:0] far_2_2601_2;    relay_conn far_2_2601_2_a(.in(far_2_2601_1[0]), .out(far_2_2601_2[0]));    relay_conn far_2_2601_2_b(.in(far_2_2601_1[1]), .out(far_2_2601_2[1]));
    assign layer_2[561] = far_2_2601_2[0] | far_2_2601_2[1]; 
    assign layer_2[562] = ~layer_1[207] | (layer_1[210] & layer_1[207]); 
    wire [1:0] far_2_2603_0;    relay_conn far_2_2603_0_a(.in(layer_1[520]), .out(far_2_2603_0[0]));    relay_conn far_2_2603_0_b(.in(layer_1[617]), .out(far_2_2603_0[1]));
    wire [1:0] far_2_2603_1;    relay_conn far_2_2603_1_a(.in(far_2_2603_0[0]), .out(far_2_2603_1[0]));    relay_conn far_2_2603_1_b(.in(far_2_2603_0[1]), .out(far_2_2603_1[1]));
    wire [1:0] far_2_2603_2;    relay_conn far_2_2603_2_a(.in(far_2_2603_1[0]), .out(far_2_2603_2[0]));    relay_conn far_2_2603_2_b(.in(far_2_2603_1[1]), .out(far_2_2603_2[1]));
    assign layer_2[563] = far_2_2603_2[0] ^ far_2_2603_2[1]; 
    wire [1:0] far_2_2604_0;    relay_conn far_2_2604_0_a(.in(layer_1[980]), .out(far_2_2604_0[0]));    relay_conn far_2_2604_0_b(.in(layer_1[863]), .out(far_2_2604_0[1]));
    wire [1:0] far_2_2604_1;    relay_conn far_2_2604_1_a(.in(far_2_2604_0[0]), .out(far_2_2604_1[0]));    relay_conn far_2_2604_1_b(.in(far_2_2604_0[1]), .out(far_2_2604_1[1]));
    wire [1:0] far_2_2604_2;    relay_conn far_2_2604_2_a(.in(far_2_2604_1[0]), .out(far_2_2604_2[0]));    relay_conn far_2_2604_2_b(.in(far_2_2604_1[1]), .out(far_2_2604_2[1]));
    assign layer_2[564] = ~far_2_2604_2[0]; 
    assign layer_2[565] = ~layer_1[124] | (layer_1[127] & layer_1[124]); 
    wire [1:0] far_2_2606_0;    relay_conn far_2_2606_0_a(.in(layer_1[765]), .out(far_2_2606_0[0]));    relay_conn far_2_2606_0_b(.in(layer_1[891]), .out(far_2_2606_0[1]));
    wire [1:0] far_2_2606_1;    relay_conn far_2_2606_1_a(.in(far_2_2606_0[0]), .out(far_2_2606_1[0]));    relay_conn far_2_2606_1_b(.in(far_2_2606_0[1]), .out(far_2_2606_1[1]));
    wire [1:0] far_2_2606_2;    relay_conn far_2_2606_2_a(.in(far_2_2606_1[0]), .out(far_2_2606_2[0]));    relay_conn far_2_2606_2_b(.in(far_2_2606_1[1]), .out(far_2_2606_2[1]));
    assign layer_2[566] = ~far_2_2606_2[0]; 
    wire [1:0] far_2_2607_0;    relay_conn far_2_2607_0_a(.in(layer_1[892]), .out(far_2_2607_0[0]));    relay_conn far_2_2607_0_b(.in(layer_1[941]), .out(far_2_2607_0[1]));
    assign layer_2[567] = ~far_2_2607_0[0] | (far_2_2607_0[0] & far_2_2607_0[1]); 
    wire [1:0] far_2_2608_0;    relay_conn far_2_2608_0_a(.in(layer_1[676]), .out(far_2_2608_0[0]));    relay_conn far_2_2608_0_b(.in(layer_1[621]), .out(far_2_2608_0[1]));
    assign layer_2[568] = far_2_2608_0[0]; 
    wire [1:0] far_2_2609_0;    relay_conn far_2_2609_0_a(.in(layer_1[768]), .out(far_2_2609_0[0]));    relay_conn far_2_2609_0_b(.in(layer_1[689]), .out(far_2_2609_0[1]));
    wire [1:0] far_2_2609_1;    relay_conn far_2_2609_1_a(.in(far_2_2609_0[0]), .out(far_2_2609_1[0]));    relay_conn far_2_2609_1_b(.in(far_2_2609_0[1]), .out(far_2_2609_1[1]));
    assign layer_2[569] = ~far_2_2609_1[1]; 
    assign layer_2[570] = layer_1[617] & layer_1[597]; 
    assign layer_2[571] = ~(layer_1[462] & layer_1[459]); 
    wire [1:0] far_2_2612_0;    relay_conn far_2_2612_0_a(.in(layer_1[779]), .out(far_2_2612_0[0]));    relay_conn far_2_2612_0_b(.in(layer_1[875]), .out(far_2_2612_0[1]));
    wire [1:0] far_2_2612_1;    relay_conn far_2_2612_1_a(.in(far_2_2612_0[0]), .out(far_2_2612_1[0]));    relay_conn far_2_2612_1_b(.in(far_2_2612_0[1]), .out(far_2_2612_1[1]));
    wire [1:0] far_2_2612_2;    relay_conn far_2_2612_2_a(.in(far_2_2612_1[0]), .out(far_2_2612_2[0]));    relay_conn far_2_2612_2_b(.in(far_2_2612_1[1]), .out(far_2_2612_2[1]));
    assign layer_2[572] = ~(far_2_2612_2[0] & far_2_2612_2[1]); 
    wire [1:0] far_2_2613_0;    relay_conn far_2_2613_0_a(.in(layer_1[596]), .out(far_2_2613_0[0]));    relay_conn far_2_2613_0_b(.in(layer_1[513]), .out(far_2_2613_0[1]));
    wire [1:0] far_2_2613_1;    relay_conn far_2_2613_1_a(.in(far_2_2613_0[0]), .out(far_2_2613_1[0]));    relay_conn far_2_2613_1_b(.in(far_2_2613_0[1]), .out(far_2_2613_1[1]));
    assign layer_2[573] = ~far_2_2613_1[1]; 
    wire [1:0] far_2_2614_0;    relay_conn far_2_2614_0_a(.in(layer_1[807]), .out(far_2_2614_0[0]));    relay_conn far_2_2614_0_b(.in(layer_1[926]), .out(far_2_2614_0[1]));
    wire [1:0] far_2_2614_1;    relay_conn far_2_2614_1_a(.in(far_2_2614_0[0]), .out(far_2_2614_1[0]));    relay_conn far_2_2614_1_b(.in(far_2_2614_0[1]), .out(far_2_2614_1[1]));
    wire [1:0] far_2_2614_2;    relay_conn far_2_2614_2_a(.in(far_2_2614_1[0]), .out(far_2_2614_2[0]));    relay_conn far_2_2614_2_b(.in(far_2_2614_1[1]), .out(far_2_2614_2[1]));
    assign layer_2[574] = far_2_2614_2[0] ^ far_2_2614_2[1]; 
    assign layer_2[575] = ~layer_1[259]; 
    wire [1:0] far_2_2616_0;    relay_conn far_2_2616_0_a(.in(layer_1[751]), .out(far_2_2616_0[0]));    relay_conn far_2_2616_0_b(.in(layer_1[632]), .out(far_2_2616_0[1]));
    wire [1:0] far_2_2616_1;    relay_conn far_2_2616_1_a(.in(far_2_2616_0[0]), .out(far_2_2616_1[0]));    relay_conn far_2_2616_1_b(.in(far_2_2616_0[1]), .out(far_2_2616_1[1]));
    wire [1:0] far_2_2616_2;    relay_conn far_2_2616_2_a(.in(far_2_2616_1[0]), .out(far_2_2616_2[0]));    relay_conn far_2_2616_2_b(.in(far_2_2616_1[1]), .out(far_2_2616_2[1]));
    assign layer_2[576] = far_2_2616_2[1]; 
    wire [1:0] far_2_2617_0;    relay_conn far_2_2617_0_a(.in(layer_1[720]), .out(far_2_2617_0[0]));    relay_conn far_2_2617_0_b(.in(layer_1[799]), .out(far_2_2617_0[1]));
    wire [1:0] far_2_2617_1;    relay_conn far_2_2617_1_a(.in(far_2_2617_0[0]), .out(far_2_2617_1[0]));    relay_conn far_2_2617_1_b(.in(far_2_2617_0[1]), .out(far_2_2617_1[1]));
    assign layer_2[577] = far_2_2617_1[1]; 
    wire [1:0] far_2_2618_0;    relay_conn far_2_2618_0_a(.in(layer_1[284]), .out(far_2_2618_0[0]));    relay_conn far_2_2618_0_b(.in(layer_1[411]), .out(far_2_2618_0[1]));
    wire [1:0] far_2_2618_1;    relay_conn far_2_2618_1_a(.in(far_2_2618_0[0]), .out(far_2_2618_1[0]));    relay_conn far_2_2618_1_b(.in(far_2_2618_0[1]), .out(far_2_2618_1[1]));
    wire [1:0] far_2_2618_2;    relay_conn far_2_2618_2_a(.in(far_2_2618_1[0]), .out(far_2_2618_2[0]));    relay_conn far_2_2618_2_b(.in(far_2_2618_1[1]), .out(far_2_2618_2[1]));
    assign layer_2[578] = ~(far_2_2618_2[0] & far_2_2618_2[1]); 
    wire [1:0] far_2_2619_0;    relay_conn far_2_2619_0_a(.in(layer_1[560]), .out(far_2_2619_0[0]));    relay_conn far_2_2619_0_b(.in(layer_1[603]), .out(far_2_2619_0[1]));
    assign layer_2[579] = far_2_2619_0[0] | far_2_2619_0[1]; 
    assign layer_2[580] = ~(layer_1[566] | layer_1[551]); 
    wire [1:0] far_2_2621_0;    relay_conn far_2_2621_0_a(.in(layer_1[925]), .out(far_2_2621_0[0]));    relay_conn far_2_2621_0_b(.in(layer_1[854]), .out(far_2_2621_0[1]));
    wire [1:0] far_2_2621_1;    relay_conn far_2_2621_1_a(.in(far_2_2621_0[0]), .out(far_2_2621_1[0]));    relay_conn far_2_2621_1_b(.in(far_2_2621_0[1]), .out(far_2_2621_1[1]));
    assign layer_2[581] = far_2_2621_1[0]; 
    wire [1:0] far_2_2622_0;    relay_conn far_2_2622_0_a(.in(layer_1[41]), .out(far_2_2622_0[0]));    relay_conn far_2_2622_0_b(.in(layer_1[134]), .out(far_2_2622_0[1]));
    wire [1:0] far_2_2622_1;    relay_conn far_2_2622_1_a(.in(far_2_2622_0[0]), .out(far_2_2622_1[0]));    relay_conn far_2_2622_1_b(.in(far_2_2622_0[1]), .out(far_2_2622_1[1]));
    assign layer_2[582] = far_2_2622_1[1] & ~far_2_2622_1[0]; 
    assign layer_2[583] = ~layer_1[400] | (layer_1[421] & layer_1[400]); 
    wire [1:0] far_2_2624_0;    relay_conn far_2_2624_0_a(.in(layer_1[482]), .out(far_2_2624_0[0]));    relay_conn far_2_2624_0_b(.in(layer_1[567]), .out(far_2_2624_0[1]));
    wire [1:0] far_2_2624_1;    relay_conn far_2_2624_1_a(.in(far_2_2624_0[0]), .out(far_2_2624_1[0]));    relay_conn far_2_2624_1_b(.in(far_2_2624_0[1]), .out(far_2_2624_1[1]));
    assign layer_2[584] = far_2_2624_1[0] & far_2_2624_1[1]; 
    wire [1:0] far_2_2625_0;    relay_conn far_2_2625_0_a(.in(layer_1[244]), .out(far_2_2625_0[0]));    relay_conn far_2_2625_0_b(.in(layer_1[284]), .out(far_2_2625_0[1]));
    assign layer_2[585] = ~far_2_2625_0[1]; 
    wire [1:0] far_2_2626_0;    relay_conn far_2_2626_0_a(.in(layer_1[340]), .out(far_2_2626_0[0]));    relay_conn far_2_2626_0_b(.in(layer_1[288]), .out(far_2_2626_0[1]));
    assign layer_2[586] = far_2_2626_0[0] | far_2_2626_0[1]; 
    wire [1:0] far_2_2627_0;    relay_conn far_2_2627_0_a(.in(layer_1[264]), .out(far_2_2627_0[0]));    relay_conn far_2_2627_0_b(.in(layer_1[346]), .out(far_2_2627_0[1]));
    wire [1:0] far_2_2627_1;    relay_conn far_2_2627_1_a(.in(far_2_2627_0[0]), .out(far_2_2627_1[0]));    relay_conn far_2_2627_1_b(.in(far_2_2627_0[1]), .out(far_2_2627_1[1]));
    assign layer_2[587] = ~(far_2_2627_1[0] & far_2_2627_1[1]); 
    assign layer_2[588] = ~(layer_1[652] | layer_1[630]); 
    assign layer_2[589] = layer_1[1006] & ~layer_1[1012]; 
    wire [1:0] far_2_2630_0;    relay_conn far_2_2630_0_a(.in(layer_1[619]), .out(far_2_2630_0[0]));    relay_conn far_2_2630_0_b(.in(layer_1[704]), .out(far_2_2630_0[1]));
    wire [1:0] far_2_2630_1;    relay_conn far_2_2630_1_a(.in(far_2_2630_0[0]), .out(far_2_2630_1[0]));    relay_conn far_2_2630_1_b(.in(far_2_2630_0[1]), .out(far_2_2630_1[1]));
    assign layer_2[590] = ~(far_2_2630_1[0] & far_2_2630_1[1]); 
    wire [1:0] far_2_2631_0;    relay_conn far_2_2631_0_a(.in(layer_1[796]), .out(far_2_2631_0[0]));    relay_conn far_2_2631_0_b(.in(layer_1[707]), .out(far_2_2631_0[1]));
    wire [1:0] far_2_2631_1;    relay_conn far_2_2631_1_a(.in(far_2_2631_0[0]), .out(far_2_2631_1[0]));    relay_conn far_2_2631_1_b(.in(far_2_2631_0[1]), .out(far_2_2631_1[1]));
    assign layer_2[591] = ~(far_2_2631_1[0] & far_2_2631_1[1]); 
    assign layer_2[592] = ~layer_1[12] | (layer_1[12] & layer_1[41]); 
    assign layer_2[593] = ~layer_1[850] | (layer_1[838] & layer_1[850]); 
    assign layer_2[594] = ~(layer_1[312] | layer_1[284]); 
    wire [1:0] far_2_2635_0;    relay_conn far_2_2635_0_a(.in(layer_1[159]), .out(far_2_2635_0[0]));    relay_conn far_2_2635_0_b(.in(layer_1[65]), .out(far_2_2635_0[1]));
    wire [1:0] far_2_2635_1;    relay_conn far_2_2635_1_a(.in(far_2_2635_0[0]), .out(far_2_2635_1[0]));    relay_conn far_2_2635_1_b(.in(far_2_2635_0[1]), .out(far_2_2635_1[1]));
    assign layer_2[595] = far_2_2635_1[1] & ~far_2_2635_1[0]; 
    wire [1:0] far_2_2636_0;    relay_conn far_2_2636_0_a(.in(layer_1[645]), .out(far_2_2636_0[0]));    relay_conn far_2_2636_0_b(.in(layer_1[724]), .out(far_2_2636_0[1]));
    wire [1:0] far_2_2636_1;    relay_conn far_2_2636_1_a(.in(far_2_2636_0[0]), .out(far_2_2636_1[0]));    relay_conn far_2_2636_1_b(.in(far_2_2636_0[1]), .out(far_2_2636_1[1]));
    assign layer_2[596] = ~far_2_2636_1[1] | (far_2_2636_1[0] & far_2_2636_1[1]); 
    wire [1:0] far_2_2637_0;    relay_conn far_2_2637_0_a(.in(layer_1[467]), .out(far_2_2637_0[0]));    relay_conn far_2_2637_0_b(.in(layer_1[364]), .out(far_2_2637_0[1]));
    wire [1:0] far_2_2637_1;    relay_conn far_2_2637_1_a(.in(far_2_2637_0[0]), .out(far_2_2637_1[0]));    relay_conn far_2_2637_1_b(.in(far_2_2637_0[1]), .out(far_2_2637_1[1]));
    wire [1:0] far_2_2637_2;    relay_conn far_2_2637_2_a(.in(far_2_2637_1[0]), .out(far_2_2637_2[0]));    relay_conn far_2_2637_2_b(.in(far_2_2637_1[1]), .out(far_2_2637_2[1]));
    assign layer_2[597] = far_2_2637_2[0] & ~far_2_2637_2[1]; 
    wire [1:0] far_2_2638_0;    relay_conn far_2_2638_0_a(.in(layer_1[584]), .out(far_2_2638_0[0]));    relay_conn far_2_2638_0_b(.in(layer_1[702]), .out(far_2_2638_0[1]));
    wire [1:0] far_2_2638_1;    relay_conn far_2_2638_1_a(.in(far_2_2638_0[0]), .out(far_2_2638_1[0]));    relay_conn far_2_2638_1_b(.in(far_2_2638_0[1]), .out(far_2_2638_1[1]));
    wire [1:0] far_2_2638_2;    relay_conn far_2_2638_2_a(.in(far_2_2638_1[0]), .out(far_2_2638_2[0]));    relay_conn far_2_2638_2_b(.in(far_2_2638_1[1]), .out(far_2_2638_2[1]));
    assign layer_2[598] = ~(far_2_2638_2[0] ^ far_2_2638_2[1]); 
    wire [1:0] far_2_2639_0;    relay_conn far_2_2639_0_a(.in(layer_1[841]), .out(far_2_2639_0[0]));    relay_conn far_2_2639_0_b(.in(layer_1[724]), .out(far_2_2639_0[1]));
    wire [1:0] far_2_2639_1;    relay_conn far_2_2639_1_a(.in(far_2_2639_0[0]), .out(far_2_2639_1[0]));    relay_conn far_2_2639_1_b(.in(far_2_2639_0[1]), .out(far_2_2639_1[1]));
    wire [1:0] far_2_2639_2;    relay_conn far_2_2639_2_a(.in(far_2_2639_1[0]), .out(far_2_2639_2[0]));    relay_conn far_2_2639_2_b(.in(far_2_2639_1[1]), .out(far_2_2639_2[1]));
    assign layer_2[599] = far_2_2639_2[0] & ~far_2_2639_2[1]; 
    wire [1:0] far_2_2640_0;    relay_conn far_2_2640_0_a(.in(layer_1[768]), .out(far_2_2640_0[0]));    relay_conn far_2_2640_0_b(.in(layer_1[680]), .out(far_2_2640_0[1]));
    wire [1:0] far_2_2640_1;    relay_conn far_2_2640_1_a(.in(far_2_2640_0[0]), .out(far_2_2640_1[0]));    relay_conn far_2_2640_1_b(.in(far_2_2640_0[1]), .out(far_2_2640_1[1]));
    assign layer_2[600] = ~(far_2_2640_1[0] & far_2_2640_1[1]); 
    wire [1:0] far_2_2641_0;    relay_conn far_2_2641_0_a(.in(layer_1[784]), .out(far_2_2641_0[0]));    relay_conn far_2_2641_0_b(.in(layer_1[702]), .out(far_2_2641_0[1]));
    wire [1:0] far_2_2641_1;    relay_conn far_2_2641_1_a(.in(far_2_2641_0[0]), .out(far_2_2641_1[0]));    relay_conn far_2_2641_1_b(.in(far_2_2641_0[1]), .out(far_2_2641_1[1]));
    assign layer_2[601] = ~far_2_2641_1[0] | (far_2_2641_1[0] & far_2_2641_1[1]); 
    wire [1:0] far_2_2642_0;    relay_conn far_2_2642_0_a(.in(layer_1[200]), .out(far_2_2642_0[0]));    relay_conn far_2_2642_0_b(.in(layer_1[95]), .out(far_2_2642_0[1]));
    wire [1:0] far_2_2642_1;    relay_conn far_2_2642_1_a(.in(far_2_2642_0[0]), .out(far_2_2642_1[0]));    relay_conn far_2_2642_1_b(.in(far_2_2642_0[1]), .out(far_2_2642_1[1]));
    wire [1:0] far_2_2642_2;    relay_conn far_2_2642_2_a(.in(far_2_2642_1[0]), .out(far_2_2642_2[0]));    relay_conn far_2_2642_2_b(.in(far_2_2642_1[1]), .out(far_2_2642_2[1]));
    assign layer_2[602] = ~far_2_2642_2[0]; 
    wire [1:0] far_2_2643_0;    relay_conn far_2_2643_0_a(.in(layer_1[596]), .out(far_2_2643_0[0]));    relay_conn far_2_2643_0_b(.in(layer_1[481]), .out(far_2_2643_0[1]));
    wire [1:0] far_2_2643_1;    relay_conn far_2_2643_1_a(.in(far_2_2643_0[0]), .out(far_2_2643_1[0]));    relay_conn far_2_2643_1_b(.in(far_2_2643_0[1]), .out(far_2_2643_1[1]));
    wire [1:0] far_2_2643_2;    relay_conn far_2_2643_2_a(.in(far_2_2643_1[0]), .out(far_2_2643_2[0]));    relay_conn far_2_2643_2_b(.in(far_2_2643_1[1]), .out(far_2_2643_2[1]));
    assign layer_2[603] = ~(far_2_2643_2[0] & far_2_2643_2[1]); 
    wire [1:0] far_2_2644_0;    relay_conn far_2_2644_0_a(.in(layer_1[647]), .out(far_2_2644_0[0]));    relay_conn far_2_2644_0_b(.in(layer_1[735]), .out(far_2_2644_0[1]));
    wire [1:0] far_2_2644_1;    relay_conn far_2_2644_1_a(.in(far_2_2644_0[0]), .out(far_2_2644_1[0]));    relay_conn far_2_2644_1_b(.in(far_2_2644_0[1]), .out(far_2_2644_1[1]));
    assign layer_2[604] = far_2_2644_1[0] ^ far_2_2644_1[1]; 
    wire [1:0] far_2_2645_0;    relay_conn far_2_2645_0_a(.in(layer_1[559]), .out(far_2_2645_0[0]));    relay_conn far_2_2645_0_b(.in(layer_1[599]), .out(far_2_2645_0[1]));
    assign layer_2[605] = ~(far_2_2645_0[0] ^ far_2_2645_0[1]); 
    wire [1:0] far_2_2646_0;    relay_conn far_2_2646_0_a(.in(layer_1[704]), .out(far_2_2646_0[0]));    relay_conn far_2_2646_0_b(.in(layer_1[603]), .out(far_2_2646_0[1]));
    wire [1:0] far_2_2646_1;    relay_conn far_2_2646_1_a(.in(far_2_2646_0[0]), .out(far_2_2646_1[0]));    relay_conn far_2_2646_1_b(.in(far_2_2646_0[1]), .out(far_2_2646_1[1]));
    wire [1:0] far_2_2646_2;    relay_conn far_2_2646_2_a(.in(far_2_2646_1[0]), .out(far_2_2646_2[0]));    relay_conn far_2_2646_2_b(.in(far_2_2646_1[1]), .out(far_2_2646_2[1]));
    assign layer_2[606] = far_2_2646_2[0] & ~far_2_2646_2[1]; 
    assign layer_2[607] = layer_1[409] & layer_1[397]; 
    wire [1:0] far_2_2648_0;    relay_conn far_2_2648_0_a(.in(layer_1[756]), .out(far_2_2648_0[0]));    relay_conn far_2_2648_0_b(.in(layer_1[685]), .out(far_2_2648_0[1]));
    wire [1:0] far_2_2648_1;    relay_conn far_2_2648_1_a(.in(far_2_2648_0[0]), .out(far_2_2648_1[0]));    relay_conn far_2_2648_1_b(.in(far_2_2648_0[1]), .out(far_2_2648_1[1]));
    assign layer_2[608] = ~(far_2_2648_1[0] | far_2_2648_1[1]); 
    wire [1:0] far_2_2649_0;    relay_conn far_2_2649_0_a(.in(layer_1[947]), .out(far_2_2649_0[0]));    relay_conn far_2_2649_0_b(.in(layer_1[881]), .out(far_2_2649_0[1]));
    wire [1:0] far_2_2649_1;    relay_conn far_2_2649_1_a(.in(far_2_2649_0[0]), .out(far_2_2649_1[0]));    relay_conn far_2_2649_1_b(.in(far_2_2649_0[1]), .out(far_2_2649_1[1]));
    assign layer_2[609] = ~far_2_2649_1[0] | (far_2_2649_1[0] & far_2_2649_1[1]); 
    assign layer_2[610] = ~layer_1[364] | (layer_1[395] & layer_1[364]); 
    wire [1:0] far_2_2651_0;    relay_conn far_2_2651_0_a(.in(layer_1[685]), .out(far_2_2651_0[0]));    relay_conn far_2_2651_0_b(.in(layer_1[742]), .out(far_2_2651_0[1]));
    assign layer_2[611] = ~(far_2_2651_0[0] ^ far_2_2651_0[1]); 
    wire [1:0] far_2_2652_0;    relay_conn far_2_2652_0_a(.in(layer_1[555]), .out(far_2_2652_0[0]));    relay_conn far_2_2652_0_b(.in(layer_1[443]), .out(far_2_2652_0[1]));
    wire [1:0] far_2_2652_1;    relay_conn far_2_2652_1_a(.in(far_2_2652_0[0]), .out(far_2_2652_1[0]));    relay_conn far_2_2652_1_b(.in(far_2_2652_0[1]), .out(far_2_2652_1[1]));
    wire [1:0] far_2_2652_2;    relay_conn far_2_2652_2_a(.in(far_2_2652_1[0]), .out(far_2_2652_2[0]));    relay_conn far_2_2652_2_b(.in(far_2_2652_1[1]), .out(far_2_2652_2[1]));
    assign layer_2[612] = ~(far_2_2652_2[0] | far_2_2652_2[1]); 
    wire [1:0] far_2_2653_0;    relay_conn far_2_2653_0_a(.in(layer_1[276]), .out(far_2_2653_0[0]));    relay_conn far_2_2653_0_b(.in(layer_1[366]), .out(far_2_2653_0[1]));
    wire [1:0] far_2_2653_1;    relay_conn far_2_2653_1_a(.in(far_2_2653_0[0]), .out(far_2_2653_1[0]));    relay_conn far_2_2653_1_b(.in(far_2_2653_0[1]), .out(far_2_2653_1[1]));
    assign layer_2[613] = ~far_2_2653_1[0] | (far_2_2653_1[0] & far_2_2653_1[1]); 
    wire [1:0] far_2_2654_0;    relay_conn far_2_2654_0_a(.in(layer_1[898]), .out(far_2_2654_0[0]));    relay_conn far_2_2654_0_b(.in(layer_1[1001]), .out(far_2_2654_0[1]));
    wire [1:0] far_2_2654_1;    relay_conn far_2_2654_1_a(.in(far_2_2654_0[0]), .out(far_2_2654_1[0]));    relay_conn far_2_2654_1_b(.in(far_2_2654_0[1]), .out(far_2_2654_1[1]));
    wire [1:0] far_2_2654_2;    relay_conn far_2_2654_2_a(.in(far_2_2654_1[0]), .out(far_2_2654_2[0]));    relay_conn far_2_2654_2_b(.in(far_2_2654_1[1]), .out(far_2_2654_2[1]));
    assign layer_2[614] = far_2_2654_2[0] | far_2_2654_2[1]; 
    wire [1:0] far_2_2655_0;    relay_conn far_2_2655_0_a(.in(layer_1[200]), .out(far_2_2655_0[0]));    relay_conn far_2_2655_0_b(.in(layer_1[325]), .out(far_2_2655_0[1]));
    wire [1:0] far_2_2655_1;    relay_conn far_2_2655_1_a(.in(far_2_2655_0[0]), .out(far_2_2655_1[0]));    relay_conn far_2_2655_1_b(.in(far_2_2655_0[1]), .out(far_2_2655_1[1]));
    wire [1:0] far_2_2655_2;    relay_conn far_2_2655_2_a(.in(far_2_2655_1[0]), .out(far_2_2655_2[0]));    relay_conn far_2_2655_2_b(.in(far_2_2655_1[1]), .out(far_2_2655_2[1]));
    assign layer_2[615] = ~far_2_2655_2[0]; 
    wire [1:0] far_2_2656_0;    relay_conn far_2_2656_0_a(.in(layer_1[75]), .out(far_2_2656_0[0]));    relay_conn far_2_2656_0_b(.in(layer_1[139]), .out(far_2_2656_0[1]));
    wire [1:0] far_2_2656_1;    relay_conn far_2_2656_1_a(.in(far_2_2656_0[0]), .out(far_2_2656_1[0]));    relay_conn far_2_2656_1_b(.in(far_2_2656_0[1]), .out(far_2_2656_1[1]));
    assign layer_2[616] = far_2_2656_1[0] | far_2_2656_1[1]; 
    assign layer_2[617] = ~layer_1[533] | (layer_1[508] & layer_1[533]); 
    wire [1:0] far_2_2658_0;    relay_conn far_2_2658_0_a(.in(layer_1[1002]), .out(far_2_2658_0[0]));    relay_conn far_2_2658_0_b(.in(layer_1[879]), .out(far_2_2658_0[1]));
    wire [1:0] far_2_2658_1;    relay_conn far_2_2658_1_a(.in(far_2_2658_0[0]), .out(far_2_2658_1[0]));    relay_conn far_2_2658_1_b(.in(far_2_2658_0[1]), .out(far_2_2658_1[1]));
    wire [1:0] far_2_2658_2;    relay_conn far_2_2658_2_a(.in(far_2_2658_1[0]), .out(far_2_2658_2[0]));    relay_conn far_2_2658_2_b(.in(far_2_2658_1[1]), .out(far_2_2658_2[1]));
    assign layer_2[618] = ~(far_2_2658_2[0] | far_2_2658_2[1]); 
    wire [1:0] far_2_2659_0;    relay_conn far_2_2659_0_a(.in(layer_1[600]), .out(far_2_2659_0[0]));    relay_conn far_2_2659_0_b(.in(layer_1[642]), .out(far_2_2659_0[1]));
    assign layer_2[619] = ~far_2_2659_0[0]; 
    wire [1:0] far_2_2660_0;    relay_conn far_2_2660_0_a(.in(layer_1[146]), .out(far_2_2660_0[0]));    relay_conn far_2_2660_0_b(.in(layer_1[204]), .out(far_2_2660_0[1]));
    assign layer_2[620] = far_2_2660_0[0] & ~far_2_2660_0[1]; 
    wire [1:0] far_2_2661_0;    relay_conn far_2_2661_0_a(.in(layer_1[286]), .out(far_2_2661_0[0]));    relay_conn far_2_2661_0_b(.in(layer_1[183]), .out(far_2_2661_0[1]));
    wire [1:0] far_2_2661_1;    relay_conn far_2_2661_1_a(.in(far_2_2661_0[0]), .out(far_2_2661_1[0]));    relay_conn far_2_2661_1_b(.in(far_2_2661_0[1]), .out(far_2_2661_1[1]));
    wire [1:0] far_2_2661_2;    relay_conn far_2_2661_2_a(.in(far_2_2661_1[0]), .out(far_2_2661_2[0]));    relay_conn far_2_2661_2_b(.in(far_2_2661_1[1]), .out(far_2_2661_2[1]));
    assign layer_2[621] = ~(far_2_2661_2[0] & far_2_2661_2[1]); 
    assign layer_2[622] = layer_1[724] & ~layer_1[701]; 
    wire [1:0] far_2_2663_0;    relay_conn far_2_2663_0_a(.in(layer_1[719]), .out(far_2_2663_0[0]));    relay_conn far_2_2663_0_b(.in(layer_1[761]), .out(far_2_2663_0[1]));
    assign layer_2[623] = ~far_2_2663_0[1] | (far_2_2663_0[0] & far_2_2663_0[1]); 
    wire [1:0] far_2_2664_0;    relay_conn far_2_2664_0_a(.in(layer_1[972]), .out(far_2_2664_0[0]));    relay_conn far_2_2664_0_b(.in(layer_1[882]), .out(far_2_2664_0[1]));
    wire [1:0] far_2_2664_1;    relay_conn far_2_2664_1_a(.in(far_2_2664_0[0]), .out(far_2_2664_1[0]));    relay_conn far_2_2664_1_b(.in(far_2_2664_0[1]), .out(far_2_2664_1[1]));
    assign layer_2[624] = ~(far_2_2664_1[0] & far_2_2664_1[1]); 
    wire [1:0] far_2_2665_0;    relay_conn far_2_2665_0_a(.in(layer_1[587]), .out(far_2_2665_0[0]));    relay_conn far_2_2665_0_b(.in(layer_1[664]), .out(far_2_2665_0[1]));
    wire [1:0] far_2_2665_1;    relay_conn far_2_2665_1_a(.in(far_2_2665_0[0]), .out(far_2_2665_1[0]));    relay_conn far_2_2665_1_b(.in(far_2_2665_0[1]), .out(far_2_2665_1[1]));
    assign layer_2[625] = far_2_2665_1[1]; 
    wire [1:0] far_2_2666_0;    relay_conn far_2_2666_0_a(.in(layer_1[929]), .out(far_2_2666_0[0]));    relay_conn far_2_2666_0_b(.in(layer_1[984]), .out(far_2_2666_0[1]));
    assign layer_2[626] = ~far_2_2666_0[1] | (far_2_2666_0[0] & far_2_2666_0[1]); 
    wire [1:0] far_2_2667_0;    relay_conn far_2_2667_0_a(.in(layer_1[910]), .out(far_2_2667_0[0]));    relay_conn far_2_2667_0_b(.in(layer_1[846]), .out(far_2_2667_0[1]));
    wire [1:0] far_2_2667_1;    relay_conn far_2_2667_1_a(.in(far_2_2667_0[0]), .out(far_2_2667_1[0]));    relay_conn far_2_2667_1_b(.in(far_2_2667_0[1]), .out(far_2_2667_1[1]));
    assign layer_2[627] = far_2_2667_1[0] | far_2_2667_1[1]; 
    wire [1:0] far_2_2668_0;    relay_conn far_2_2668_0_a(.in(layer_1[525]), .out(far_2_2668_0[0]));    relay_conn far_2_2668_0_b(.in(layer_1[436]), .out(far_2_2668_0[1]));
    wire [1:0] far_2_2668_1;    relay_conn far_2_2668_1_a(.in(far_2_2668_0[0]), .out(far_2_2668_1[0]));    relay_conn far_2_2668_1_b(.in(far_2_2668_0[1]), .out(far_2_2668_1[1]));
    assign layer_2[628] = ~(far_2_2668_1[0] | far_2_2668_1[1]); 
    wire [1:0] far_2_2669_0;    relay_conn far_2_2669_0_a(.in(layer_1[566]), .out(far_2_2669_0[0]));    relay_conn far_2_2669_0_b(.in(layer_1[514]), .out(far_2_2669_0[1]));
    assign layer_2[629] = ~far_2_2669_0[0]; 
    assign layer_2[630] = ~layer_1[483] | (layer_1[497] & layer_1[483]); 
    wire [1:0] far_2_2671_0;    relay_conn far_2_2671_0_a(.in(layer_1[656]), .out(far_2_2671_0[0]));    relay_conn far_2_2671_0_b(.in(layer_1[623]), .out(far_2_2671_0[1]));
    assign layer_2[631] = ~(far_2_2671_0[0] | far_2_2671_0[1]); 
    wire [1:0] far_2_2672_0;    relay_conn far_2_2672_0_a(.in(layer_1[12]), .out(far_2_2672_0[0]));    relay_conn far_2_2672_0_b(.in(layer_1[83]), .out(far_2_2672_0[1]));
    wire [1:0] far_2_2672_1;    relay_conn far_2_2672_1_a(.in(far_2_2672_0[0]), .out(far_2_2672_1[0]));    relay_conn far_2_2672_1_b(.in(far_2_2672_0[1]), .out(far_2_2672_1[1]));
    assign layer_2[632] = ~far_2_2672_1[0] | (far_2_2672_1[0] & far_2_2672_1[1]); 
    assign layer_2[633] = layer_1[577] & layer_1[608]; 
    wire [1:0] far_2_2674_0;    relay_conn far_2_2674_0_a(.in(layer_1[559]), .out(far_2_2674_0[0]));    relay_conn far_2_2674_0_b(.in(layer_1[607]), .out(far_2_2674_0[1]));
    assign layer_2[634] = ~(far_2_2674_0[0] & far_2_2674_0[1]); 
    assign layer_2[635] = layer_1[701] & layer_1[705]; 
    wire [1:0] far_2_2676_0;    relay_conn far_2_2676_0_a(.in(layer_1[865]), .out(far_2_2676_0[0]));    relay_conn far_2_2676_0_b(.in(layer_1[962]), .out(far_2_2676_0[1]));
    wire [1:0] far_2_2676_1;    relay_conn far_2_2676_1_a(.in(far_2_2676_0[0]), .out(far_2_2676_1[0]));    relay_conn far_2_2676_1_b(.in(far_2_2676_0[1]), .out(far_2_2676_1[1]));
    wire [1:0] far_2_2676_2;    relay_conn far_2_2676_2_a(.in(far_2_2676_1[0]), .out(far_2_2676_2[0]));    relay_conn far_2_2676_2_b(.in(far_2_2676_1[1]), .out(far_2_2676_2[1]));
    assign layer_2[636] = far_2_2676_2[0]; 
    wire [1:0] far_2_2677_0;    relay_conn far_2_2677_0_a(.in(layer_1[889]), .out(far_2_2677_0[0]));    relay_conn far_2_2677_0_b(.in(layer_1[988]), .out(far_2_2677_0[1]));
    wire [1:0] far_2_2677_1;    relay_conn far_2_2677_1_a(.in(far_2_2677_0[0]), .out(far_2_2677_1[0]));    relay_conn far_2_2677_1_b(.in(far_2_2677_0[1]), .out(far_2_2677_1[1]));
    wire [1:0] far_2_2677_2;    relay_conn far_2_2677_2_a(.in(far_2_2677_1[0]), .out(far_2_2677_2[0]));    relay_conn far_2_2677_2_b(.in(far_2_2677_1[1]), .out(far_2_2677_2[1]));
    assign layer_2[637] = far_2_2677_2[1] & ~far_2_2677_2[0]; 
    wire [1:0] far_2_2678_0;    relay_conn far_2_2678_0_a(.in(layer_1[503]), .out(far_2_2678_0[0]));    relay_conn far_2_2678_0_b(.in(layer_1[423]), .out(far_2_2678_0[1]));
    wire [1:0] far_2_2678_1;    relay_conn far_2_2678_1_a(.in(far_2_2678_0[0]), .out(far_2_2678_1[0]));    relay_conn far_2_2678_1_b(.in(far_2_2678_0[1]), .out(far_2_2678_1[1]));
    assign layer_2[638] = far_2_2678_1[0]; 
    wire [1:0] far_2_2679_0;    relay_conn far_2_2679_0_a(.in(layer_1[867]), .out(far_2_2679_0[0]));    relay_conn far_2_2679_0_b(.in(layer_1[822]), .out(far_2_2679_0[1]));
    assign layer_2[639] = ~far_2_2679_0[0] | (far_2_2679_0[0] & far_2_2679_0[1]); 
    wire [1:0] far_2_2680_0;    relay_conn far_2_2680_0_a(.in(layer_1[1008]), .out(far_2_2680_0[0]));    relay_conn far_2_2680_0_b(.in(layer_1[941]), .out(far_2_2680_0[1]));
    wire [1:0] far_2_2680_1;    relay_conn far_2_2680_1_a(.in(far_2_2680_0[0]), .out(far_2_2680_1[0]));    relay_conn far_2_2680_1_b(.in(far_2_2680_0[1]), .out(far_2_2680_1[1]));
    assign layer_2[640] = ~far_2_2680_1[0] | (far_2_2680_1[0] & far_2_2680_1[1]); 
    assign layer_2[641] = ~(layer_1[102] ^ layer_1[115]); 
    wire [1:0] far_2_2682_0;    relay_conn far_2_2682_0_a(.in(layer_1[267]), .out(far_2_2682_0[0]));    relay_conn far_2_2682_0_b(.in(layer_1[140]), .out(far_2_2682_0[1]));
    wire [1:0] far_2_2682_1;    relay_conn far_2_2682_1_a(.in(far_2_2682_0[0]), .out(far_2_2682_1[0]));    relay_conn far_2_2682_1_b(.in(far_2_2682_0[1]), .out(far_2_2682_1[1]));
    wire [1:0] far_2_2682_2;    relay_conn far_2_2682_2_a(.in(far_2_2682_1[0]), .out(far_2_2682_2[0]));    relay_conn far_2_2682_2_b(.in(far_2_2682_1[1]), .out(far_2_2682_2[1]));
    assign layer_2[642] = far_2_2682_2[0] ^ far_2_2682_2[1]; 
    wire [1:0] far_2_2683_0;    relay_conn far_2_2683_0_a(.in(layer_1[280]), .out(far_2_2683_0[0]));    relay_conn far_2_2683_0_b(.in(layer_1[322]), .out(far_2_2683_0[1]));
    assign layer_2[643] = ~far_2_2683_0[1]; 
    wire [1:0] far_2_2684_0;    relay_conn far_2_2684_0_a(.in(layer_1[409]), .out(far_2_2684_0[0]));    relay_conn far_2_2684_0_b(.in(layer_1[313]), .out(far_2_2684_0[1]));
    wire [1:0] far_2_2684_1;    relay_conn far_2_2684_1_a(.in(far_2_2684_0[0]), .out(far_2_2684_1[0]));    relay_conn far_2_2684_1_b(.in(far_2_2684_0[1]), .out(far_2_2684_1[1]));
    wire [1:0] far_2_2684_2;    relay_conn far_2_2684_2_a(.in(far_2_2684_1[0]), .out(far_2_2684_2[0]));    relay_conn far_2_2684_2_b(.in(far_2_2684_1[1]), .out(far_2_2684_2[1]));
    assign layer_2[644] = far_2_2684_2[0] & far_2_2684_2[1]; 
    assign layer_2[645] = layer_1[642] | layer_1[619]; 
    wire [1:0] far_2_2686_0;    relay_conn far_2_2686_0_a(.in(layer_1[815]), .out(far_2_2686_0[0]));    relay_conn far_2_2686_0_b(.in(layer_1[721]), .out(far_2_2686_0[1]));
    wire [1:0] far_2_2686_1;    relay_conn far_2_2686_1_a(.in(far_2_2686_0[0]), .out(far_2_2686_1[0]));    relay_conn far_2_2686_1_b(.in(far_2_2686_0[1]), .out(far_2_2686_1[1]));
    assign layer_2[646] = ~far_2_2686_1[1]; 
    wire [1:0] far_2_2687_0;    relay_conn far_2_2687_0_a(.in(layer_1[22]), .out(far_2_2687_0[0]));    relay_conn far_2_2687_0_b(.in(layer_1[133]), .out(far_2_2687_0[1]));
    wire [1:0] far_2_2687_1;    relay_conn far_2_2687_1_a(.in(far_2_2687_0[0]), .out(far_2_2687_1[0]));    relay_conn far_2_2687_1_b(.in(far_2_2687_0[1]), .out(far_2_2687_1[1]));
    wire [1:0] far_2_2687_2;    relay_conn far_2_2687_2_a(.in(far_2_2687_1[0]), .out(far_2_2687_2[0]));    relay_conn far_2_2687_2_b(.in(far_2_2687_1[1]), .out(far_2_2687_2[1]));
    assign layer_2[647] = far_2_2687_2[0] & ~far_2_2687_2[1]; 
    wire [1:0] far_2_2688_0;    relay_conn far_2_2688_0_a(.in(layer_1[241]), .out(far_2_2688_0[0]));    relay_conn far_2_2688_0_b(.in(layer_1[319]), .out(far_2_2688_0[1]));
    wire [1:0] far_2_2688_1;    relay_conn far_2_2688_1_a(.in(far_2_2688_0[0]), .out(far_2_2688_1[0]));    relay_conn far_2_2688_1_b(.in(far_2_2688_0[1]), .out(far_2_2688_1[1]));
    assign layer_2[648] = ~far_2_2688_1[1]; 
    assign layer_2[649] = ~(layer_1[722] | layer_1[710]); 
    wire [1:0] far_2_2690_0;    relay_conn far_2_2690_0_a(.in(layer_1[446]), .out(far_2_2690_0[0]));    relay_conn far_2_2690_0_b(.in(layer_1[491]), .out(far_2_2690_0[1]));
    assign layer_2[650] = ~(far_2_2690_0[0] & far_2_2690_0[1]); 
    assign layer_2[651] = ~(layer_1[690] | layer_1[715]); 
    assign layer_2[652] = layer_1[204] & ~layer_1[231]; 
    wire [1:0] far_2_2693_0;    relay_conn far_2_2693_0_a(.in(layer_1[299]), .out(far_2_2693_0[0]));    relay_conn far_2_2693_0_b(.in(layer_1[241]), .out(far_2_2693_0[1]));
    assign layer_2[653] = far_2_2693_0[0] & ~far_2_2693_0[1]; 
    wire [1:0] far_2_2694_0;    relay_conn far_2_2694_0_a(.in(layer_1[348]), .out(far_2_2694_0[0]));    relay_conn far_2_2694_0_b(.in(layer_1[288]), .out(far_2_2694_0[1]));
    assign layer_2[654] = ~far_2_2694_0[0] | (far_2_2694_0[0] & far_2_2694_0[1]); 
    wire [1:0] far_2_2695_0;    relay_conn far_2_2695_0_a(.in(layer_1[95]), .out(far_2_2695_0[0]));    relay_conn far_2_2695_0_b(.in(layer_1[55]), .out(far_2_2695_0[1]));
    assign layer_2[655] = ~far_2_2695_0[0] | (far_2_2695_0[0] & far_2_2695_0[1]); 
    wire [1:0] far_2_2696_0;    relay_conn far_2_2696_0_a(.in(layer_1[676]), .out(far_2_2696_0[0]));    relay_conn far_2_2696_0_b(.in(layer_1[553]), .out(far_2_2696_0[1]));
    wire [1:0] far_2_2696_1;    relay_conn far_2_2696_1_a(.in(far_2_2696_0[0]), .out(far_2_2696_1[0]));    relay_conn far_2_2696_1_b(.in(far_2_2696_0[1]), .out(far_2_2696_1[1]));
    wire [1:0] far_2_2696_2;    relay_conn far_2_2696_2_a(.in(far_2_2696_1[0]), .out(far_2_2696_2[0]));    relay_conn far_2_2696_2_b(.in(far_2_2696_1[1]), .out(far_2_2696_2[1]));
    assign layer_2[656] = far_2_2696_2[0] & ~far_2_2696_2[1]; 
    wire [1:0] far_2_2697_0;    relay_conn far_2_2697_0_a(.in(layer_1[390]), .out(far_2_2697_0[0]));    relay_conn far_2_2697_0_b(.in(layer_1[309]), .out(far_2_2697_0[1]));
    wire [1:0] far_2_2697_1;    relay_conn far_2_2697_1_a(.in(far_2_2697_0[0]), .out(far_2_2697_1[0]));    relay_conn far_2_2697_1_b(.in(far_2_2697_0[1]), .out(far_2_2697_1[1]));
    assign layer_2[657] = far_2_2697_1[0] | far_2_2697_1[1]; 
    wire [1:0] far_2_2698_0;    relay_conn far_2_2698_0_a(.in(layer_1[312]), .out(far_2_2698_0[0]));    relay_conn far_2_2698_0_b(.in(layer_1[189]), .out(far_2_2698_0[1]));
    wire [1:0] far_2_2698_1;    relay_conn far_2_2698_1_a(.in(far_2_2698_0[0]), .out(far_2_2698_1[0]));    relay_conn far_2_2698_1_b(.in(far_2_2698_0[1]), .out(far_2_2698_1[1]));
    wire [1:0] far_2_2698_2;    relay_conn far_2_2698_2_a(.in(far_2_2698_1[0]), .out(far_2_2698_2[0]));    relay_conn far_2_2698_2_b(.in(far_2_2698_1[1]), .out(far_2_2698_2[1]));
    assign layer_2[658] = ~far_2_2698_2[1]; 
    assign layer_2[659] = layer_1[280] | layer_1[284]; 
    wire [1:0] far_2_2700_0;    relay_conn far_2_2700_0_a(.in(layer_1[910]), .out(far_2_2700_0[0]));    relay_conn far_2_2700_0_b(.in(layer_1[871]), .out(far_2_2700_0[1]));
    assign layer_2[660] = far_2_2700_0[0] & far_2_2700_0[1]; 
    wire [1:0] far_2_2701_0;    relay_conn far_2_2701_0_a(.in(layer_1[520]), .out(far_2_2701_0[0]));    relay_conn far_2_2701_0_b(.in(layer_1[559]), .out(far_2_2701_0[1]));
    assign layer_2[661] = ~(far_2_2701_0[0] & far_2_2701_0[1]); 
    wire [1:0] far_2_2702_0;    relay_conn far_2_2702_0_a(.in(layer_1[596]), .out(far_2_2702_0[0]));    relay_conn far_2_2702_0_b(.in(layer_1[528]), .out(far_2_2702_0[1]));
    wire [1:0] far_2_2702_1;    relay_conn far_2_2702_1_a(.in(far_2_2702_0[0]), .out(far_2_2702_1[0]));    relay_conn far_2_2702_1_b(.in(far_2_2702_0[1]), .out(far_2_2702_1[1]));
    assign layer_2[662] = far_2_2702_1[1] & ~far_2_2702_1[0]; 
    wire [1:0] far_2_2703_0;    relay_conn far_2_2703_0_a(.in(layer_1[882]), .out(far_2_2703_0[0]));    relay_conn far_2_2703_0_b(.in(layer_1[776]), .out(far_2_2703_0[1]));
    wire [1:0] far_2_2703_1;    relay_conn far_2_2703_1_a(.in(far_2_2703_0[0]), .out(far_2_2703_1[0]));    relay_conn far_2_2703_1_b(.in(far_2_2703_0[1]), .out(far_2_2703_1[1]));
    wire [1:0] far_2_2703_2;    relay_conn far_2_2703_2_a(.in(far_2_2703_1[0]), .out(far_2_2703_2[0]));    relay_conn far_2_2703_2_b(.in(far_2_2703_1[1]), .out(far_2_2703_2[1]));
    assign layer_2[663] = far_2_2703_2[0] & ~far_2_2703_2[1]; 
    assign layer_2[664] = ~(layer_1[404] & layer_1[426]); 
    wire [1:0] far_2_2705_0;    relay_conn far_2_2705_0_a(.in(layer_1[352]), .out(far_2_2705_0[0]));    relay_conn far_2_2705_0_b(.in(layer_1[258]), .out(far_2_2705_0[1]));
    wire [1:0] far_2_2705_1;    relay_conn far_2_2705_1_a(.in(far_2_2705_0[0]), .out(far_2_2705_1[0]));    relay_conn far_2_2705_1_b(.in(far_2_2705_0[1]), .out(far_2_2705_1[1]));
    assign layer_2[665] = far_2_2705_1[0]; 
    wire [1:0] far_2_2706_0;    relay_conn far_2_2706_0_a(.in(layer_1[207]), .out(far_2_2706_0[0]));    relay_conn far_2_2706_0_b(.in(layer_1[329]), .out(far_2_2706_0[1]));
    wire [1:0] far_2_2706_1;    relay_conn far_2_2706_1_a(.in(far_2_2706_0[0]), .out(far_2_2706_1[0]));    relay_conn far_2_2706_1_b(.in(far_2_2706_0[1]), .out(far_2_2706_1[1]));
    wire [1:0] far_2_2706_2;    relay_conn far_2_2706_2_a(.in(far_2_2706_1[0]), .out(far_2_2706_2[0]));    relay_conn far_2_2706_2_b(.in(far_2_2706_1[1]), .out(far_2_2706_2[1]));
    assign layer_2[666] = ~(far_2_2706_2[0] | far_2_2706_2[1]); 
    wire [1:0] far_2_2707_0;    relay_conn far_2_2707_0_a(.in(layer_1[763]), .out(far_2_2707_0[0]));    relay_conn far_2_2707_0_b(.in(layer_1[875]), .out(far_2_2707_0[1]));
    wire [1:0] far_2_2707_1;    relay_conn far_2_2707_1_a(.in(far_2_2707_0[0]), .out(far_2_2707_1[0]));    relay_conn far_2_2707_1_b(.in(far_2_2707_0[1]), .out(far_2_2707_1[1]));
    wire [1:0] far_2_2707_2;    relay_conn far_2_2707_2_a(.in(far_2_2707_1[0]), .out(far_2_2707_2[0]));    relay_conn far_2_2707_2_b(.in(far_2_2707_1[1]), .out(far_2_2707_2[1]));
    assign layer_2[667] = ~far_2_2707_2[1]; 
    assign layer_2[668] = layer_1[21] ^ layer_1[11]; 
    wire [1:0] far_2_2709_0;    relay_conn far_2_2709_0_a(.in(layer_1[984]), .out(far_2_2709_0[0]));    relay_conn far_2_2709_0_b(.in(layer_1[888]), .out(far_2_2709_0[1]));
    wire [1:0] far_2_2709_1;    relay_conn far_2_2709_1_a(.in(far_2_2709_0[0]), .out(far_2_2709_1[0]));    relay_conn far_2_2709_1_b(.in(far_2_2709_0[1]), .out(far_2_2709_1[1]));
    wire [1:0] far_2_2709_2;    relay_conn far_2_2709_2_a(.in(far_2_2709_1[0]), .out(far_2_2709_2[0]));    relay_conn far_2_2709_2_b(.in(far_2_2709_1[1]), .out(far_2_2709_2[1]));
    assign layer_2[669] = ~far_2_2709_2[0] | (far_2_2709_2[0] & far_2_2709_2[1]); 
    wire [1:0] far_2_2710_0;    relay_conn far_2_2710_0_a(.in(layer_1[952]), .out(far_2_2710_0[0]));    relay_conn far_2_2710_0_b(.in(layer_1[867]), .out(far_2_2710_0[1]));
    wire [1:0] far_2_2710_1;    relay_conn far_2_2710_1_a(.in(far_2_2710_0[0]), .out(far_2_2710_1[0]));    relay_conn far_2_2710_1_b(.in(far_2_2710_0[1]), .out(far_2_2710_1[1]));
    assign layer_2[670] = far_2_2710_1[0] & ~far_2_2710_1[1]; 
    assign layer_2[671] = layer_1[780] & ~layer_1[810]; 
    assign layer_2[672] = layer_1[176]; 
    wire [1:0] far_2_2713_0;    relay_conn far_2_2713_0_a(.in(layer_1[289]), .out(far_2_2713_0[0]));    relay_conn far_2_2713_0_b(.in(layer_1[358]), .out(far_2_2713_0[1]));
    wire [1:0] far_2_2713_1;    relay_conn far_2_2713_1_a(.in(far_2_2713_0[0]), .out(far_2_2713_1[0]));    relay_conn far_2_2713_1_b(.in(far_2_2713_0[1]), .out(far_2_2713_1[1]));
    assign layer_2[673] = ~(far_2_2713_1[0] | far_2_2713_1[1]); 
    wire [1:0] far_2_2714_0;    relay_conn far_2_2714_0_a(.in(layer_1[569]), .out(far_2_2714_0[0]));    relay_conn far_2_2714_0_b(.in(layer_1[647]), .out(far_2_2714_0[1]));
    wire [1:0] far_2_2714_1;    relay_conn far_2_2714_1_a(.in(far_2_2714_0[0]), .out(far_2_2714_1[0]));    relay_conn far_2_2714_1_b(.in(far_2_2714_0[1]), .out(far_2_2714_1[1]));
    assign layer_2[674] = far_2_2714_1[0] & far_2_2714_1[1]; 
    wire [1:0] far_2_2715_0;    relay_conn far_2_2715_0_a(.in(layer_1[521]), .out(far_2_2715_0[0]));    relay_conn far_2_2715_0_b(.in(layer_1[439]), .out(far_2_2715_0[1]));
    wire [1:0] far_2_2715_1;    relay_conn far_2_2715_1_a(.in(far_2_2715_0[0]), .out(far_2_2715_1[0]));    relay_conn far_2_2715_1_b(.in(far_2_2715_0[1]), .out(far_2_2715_1[1]));
    assign layer_2[675] = far_2_2715_1[0] | far_2_2715_1[1]; 
    wire [1:0] far_2_2716_0;    relay_conn far_2_2716_0_a(.in(layer_1[174]), .out(far_2_2716_0[0]));    relay_conn far_2_2716_0_b(.in(layer_1[240]), .out(far_2_2716_0[1]));
    wire [1:0] far_2_2716_1;    relay_conn far_2_2716_1_a(.in(far_2_2716_0[0]), .out(far_2_2716_1[0]));    relay_conn far_2_2716_1_b(.in(far_2_2716_0[1]), .out(far_2_2716_1[1]));
    assign layer_2[676] = far_2_2716_1[1]; 
    assign layer_2[677] = layer_1[837] & ~layer_1[836]; 
    wire [1:0] far_2_2718_0;    relay_conn far_2_2718_0_a(.in(layer_1[747]), .out(far_2_2718_0[0]));    relay_conn far_2_2718_0_b(.in(layer_1[619]), .out(far_2_2718_0[1]));
    wire [1:0] far_2_2718_1;    relay_conn far_2_2718_1_a(.in(far_2_2718_0[0]), .out(far_2_2718_1[0]));    relay_conn far_2_2718_1_b(.in(far_2_2718_0[1]), .out(far_2_2718_1[1]));
    wire [1:0] far_2_2718_2;    relay_conn far_2_2718_2_a(.in(far_2_2718_1[0]), .out(far_2_2718_2[0]));    relay_conn far_2_2718_2_b(.in(far_2_2718_1[1]), .out(far_2_2718_2[1]));
    wire [1:0] far_2_2718_3;    relay_conn far_2_2718_3_a(.in(far_2_2718_2[0]), .out(far_2_2718_3[0]));    relay_conn far_2_2718_3_b(.in(far_2_2718_2[1]), .out(far_2_2718_3[1]));
    assign layer_2[678] = ~far_2_2718_3[0] | (far_2_2718_3[0] & far_2_2718_3[1]); 
    wire [1:0] far_2_2719_0;    relay_conn far_2_2719_0_a(.in(layer_1[532]), .out(far_2_2719_0[0]));    relay_conn far_2_2719_0_b(.in(layer_1[419]), .out(far_2_2719_0[1]));
    wire [1:0] far_2_2719_1;    relay_conn far_2_2719_1_a(.in(far_2_2719_0[0]), .out(far_2_2719_1[0]));    relay_conn far_2_2719_1_b(.in(far_2_2719_0[1]), .out(far_2_2719_1[1]));
    wire [1:0] far_2_2719_2;    relay_conn far_2_2719_2_a(.in(far_2_2719_1[0]), .out(far_2_2719_2[0]));    relay_conn far_2_2719_2_b(.in(far_2_2719_1[1]), .out(far_2_2719_2[1]));
    assign layer_2[679] = far_2_2719_2[1] & ~far_2_2719_2[0]; 
    assign layer_2[680] = layer_1[40] | layer_1[32]; 
    assign layer_2[681] = ~layer_1[248]; 
    wire [1:0] far_2_2722_0;    relay_conn far_2_2722_0_a(.in(layer_1[646]), .out(far_2_2722_0[0]));    relay_conn far_2_2722_0_b(.in(layer_1[743]), .out(far_2_2722_0[1]));
    wire [1:0] far_2_2722_1;    relay_conn far_2_2722_1_a(.in(far_2_2722_0[0]), .out(far_2_2722_1[0]));    relay_conn far_2_2722_1_b(.in(far_2_2722_0[1]), .out(far_2_2722_1[1]));
    wire [1:0] far_2_2722_2;    relay_conn far_2_2722_2_a(.in(far_2_2722_1[0]), .out(far_2_2722_2[0]));    relay_conn far_2_2722_2_b(.in(far_2_2722_1[1]), .out(far_2_2722_2[1]));
    assign layer_2[682] = ~(far_2_2722_2[0] & far_2_2722_2[1]); 
    wire [1:0] far_2_2723_0;    relay_conn far_2_2723_0_a(.in(layer_1[517]), .out(far_2_2723_0[0]));    relay_conn far_2_2723_0_b(.in(layer_1[428]), .out(far_2_2723_0[1]));
    wire [1:0] far_2_2723_1;    relay_conn far_2_2723_1_a(.in(far_2_2723_0[0]), .out(far_2_2723_1[0]));    relay_conn far_2_2723_1_b(.in(far_2_2723_0[1]), .out(far_2_2723_1[1]));
    assign layer_2[683] = ~far_2_2723_1[1]; 
    wire [1:0] far_2_2724_0;    relay_conn far_2_2724_0_a(.in(layer_1[927]), .out(far_2_2724_0[0]));    relay_conn far_2_2724_0_b(.in(layer_1[825]), .out(far_2_2724_0[1]));
    wire [1:0] far_2_2724_1;    relay_conn far_2_2724_1_a(.in(far_2_2724_0[0]), .out(far_2_2724_1[0]));    relay_conn far_2_2724_1_b(.in(far_2_2724_0[1]), .out(far_2_2724_1[1]));
    wire [1:0] far_2_2724_2;    relay_conn far_2_2724_2_a(.in(far_2_2724_1[0]), .out(far_2_2724_2[0]));    relay_conn far_2_2724_2_b(.in(far_2_2724_1[1]), .out(far_2_2724_2[1]));
    assign layer_2[684] = ~far_2_2724_2[0]; 
    wire [1:0] far_2_2725_0;    relay_conn far_2_2725_0_a(.in(layer_1[833]), .out(far_2_2725_0[0]));    relay_conn far_2_2725_0_b(.in(layer_1[727]), .out(far_2_2725_0[1]));
    wire [1:0] far_2_2725_1;    relay_conn far_2_2725_1_a(.in(far_2_2725_0[0]), .out(far_2_2725_1[0]));    relay_conn far_2_2725_1_b(.in(far_2_2725_0[1]), .out(far_2_2725_1[1]));
    wire [1:0] far_2_2725_2;    relay_conn far_2_2725_2_a(.in(far_2_2725_1[0]), .out(far_2_2725_2[0]));    relay_conn far_2_2725_2_b(.in(far_2_2725_1[1]), .out(far_2_2725_2[1]));
    assign layer_2[685] = far_2_2725_2[1]; 
    wire [1:0] far_2_2726_0;    relay_conn far_2_2726_0_a(.in(layer_1[768]), .out(far_2_2726_0[0]));    relay_conn far_2_2726_0_b(.in(layer_1[855]), .out(far_2_2726_0[1]));
    wire [1:0] far_2_2726_1;    relay_conn far_2_2726_1_a(.in(far_2_2726_0[0]), .out(far_2_2726_1[0]));    relay_conn far_2_2726_1_b(.in(far_2_2726_0[1]), .out(far_2_2726_1[1]));
    assign layer_2[686] = ~far_2_2726_1[0]; 
    wire [1:0] far_2_2727_0;    relay_conn far_2_2727_0_a(.in(layer_1[352]), .out(far_2_2727_0[0]));    relay_conn far_2_2727_0_b(.in(layer_1[419]), .out(far_2_2727_0[1]));
    wire [1:0] far_2_2727_1;    relay_conn far_2_2727_1_a(.in(far_2_2727_0[0]), .out(far_2_2727_1[0]));    relay_conn far_2_2727_1_b(.in(far_2_2727_0[1]), .out(far_2_2727_1[1]));
    assign layer_2[687] = ~far_2_2727_1[0] | (far_2_2727_1[0] & far_2_2727_1[1]); 
    wire [1:0] far_2_2728_0;    relay_conn far_2_2728_0_a(.in(layer_1[867]), .out(far_2_2728_0[0]));    relay_conn far_2_2728_0_b(.in(layer_1[767]), .out(far_2_2728_0[1]));
    wire [1:0] far_2_2728_1;    relay_conn far_2_2728_1_a(.in(far_2_2728_0[0]), .out(far_2_2728_1[0]));    relay_conn far_2_2728_1_b(.in(far_2_2728_0[1]), .out(far_2_2728_1[1]));
    wire [1:0] far_2_2728_2;    relay_conn far_2_2728_2_a(.in(far_2_2728_1[0]), .out(far_2_2728_2[0]));    relay_conn far_2_2728_2_b(.in(far_2_2728_1[1]), .out(far_2_2728_2[1]));
    assign layer_2[688] = far_2_2728_2[0] & far_2_2728_2[1]; 
    wire [1:0] far_2_2729_0;    relay_conn far_2_2729_0_a(.in(layer_1[630]), .out(far_2_2729_0[0]));    relay_conn far_2_2729_0_b(.in(layer_1[558]), .out(far_2_2729_0[1]));
    wire [1:0] far_2_2729_1;    relay_conn far_2_2729_1_a(.in(far_2_2729_0[0]), .out(far_2_2729_1[0]));    relay_conn far_2_2729_1_b(.in(far_2_2729_0[1]), .out(far_2_2729_1[1]));
    assign layer_2[689] = far_2_2729_1[0] & ~far_2_2729_1[1]; 
    wire [1:0] far_2_2730_0;    relay_conn far_2_2730_0_a(.in(layer_1[855]), .out(far_2_2730_0[0]));    relay_conn far_2_2730_0_b(.in(layer_1[977]), .out(far_2_2730_0[1]));
    wire [1:0] far_2_2730_1;    relay_conn far_2_2730_1_a(.in(far_2_2730_0[0]), .out(far_2_2730_1[0]));    relay_conn far_2_2730_1_b(.in(far_2_2730_0[1]), .out(far_2_2730_1[1]));
    wire [1:0] far_2_2730_2;    relay_conn far_2_2730_2_a(.in(far_2_2730_1[0]), .out(far_2_2730_2[0]));    relay_conn far_2_2730_2_b(.in(far_2_2730_1[1]), .out(far_2_2730_2[1]));
    assign layer_2[690] = ~(far_2_2730_2[0] | far_2_2730_2[1]); 
    wire [1:0] far_2_2731_0;    relay_conn far_2_2731_0_a(.in(layer_1[557]), .out(far_2_2731_0[0]));    relay_conn far_2_2731_0_b(.in(layer_1[597]), .out(far_2_2731_0[1]));
    assign layer_2[691] = ~(far_2_2731_0[0] & far_2_2731_0[1]); 
    assign layer_2[692] = ~(layer_1[833] ^ layer_1[838]); 
    wire [1:0] far_2_2733_0;    relay_conn far_2_2733_0_a(.in(layer_1[57]), .out(far_2_2733_0[0]));    relay_conn far_2_2733_0_b(.in(layer_1[184]), .out(far_2_2733_0[1]));
    wire [1:0] far_2_2733_1;    relay_conn far_2_2733_1_a(.in(far_2_2733_0[0]), .out(far_2_2733_1[0]));    relay_conn far_2_2733_1_b(.in(far_2_2733_0[1]), .out(far_2_2733_1[1]));
    wire [1:0] far_2_2733_2;    relay_conn far_2_2733_2_a(.in(far_2_2733_1[0]), .out(far_2_2733_2[0]));    relay_conn far_2_2733_2_b(.in(far_2_2733_1[1]), .out(far_2_2733_2[1]));
    assign layer_2[693] = far_2_2733_2[0] | far_2_2733_2[1]; 
    wire [1:0] far_2_2734_0;    relay_conn far_2_2734_0_a(.in(layer_1[419]), .out(far_2_2734_0[0]));    relay_conn far_2_2734_0_b(.in(layer_1[455]), .out(far_2_2734_0[1]));
    assign layer_2[694] = ~far_2_2734_0[0] | (far_2_2734_0[0] & far_2_2734_0[1]); 
    assign layer_2[695] = layer_1[558] & layer_1[547]; 
    wire [1:0] far_2_2736_0;    relay_conn far_2_2736_0_a(.in(layer_1[469]), .out(far_2_2736_0[0]));    relay_conn far_2_2736_0_b(.in(layer_1[514]), .out(far_2_2736_0[1]));
    assign layer_2[696] = ~(far_2_2736_0[0] & far_2_2736_0[1]); 
    assign layer_2[697] = layer_1[959]; 
    wire [1:0] far_2_2738_0;    relay_conn far_2_2738_0_a(.in(layer_1[513]), .out(far_2_2738_0[0]));    relay_conn far_2_2738_0_b(.in(layer_1[562]), .out(far_2_2738_0[1]));
    assign layer_2[698] = ~far_2_2738_0[0]; 
    wire [1:0] far_2_2739_0;    relay_conn far_2_2739_0_a(.in(layer_1[795]), .out(far_2_2739_0[0]));    relay_conn far_2_2739_0_b(.in(layer_1[864]), .out(far_2_2739_0[1]));
    wire [1:0] far_2_2739_1;    relay_conn far_2_2739_1_a(.in(far_2_2739_0[0]), .out(far_2_2739_1[0]));    relay_conn far_2_2739_1_b(.in(far_2_2739_0[1]), .out(far_2_2739_1[1]));
    assign layer_2[699] = ~(far_2_2739_1[0] ^ far_2_2739_1[1]); 
    wire [1:0] far_2_2740_0;    relay_conn far_2_2740_0_a(.in(layer_1[1008]), .out(far_2_2740_0[0]));    relay_conn far_2_2740_0_b(.in(layer_1[949]), .out(far_2_2740_0[1]));
    assign layer_2[700] = ~far_2_2740_0[1] | (far_2_2740_0[0] & far_2_2740_0[1]); 
    wire [1:0] far_2_2741_0;    relay_conn far_2_2741_0_a(.in(layer_1[248]), .out(far_2_2741_0[0]));    relay_conn far_2_2741_0_b(.in(layer_1[188]), .out(far_2_2741_0[1]));
    assign layer_2[701] = ~far_2_2741_0[0] | (far_2_2741_0[0] & far_2_2741_0[1]); 
    assign layer_2[702] = ~layer_1[949] | (layer_1[949] & layer_1[962]); 
    wire [1:0] far_2_2743_0;    relay_conn far_2_2743_0_a(.in(layer_1[548]), .out(far_2_2743_0[0]));    relay_conn far_2_2743_0_b(.in(layer_1[474]), .out(far_2_2743_0[1]));
    wire [1:0] far_2_2743_1;    relay_conn far_2_2743_1_a(.in(far_2_2743_0[0]), .out(far_2_2743_1[0]));    relay_conn far_2_2743_1_b(.in(far_2_2743_0[1]), .out(far_2_2743_1[1]));
    assign layer_2[703] = ~(far_2_2743_1[0] | far_2_2743_1[1]); 
    wire [1:0] far_2_2744_0;    relay_conn far_2_2744_0_a(.in(layer_1[851]), .out(far_2_2744_0[0]));    relay_conn far_2_2744_0_b(.in(layer_1[783]), .out(far_2_2744_0[1]));
    wire [1:0] far_2_2744_1;    relay_conn far_2_2744_1_a(.in(far_2_2744_0[0]), .out(far_2_2744_1[0]));    relay_conn far_2_2744_1_b(.in(far_2_2744_0[1]), .out(far_2_2744_1[1]));
    assign layer_2[704] = far_2_2744_1[0] ^ far_2_2744_1[1]; 
    wire [1:0] far_2_2745_0;    relay_conn far_2_2745_0_a(.in(layer_1[188]), .out(far_2_2745_0[0]));    relay_conn far_2_2745_0_b(.in(layer_1[261]), .out(far_2_2745_0[1]));
    wire [1:0] far_2_2745_1;    relay_conn far_2_2745_1_a(.in(far_2_2745_0[0]), .out(far_2_2745_1[0]));    relay_conn far_2_2745_1_b(.in(far_2_2745_0[1]), .out(far_2_2745_1[1]));
    assign layer_2[705] = ~far_2_2745_1[0]; 
    wire [1:0] far_2_2746_0;    relay_conn far_2_2746_0_a(.in(layer_1[169]), .out(far_2_2746_0[0]));    relay_conn far_2_2746_0_b(.in(layer_1[75]), .out(far_2_2746_0[1]));
    wire [1:0] far_2_2746_1;    relay_conn far_2_2746_1_a(.in(far_2_2746_0[0]), .out(far_2_2746_1[0]));    relay_conn far_2_2746_1_b(.in(far_2_2746_0[1]), .out(far_2_2746_1[1]));
    assign layer_2[706] = ~far_2_2746_1[0] | (far_2_2746_1[0] & far_2_2746_1[1]); 
    wire [1:0] far_2_2747_0;    relay_conn far_2_2747_0_a(.in(layer_1[563]), .out(far_2_2747_0[0]));    relay_conn far_2_2747_0_b(.in(layer_1[518]), .out(far_2_2747_0[1]));
    assign layer_2[707] = ~(far_2_2747_0[0] | far_2_2747_0[1]); 
    wire [1:0] far_2_2748_0;    relay_conn far_2_2748_0_a(.in(layer_1[248]), .out(far_2_2748_0[0]));    relay_conn far_2_2748_0_b(.in(layer_1[135]), .out(far_2_2748_0[1]));
    wire [1:0] far_2_2748_1;    relay_conn far_2_2748_1_a(.in(far_2_2748_0[0]), .out(far_2_2748_1[0]));    relay_conn far_2_2748_1_b(.in(far_2_2748_0[1]), .out(far_2_2748_1[1]));
    wire [1:0] far_2_2748_2;    relay_conn far_2_2748_2_a(.in(far_2_2748_1[0]), .out(far_2_2748_2[0]));    relay_conn far_2_2748_2_b(.in(far_2_2748_1[1]), .out(far_2_2748_2[1]));
    assign layer_2[708] = ~far_2_2748_2[0] | (far_2_2748_2[0] & far_2_2748_2[1]); 
    assign layer_2[709] = layer_1[248] & ~layer_1[217]; 
    wire [1:0] far_2_2750_0;    relay_conn far_2_2750_0_a(.in(layer_1[223]), .out(far_2_2750_0[0]));    relay_conn far_2_2750_0_b(.in(layer_1[294]), .out(far_2_2750_0[1]));
    wire [1:0] far_2_2750_1;    relay_conn far_2_2750_1_a(.in(far_2_2750_0[0]), .out(far_2_2750_1[0]));    relay_conn far_2_2750_1_b(.in(far_2_2750_0[1]), .out(far_2_2750_1[1]));
    assign layer_2[710] = far_2_2750_1[0] | far_2_2750_1[1]; 
    wire [1:0] far_2_2751_0;    relay_conn far_2_2751_0_a(.in(layer_1[661]), .out(far_2_2751_0[0]));    relay_conn far_2_2751_0_b(.in(layer_1[746]), .out(far_2_2751_0[1]));
    wire [1:0] far_2_2751_1;    relay_conn far_2_2751_1_a(.in(far_2_2751_0[0]), .out(far_2_2751_1[0]));    relay_conn far_2_2751_1_b(.in(far_2_2751_0[1]), .out(far_2_2751_1[1]));
    assign layer_2[711] = far_2_2751_1[0] ^ far_2_2751_1[1]; 
    wire [1:0] far_2_2752_0;    relay_conn far_2_2752_0_a(.in(layer_1[220]), .out(far_2_2752_0[0]));    relay_conn far_2_2752_0_b(.in(layer_1[104]), .out(far_2_2752_0[1]));
    wire [1:0] far_2_2752_1;    relay_conn far_2_2752_1_a(.in(far_2_2752_0[0]), .out(far_2_2752_1[0]));    relay_conn far_2_2752_1_b(.in(far_2_2752_0[1]), .out(far_2_2752_1[1]));
    wire [1:0] far_2_2752_2;    relay_conn far_2_2752_2_a(.in(far_2_2752_1[0]), .out(far_2_2752_2[0]));    relay_conn far_2_2752_2_b(.in(far_2_2752_1[1]), .out(far_2_2752_2[1]));
    assign layer_2[712] = ~far_2_2752_2[0] | (far_2_2752_2[0] & far_2_2752_2[1]); 
    wire [1:0] far_2_2753_0;    relay_conn far_2_2753_0_a(.in(layer_1[55]), .out(far_2_2753_0[0]));    relay_conn far_2_2753_0_b(.in(layer_1[152]), .out(far_2_2753_0[1]));
    wire [1:0] far_2_2753_1;    relay_conn far_2_2753_1_a(.in(far_2_2753_0[0]), .out(far_2_2753_1[0]));    relay_conn far_2_2753_1_b(.in(far_2_2753_0[1]), .out(far_2_2753_1[1]));
    wire [1:0] far_2_2753_2;    relay_conn far_2_2753_2_a(.in(far_2_2753_1[0]), .out(far_2_2753_2[0]));    relay_conn far_2_2753_2_b(.in(far_2_2753_1[1]), .out(far_2_2753_2[1]));
    assign layer_2[713] = far_2_2753_2[0] & far_2_2753_2[1]; 
    wire [1:0] far_2_2754_0;    relay_conn far_2_2754_0_a(.in(layer_1[525]), .out(far_2_2754_0[0]));    relay_conn far_2_2754_0_b(.in(layer_1[622]), .out(far_2_2754_0[1]));
    wire [1:0] far_2_2754_1;    relay_conn far_2_2754_1_a(.in(far_2_2754_0[0]), .out(far_2_2754_1[0]));    relay_conn far_2_2754_1_b(.in(far_2_2754_0[1]), .out(far_2_2754_1[1]));
    wire [1:0] far_2_2754_2;    relay_conn far_2_2754_2_a(.in(far_2_2754_1[0]), .out(far_2_2754_2[0]));    relay_conn far_2_2754_2_b(.in(far_2_2754_1[1]), .out(far_2_2754_2[1]));
    assign layer_2[714] = ~far_2_2754_2[0] | (far_2_2754_2[0] & far_2_2754_2[1]); 
    wire [1:0] far_2_2755_0;    relay_conn far_2_2755_0_a(.in(layer_1[514]), .out(far_2_2755_0[0]));    relay_conn far_2_2755_0_b(.in(layer_1[595]), .out(far_2_2755_0[1]));
    wire [1:0] far_2_2755_1;    relay_conn far_2_2755_1_a(.in(far_2_2755_0[0]), .out(far_2_2755_1[0]));    relay_conn far_2_2755_1_b(.in(far_2_2755_0[1]), .out(far_2_2755_1[1]));
    assign layer_2[715] = far_2_2755_1[0] & far_2_2755_1[1]; 
    wire [1:0] far_2_2756_0;    relay_conn far_2_2756_0_a(.in(layer_1[598]), .out(far_2_2756_0[0]));    relay_conn far_2_2756_0_b(.in(layer_1[497]), .out(far_2_2756_0[1]));
    wire [1:0] far_2_2756_1;    relay_conn far_2_2756_1_a(.in(far_2_2756_0[0]), .out(far_2_2756_1[0]));    relay_conn far_2_2756_1_b(.in(far_2_2756_0[1]), .out(far_2_2756_1[1]));
    wire [1:0] far_2_2756_2;    relay_conn far_2_2756_2_a(.in(far_2_2756_1[0]), .out(far_2_2756_2[0]));    relay_conn far_2_2756_2_b(.in(far_2_2756_1[1]), .out(far_2_2756_2[1]));
    assign layer_2[716] = far_2_2756_2[0]; 
    wire [1:0] far_2_2757_0;    relay_conn far_2_2757_0_a(.in(layer_1[731]), .out(far_2_2757_0[0]));    relay_conn far_2_2757_0_b(.in(layer_1[795]), .out(far_2_2757_0[1]));
    wire [1:0] far_2_2757_1;    relay_conn far_2_2757_1_a(.in(far_2_2757_0[0]), .out(far_2_2757_1[0]));    relay_conn far_2_2757_1_b(.in(far_2_2757_0[1]), .out(far_2_2757_1[1]));
    assign layer_2[717] = far_2_2757_1[0]; 
    wire [1:0] far_2_2758_0;    relay_conn far_2_2758_0_a(.in(layer_1[669]), .out(far_2_2758_0[0]));    relay_conn far_2_2758_0_b(.in(layer_1[796]), .out(far_2_2758_0[1]));
    wire [1:0] far_2_2758_1;    relay_conn far_2_2758_1_a(.in(far_2_2758_0[0]), .out(far_2_2758_1[0]));    relay_conn far_2_2758_1_b(.in(far_2_2758_0[1]), .out(far_2_2758_1[1]));
    wire [1:0] far_2_2758_2;    relay_conn far_2_2758_2_a(.in(far_2_2758_1[0]), .out(far_2_2758_2[0]));    relay_conn far_2_2758_2_b(.in(far_2_2758_1[1]), .out(far_2_2758_2[1]));
    assign layer_2[718] = ~far_2_2758_2[1]; 
    wire [1:0] far_2_2759_0;    relay_conn far_2_2759_0_a(.in(layer_1[674]), .out(far_2_2759_0[0]));    relay_conn far_2_2759_0_b(.in(layer_1[620]), .out(far_2_2759_0[1]));
    assign layer_2[719] = ~far_2_2759_0[1] | (far_2_2759_0[0] & far_2_2759_0[1]); 
    wire [1:0] far_2_2760_0;    relay_conn far_2_2760_0_a(.in(layer_1[680]), .out(far_2_2760_0[0]));    relay_conn far_2_2760_0_b(.in(layer_1[720]), .out(far_2_2760_0[1]));
    assign layer_2[720] = far_2_2760_0[1] & ~far_2_2760_0[0]; 
    wire [1:0] far_2_2761_0;    relay_conn far_2_2761_0_a(.in(layer_1[166]), .out(far_2_2761_0[0]));    relay_conn far_2_2761_0_b(.in(layer_1[95]), .out(far_2_2761_0[1]));
    wire [1:0] far_2_2761_1;    relay_conn far_2_2761_1_a(.in(far_2_2761_0[0]), .out(far_2_2761_1[0]));    relay_conn far_2_2761_1_b(.in(far_2_2761_0[1]), .out(far_2_2761_1[1]));
    assign layer_2[721] = ~far_2_2761_1[0] | (far_2_2761_1[0] & far_2_2761_1[1]); 
    wire [1:0] far_2_2762_0;    relay_conn far_2_2762_0_a(.in(layer_1[67]), .out(far_2_2762_0[0]));    relay_conn far_2_2762_0_b(.in(layer_1[6]), .out(far_2_2762_0[1]));
    assign layer_2[722] = far_2_2762_0[0]; 
    wire [1:0] far_2_2763_0;    relay_conn far_2_2763_0_a(.in(layer_1[671]), .out(far_2_2763_0[0]));    relay_conn far_2_2763_0_b(.in(layer_1[589]), .out(far_2_2763_0[1]));
    wire [1:0] far_2_2763_1;    relay_conn far_2_2763_1_a(.in(far_2_2763_0[0]), .out(far_2_2763_1[0]));    relay_conn far_2_2763_1_b(.in(far_2_2763_0[1]), .out(far_2_2763_1[1]));
    assign layer_2[723] = ~(far_2_2763_1[0] | far_2_2763_1[1]); 
    wire [1:0] far_2_2764_0;    relay_conn far_2_2764_0_a(.in(layer_1[105]), .out(far_2_2764_0[0]));    relay_conn far_2_2764_0_b(.in(layer_1[8]), .out(far_2_2764_0[1]));
    wire [1:0] far_2_2764_1;    relay_conn far_2_2764_1_a(.in(far_2_2764_0[0]), .out(far_2_2764_1[0]));    relay_conn far_2_2764_1_b(.in(far_2_2764_0[1]), .out(far_2_2764_1[1]));
    wire [1:0] far_2_2764_2;    relay_conn far_2_2764_2_a(.in(far_2_2764_1[0]), .out(far_2_2764_2[0]));    relay_conn far_2_2764_2_b(.in(far_2_2764_1[1]), .out(far_2_2764_2[1]));
    assign layer_2[724] = ~far_2_2764_2[0]; 
    wire [1:0] far_2_2765_0;    relay_conn far_2_2765_0_a(.in(layer_1[877]), .out(far_2_2765_0[0]));    relay_conn far_2_2765_0_b(.in(layer_1[796]), .out(far_2_2765_0[1]));
    wire [1:0] far_2_2765_1;    relay_conn far_2_2765_1_a(.in(far_2_2765_0[0]), .out(far_2_2765_1[0]));    relay_conn far_2_2765_1_b(.in(far_2_2765_0[1]), .out(far_2_2765_1[1]));
    assign layer_2[725] = ~far_2_2765_1[1] | (far_2_2765_1[0] & far_2_2765_1[1]); 
    assign layer_2[726] = ~layer_1[207] | (layer_1[207] & layer_1[218]); 
    assign layer_2[727] = layer_1[221]; 
    wire [1:0] far_2_2768_0;    relay_conn far_2_2768_0_a(.in(layer_1[520]), .out(far_2_2768_0[0]));    relay_conn far_2_2768_0_b(.in(layer_1[444]), .out(far_2_2768_0[1]));
    wire [1:0] far_2_2768_1;    relay_conn far_2_2768_1_a(.in(far_2_2768_0[0]), .out(far_2_2768_1[0]));    relay_conn far_2_2768_1_b(.in(far_2_2768_0[1]), .out(far_2_2768_1[1]));
    assign layer_2[728] = far_2_2768_1[1]; 
    assign layer_2[729] = layer_1[842] | layer_1[844]; 
    assign layer_2[730] = layer_1[958] & ~layer_1[932]; 
    wire [1:0] far_2_2771_0;    relay_conn far_2_2771_0_a(.in(layer_1[139]), .out(far_2_2771_0[0]));    relay_conn far_2_2771_0_b(.in(layer_1[70]), .out(far_2_2771_0[1]));
    wire [1:0] far_2_2771_1;    relay_conn far_2_2771_1_a(.in(far_2_2771_0[0]), .out(far_2_2771_1[0]));    relay_conn far_2_2771_1_b(.in(far_2_2771_0[1]), .out(far_2_2771_1[1]));
    assign layer_2[731] = far_2_2771_1[0] & far_2_2771_1[1]; 
    wire [1:0] far_2_2772_0;    relay_conn far_2_2772_0_a(.in(layer_1[89]), .out(far_2_2772_0[0]));    relay_conn far_2_2772_0_b(.in(layer_1[141]), .out(far_2_2772_0[1]));
    assign layer_2[732] = far_2_2772_0[0] & ~far_2_2772_0[1]; 
    wire [1:0] far_2_2773_0;    relay_conn far_2_2773_0_a(.in(layer_1[538]), .out(far_2_2773_0[0]));    relay_conn far_2_2773_0_b(.in(layer_1[617]), .out(far_2_2773_0[1]));
    wire [1:0] far_2_2773_1;    relay_conn far_2_2773_1_a(.in(far_2_2773_0[0]), .out(far_2_2773_1[0]));    relay_conn far_2_2773_1_b(.in(far_2_2773_0[1]), .out(far_2_2773_1[1]));
    assign layer_2[733] = far_2_2773_1[0] & ~far_2_2773_1[1]; 
    wire [1:0] far_2_2774_0;    relay_conn far_2_2774_0_a(.in(layer_1[796]), .out(far_2_2774_0[0]));    relay_conn far_2_2774_0_b(.in(layer_1[743]), .out(far_2_2774_0[1]));
    assign layer_2[734] = far_2_2774_0[1] & ~far_2_2774_0[0]; 
    wire [1:0] far_2_2775_0;    relay_conn far_2_2775_0_a(.in(layer_1[1008]), .out(far_2_2775_0[0]));    relay_conn far_2_2775_0_b(.in(layer_1[913]), .out(far_2_2775_0[1]));
    wire [1:0] far_2_2775_1;    relay_conn far_2_2775_1_a(.in(far_2_2775_0[0]), .out(far_2_2775_1[0]));    relay_conn far_2_2775_1_b(.in(far_2_2775_0[1]), .out(far_2_2775_1[1]));
    assign layer_2[735] = far_2_2775_1[1]; 
    assign layer_2[736] = ~layer_1[115]; 
    assign layer_2[737] = layer_1[368] & ~layer_1[342]; 
    wire [1:0] far_2_2778_0;    relay_conn far_2_2778_0_a(.in(layer_1[927]), .out(far_2_2778_0[0]));    relay_conn far_2_2778_0_b(.in(layer_1[874]), .out(far_2_2778_0[1]));
    assign layer_2[738] = far_2_2778_0[1]; 
    wire [1:0] far_2_2779_0;    relay_conn far_2_2779_0_a(.in(layer_1[787]), .out(far_2_2779_0[0]));    relay_conn far_2_2779_0_b(.in(layer_1[700]), .out(far_2_2779_0[1]));
    wire [1:0] far_2_2779_1;    relay_conn far_2_2779_1_a(.in(far_2_2779_0[0]), .out(far_2_2779_1[0]));    relay_conn far_2_2779_1_b(.in(far_2_2779_0[1]), .out(far_2_2779_1[1]));
    assign layer_2[739] = ~far_2_2779_1[0] | (far_2_2779_1[0] & far_2_2779_1[1]); 
    wire [1:0] far_2_2780_0;    relay_conn far_2_2780_0_a(.in(layer_1[615]), .out(far_2_2780_0[0]));    relay_conn far_2_2780_0_b(.in(layer_1[567]), .out(far_2_2780_0[1]));
    assign layer_2[740] = ~far_2_2780_0[1] | (far_2_2780_0[0] & far_2_2780_0[1]); 
    wire [1:0] far_2_2781_0;    relay_conn far_2_2781_0_a(.in(layer_1[882]), .out(far_2_2781_0[0]));    relay_conn far_2_2781_0_b(.in(layer_1[980]), .out(far_2_2781_0[1]));
    wire [1:0] far_2_2781_1;    relay_conn far_2_2781_1_a(.in(far_2_2781_0[0]), .out(far_2_2781_1[0]));    relay_conn far_2_2781_1_b(.in(far_2_2781_0[1]), .out(far_2_2781_1[1]));
    wire [1:0] far_2_2781_2;    relay_conn far_2_2781_2_a(.in(far_2_2781_1[0]), .out(far_2_2781_2[0]));    relay_conn far_2_2781_2_b(.in(far_2_2781_1[1]), .out(far_2_2781_2[1]));
    assign layer_2[741] = ~far_2_2781_2[0]; 
    wire [1:0] far_2_2782_0;    relay_conn far_2_2782_0_a(.in(layer_1[898]), .out(far_2_2782_0[0]));    relay_conn far_2_2782_0_b(.in(layer_1[935]), .out(far_2_2782_0[1]));
    assign layer_2[742] = ~far_2_2782_0[0]; 
    assign layer_2[743] = layer_1[63] | layer_1[58]; 
    assign layer_2[744] = layer_1[341] & layer_1[316]; 
    wire [1:0] far_2_2785_0;    relay_conn far_2_2785_0_a(.in(layer_1[257]), .out(far_2_2785_0[0]));    relay_conn far_2_2785_0_b(.in(layer_1[141]), .out(far_2_2785_0[1]));
    wire [1:0] far_2_2785_1;    relay_conn far_2_2785_1_a(.in(far_2_2785_0[0]), .out(far_2_2785_1[0]));    relay_conn far_2_2785_1_b(.in(far_2_2785_0[1]), .out(far_2_2785_1[1]));
    wire [1:0] far_2_2785_2;    relay_conn far_2_2785_2_a(.in(far_2_2785_1[0]), .out(far_2_2785_2[0]));    relay_conn far_2_2785_2_b(.in(far_2_2785_1[1]), .out(far_2_2785_2[1]));
    assign layer_2[745] = ~far_2_2785_2[1] | (far_2_2785_2[0] & far_2_2785_2[1]); 
    wire [1:0] far_2_2786_0;    relay_conn far_2_2786_0_a(.in(layer_1[877]), .out(far_2_2786_0[0]));    relay_conn far_2_2786_0_b(.in(layer_1[828]), .out(far_2_2786_0[1]));
    assign layer_2[746] = ~(far_2_2786_0[0] | far_2_2786_0[1]); 
    wire [1:0] far_2_2787_0;    relay_conn far_2_2787_0_a(.in(layer_1[507]), .out(far_2_2787_0[0]));    relay_conn far_2_2787_0_b(.in(layer_1[567]), .out(far_2_2787_0[1]));
    assign layer_2[747] = far_2_2787_0[0] & far_2_2787_0[1]; 
    assign layer_2[748] = layer_1[988]; 
    wire [1:0] far_2_2789_0;    relay_conn far_2_2789_0_a(.in(layer_1[838]), .out(far_2_2789_0[0]));    relay_conn far_2_2789_0_b(.in(layer_1[801]), .out(far_2_2789_0[1]));
    assign layer_2[749] = ~(far_2_2789_0[0] | far_2_2789_0[1]); 
    wire [1:0] far_2_2790_0;    relay_conn far_2_2790_0_a(.in(layer_1[531]), .out(far_2_2790_0[0]));    relay_conn far_2_2790_0_b(.in(layer_1[460]), .out(far_2_2790_0[1]));
    wire [1:0] far_2_2790_1;    relay_conn far_2_2790_1_a(.in(far_2_2790_0[0]), .out(far_2_2790_1[0]));    relay_conn far_2_2790_1_b(.in(far_2_2790_0[1]), .out(far_2_2790_1[1]));
    assign layer_2[750] = far_2_2790_1[0] & far_2_2790_1[1]; 
    wire [1:0] far_2_2791_0;    relay_conn far_2_2791_0_a(.in(layer_1[612]), .out(far_2_2791_0[0]));    relay_conn far_2_2791_0_b(.in(layer_1[720]), .out(far_2_2791_0[1]));
    wire [1:0] far_2_2791_1;    relay_conn far_2_2791_1_a(.in(far_2_2791_0[0]), .out(far_2_2791_1[0]));    relay_conn far_2_2791_1_b(.in(far_2_2791_0[1]), .out(far_2_2791_1[1]));
    wire [1:0] far_2_2791_2;    relay_conn far_2_2791_2_a(.in(far_2_2791_1[0]), .out(far_2_2791_2[0]));    relay_conn far_2_2791_2_b(.in(far_2_2791_1[1]), .out(far_2_2791_2[1]));
    assign layer_2[751] = ~(far_2_2791_2[0] & far_2_2791_2[1]); 
    wire [1:0] far_2_2792_0;    relay_conn far_2_2792_0_a(.in(layer_1[796]), .out(far_2_2792_0[0]));    relay_conn far_2_2792_0_b(.in(layer_1[735]), .out(far_2_2792_0[1]));
    assign layer_2[752] = ~(far_2_2792_0[0] ^ far_2_2792_0[1]); 
    wire [1:0] far_2_2793_0;    relay_conn far_2_2793_0_a(.in(layer_1[97]), .out(far_2_2793_0[0]));    relay_conn far_2_2793_0_b(.in(layer_1[139]), .out(far_2_2793_0[1]));
    assign layer_2[753] = far_2_2793_0[0] ^ far_2_2793_0[1]; 
    wire [1:0] far_2_2794_0;    relay_conn far_2_2794_0_a(.in(layer_1[603]), .out(far_2_2794_0[0]));    relay_conn far_2_2794_0_b(.in(layer_1[648]), .out(far_2_2794_0[1]));
    assign layer_2[754] = far_2_2794_0[0] & far_2_2794_0[1]; 
    assign layer_2[755] = layer_1[780] & ~layer_1[796]; 
    wire [1:0] far_2_2796_0;    relay_conn far_2_2796_0_a(.in(layer_1[285]), .out(far_2_2796_0[0]));    relay_conn far_2_2796_0_b(.in(layer_1[401]), .out(far_2_2796_0[1]));
    wire [1:0] far_2_2796_1;    relay_conn far_2_2796_1_a(.in(far_2_2796_0[0]), .out(far_2_2796_1[0]));    relay_conn far_2_2796_1_b(.in(far_2_2796_0[1]), .out(far_2_2796_1[1]));
    wire [1:0] far_2_2796_2;    relay_conn far_2_2796_2_a(.in(far_2_2796_1[0]), .out(far_2_2796_2[0]));    relay_conn far_2_2796_2_b(.in(far_2_2796_1[1]), .out(far_2_2796_2[1]));
    assign layer_2[756] = far_2_2796_2[0] & ~far_2_2796_2[1]; 
    wire [1:0] far_2_2797_0;    relay_conn far_2_2797_0_a(.in(layer_1[696]), .out(far_2_2797_0[0]));    relay_conn far_2_2797_0_b(.in(layer_1[771]), .out(far_2_2797_0[1]));
    wire [1:0] far_2_2797_1;    relay_conn far_2_2797_1_a(.in(far_2_2797_0[0]), .out(far_2_2797_1[0]));    relay_conn far_2_2797_1_b(.in(far_2_2797_0[1]), .out(far_2_2797_1[1]));
    assign layer_2[757] = far_2_2797_1[0] | far_2_2797_1[1]; 
    wire [1:0] far_2_2798_0;    relay_conn far_2_2798_0_a(.in(layer_1[734]), .out(far_2_2798_0[0]));    relay_conn far_2_2798_0_b(.in(layer_1[652]), .out(far_2_2798_0[1]));
    wire [1:0] far_2_2798_1;    relay_conn far_2_2798_1_a(.in(far_2_2798_0[0]), .out(far_2_2798_1[0]));    relay_conn far_2_2798_1_b(.in(far_2_2798_0[1]), .out(far_2_2798_1[1]));
    assign layer_2[758] = ~(far_2_2798_1[0] & far_2_2798_1[1]); 
    wire [1:0] far_2_2799_0;    relay_conn far_2_2799_0_a(.in(layer_1[701]), .out(far_2_2799_0[0]));    relay_conn far_2_2799_0_b(.in(layer_1[817]), .out(far_2_2799_0[1]));
    wire [1:0] far_2_2799_1;    relay_conn far_2_2799_1_a(.in(far_2_2799_0[0]), .out(far_2_2799_1[0]));    relay_conn far_2_2799_1_b(.in(far_2_2799_0[1]), .out(far_2_2799_1[1]));
    wire [1:0] far_2_2799_2;    relay_conn far_2_2799_2_a(.in(far_2_2799_1[0]), .out(far_2_2799_2[0]));    relay_conn far_2_2799_2_b(.in(far_2_2799_1[1]), .out(far_2_2799_2[1]));
    assign layer_2[759] = far_2_2799_2[0] ^ far_2_2799_2[1]; 
    assign layer_2[760] = layer_1[980] & ~layer_1[986]; 
    wire [1:0] far_2_2801_0;    relay_conn far_2_2801_0_a(.in(layer_1[293]), .out(far_2_2801_0[0]));    relay_conn far_2_2801_0_b(.in(layer_1[259]), .out(far_2_2801_0[1]));
    assign layer_2[761] = ~far_2_2801_0[0]; 
    wire [1:0] far_2_2802_0;    relay_conn far_2_2802_0_a(.in(layer_1[795]), .out(far_2_2802_0[0]));    relay_conn far_2_2802_0_b(.in(layer_1[869]), .out(far_2_2802_0[1]));
    wire [1:0] far_2_2802_1;    relay_conn far_2_2802_1_a(.in(far_2_2802_0[0]), .out(far_2_2802_1[0]));    relay_conn far_2_2802_1_b(.in(far_2_2802_0[1]), .out(far_2_2802_1[1]));
    assign layer_2[762] = ~(far_2_2802_1[0] ^ far_2_2802_1[1]); 
    wire [1:0] far_2_2803_0;    relay_conn far_2_2803_0_a(.in(layer_1[430]), .out(far_2_2803_0[0]));    relay_conn far_2_2803_0_b(.in(layer_1[533]), .out(far_2_2803_0[1]));
    wire [1:0] far_2_2803_1;    relay_conn far_2_2803_1_a(.in(far_2_2803_0[0]), .out(far_2_2803_1[0]));    relay_conn far_2_2803_1_b(.in(far_2_2803_0[1]), .out(far_2_2803_1[1]));
    wire [1:0] far_2_2803_2;    relay_conn far_2_2803_2_a(.in(far_2_2803_1[0]), .out(far_2_2803_2[0]));    relay_conn far_2_2803_2_b(.in(far_2_2803_1[1]), .out(far_2_2803_2[1]));
    assign layer_2[763] = far_2_2803_2[0] & far_2_2803_2[1]; 
    wire [1:0] far_2_2804_0;    relay_conn far_2_2804_0_a(.in(layer_1[429]), .out(far_2_2804_0[0]));    relay_conn far_2_2804_0_b(.in(layer_1[363]), .out(far_2_2804_0[1]));
    wire [1:0] far_2_2804_1;    relay_conn far_2_2804_1_a(.in(far_2_2804_0[0]), .out(far_2_2804_1[0]));    relay_conn far_2_2804_1_b(.in(far_2_2804_0[1]), .out(far_2_2804_1[1]));
    assign layer_2[764] = ~(far_2_2804_1[0] | far_2_2804_1[1]); 
    assign layer_2[765] = layer_1[563] & ~layer_1[585]; 
    assign layer_2[766] = layer_1[64]; 
    assign layer_2[767] = ~layer_1[967]; 
    wire [1:0] far_2_2808_0;    relay_conn far_2_2808_0_a(.in(layer_1[291]), .out(far_2_2808_0[0]));    relay_conn far_2_2808_0_b(.in(layer_1[232]), .out(far_2_2808_0[1]));
    assign layer_2[768] = ~(far_2_2808_0[0] & far_2_2808_0[1]); 
    wire [1:0] far_2_2809_0;    relay_conn far_2_2809_0_a(.in(layer_1[77]), .out(far_2_2809_0[0]));    relay_conn far_2_2809_0_b(.in(layer_1[133]), .out(far_2_2809_0[1]));
    assign layer_2[769] = ~far_2_2809_0[0]; 
    wire [1:0] far_2_2810_0;    relay_conn far_2_2810_0_a(.in(layer_1[428]), .out(far_2_2810_0[0]));    relay_conn far_2_2810_0_b(.in(layer_1[358]), .out(far_2_2810_0[1]));
    wire [1:0] far_2_2810_1;    relay_conn far_2_2810_1_a(.in(far_2_2810_0[0]), .out(far_2_2810_1[0]));    relay_conn far_2_2810_1_b(.in(far_2_2810_0[1]), .out(far_2_2810_1[1]));
    assign layer_2[770] = far_2_2810_1[1]; 
    wire [1:0] far_2_2811_0;    relay_conn far_2_2811_0_a(.in(layer_1[173]), .out(far_2_2811_0[0]));    relay_conn far_2_2811_0_b(.in(layer_1[267]), .out(far_2_2811_0[1]));
    wire [1:0] far_2_2811_1;    relay_conn far_2_2811_1_a(.in(far_2_2811_0[0]), .out(far_2_2811_1[0]));    relay_conn far_2_2811_1_b(.in(far_2_2811_0[1]), .out(far_2_2811_1[1]));
    assign layer_2[771] = ~(far_2_2811_1[0] & far_2_2811_1[1]); 
    wire [1:0] far_2_2812_0;    relay_conn far_2_2812_0_a(.in(layer_1[307]), .out(far_2_2812_0[0]));    relay_conn far_2_2812_0_b(.in(layer_1[409]), .out(far_2_2812_0[1]));
    wire [1:0] far_2_2812_1;    relay_conn far_2_2812_1_a(.in(far_2_2812_0[0]), .out(far_2_2812_1[0]));    relay_conn far_2_2812_1_b(.in(far_2_2812_0[1]), .out(far_2_2812_1[1]));
    wire [1:0] far_2_2812_2;    relay_conn far_2_2812_2_a(.in(far_2_2812_1[0]), .out(far_2_2812_2[0]));    relay_conn far_2_2812_2_b(.in(far_2_2812_1[1]), .out(far_2_2812_2[1]));
    assign layer_2[772] = ~far_2_2812_2[1]; 
    wire [1:0] far_2_2813_0;    relay_conn far_2_2813_0_a(.in(layer_1[985]), .out(far_2_2813_0[0]));    relay_conn far_2_2813_0_b(.in(layer_1[950]), .out(far_2_2813_0[1]));
    assign layer_2[773] = ~(far_2_2813_0[0] & far_2_2813_0[1]); 
    wire [1:0] far_2_2814_0;    relay_conn far_2_2814_0_a(.in(layer_1[113]), .out(far_2_2814_0[0]));    relay_conn far_2_2814_0_b(.in(layer_1[213]), .out(far_2_2814_0[1]));
    wire [1:0] far_2_2814_1;    relay_conn far_2_2814_1_a(.in(far_2_2814_0[0]), .out(far_2_2814_1[0]));    relay_conn far_2_2814_1_b(.in(far_2_2814_0[1]), .out(far_2_2814_1[1]));
    wire [1:0] far_2_2814_2;    relay_conn far_2_2814_2_a(.in(far_2_2814_1[0]), .out(far_2_2814_2[0]));    relay_conn far_2_2814_2_b(.in(far_2_2814_1[1]), .out(far_2_2814_2[1]));
    assign layer_2[774] = far_2_2814_2[1] & ~far_2_2814_2[0]; 
    wire [1:0] far_2_2815_0;    relay_conn far_2_2815_0_a(.in(layer_1[740]), .out(far_2_2815_0[0]));    relay_conn far_2_2815_0_b(.in(layer_1[673]), .out(far_2_2815_0[1]));
    wire [1:0] far_2_2815_1;    relay_conn far_2_2815_1_a(.in(far_2_2815_0[0]), .out(far_2_2815_1[0]));    relay_conn far_2_2815_1_b(.in(far_2_2815_0[1]), .out(far_2_2815_1[1]));
    assign layer_2[775] = far_2_2815_1[1] & ~far_2_2815_1[0]; 
    wire [1:0] far_2_2816_0;    relay_conn far_2_2816_0_a(.in(layer_1[1018]), .out(far_2_2816_0[0]));    relay_conn far_2_2816_0_b(.in(layer_1[917]), .out(far_2_2816_0[1]));
    wire [1:0] far_2_2816_1;    relay_conn far_2_2816_1_a(.in(far_2_2816_0[0]), .out(far_2_2816_1[0]));    relay_conn far_2_2816_1_b(.in(far_2_2816_0[1]), .out(far_2_2816_1[1]));
    wire [1:0] far_2_2816_2;    relay_conn far_2_2816_2_a(.in(far_2_2816_1[0]), .out(far_2_2816_2[0]));    relay_conn far_2_2816_2_b(.in(far_2_2816_1[1]), .out(far_2_2816_2[1]));
    assign layer_2[776] = far_2_2816_2[0]; 
    assign layer_2[777] = ~layer_1[162]; 
    wire [1:0] far_2_2818_0;    relay_conn far_2_2818_0_a(.in(layer_1[444]), .out(far_2_2818_0[0]));    relay_conn far_2_2818_0_b(.in(layer_1[404]), .out(far_2_2818_0[1]));
    assign layer_2[778] = far_2_2818_0[0] ^ far_2_2818_0[1]; 
    wire [1:0] far_2_2819_0;    relay_conn far_2_2819_0_a(.in(layer_1[444]), .out(far_2_2819_0[0]));    relay_conn far_2_2819_0_b(.in(layer_1[364]), .out(far_2_2819_0[1]));
    wire [1:0] far_2_2819_1;    relay_conn far_2_2819_1_a(.in(far_2_2819_0[0]), .out(far_2_2819_1[0]));    relay_conn far_2_2819_1_b(.in(far_2_2819_0[1]), .out(far_2_2819_1[1]));
    assign layer_2[779] = far_2_2819_1[0] & ~far_2_2819_1[1]; 
    wire [1:0] far_2_2820_0;    relay_conn far_2_2820_0_a(.in(layer_1[408]), .out(far_2_2820_0[0]));    relay_conn far_2_2820_0_b(.in(layer_1[353]), .out(far_2_2820_0[1]));
    assign layer_2[780] = ~(far_2_2820_0[0] | far_2_2820_0[1]); 
    assign layer_2[781] = layer_1[132] & ~layer_1[141]; 
    wire [1:0] far_2_2822_0;    relay_conn far_2_2822_0_a(.in(layer_1[796]), .out(far_2_2822_0[0]));    relay_conn far_2_2822_0_b(.in(layer_1[724]), .out(far_2_2822_0[1]));
    wire [1:0] far_2_2822_1;    relay_conn far_2_2822_1_a(.in(far_2_2822_0[0]), .out(far_2_2822_1[0]));    relay_conn far_2_2822_1_b(.in(far_2_2822_0[1]), .out(far_2_2822_1[1]));
    assign layer_2[782] = ~(far_2_2822_1[0] & far_2_2822_1[1]); 
    wire [1:0] far_2_2823_0;    relay_conn far_2_2823_0_a(.in(layer_1[758]), .out(far_2_2823_0[0]));    relay_conn far_2_2823_0_b(.in(layer_1[837]), .out(far_2_2823_0[1]));
    wire [1:0] far_2_2823_1;    relay_conn far_2_2823_1_a(.in(far_2_2823_0[0]), .out(far_2_2823_1[0]));    relay_conn far_2_2823_1_b(.in(far_2_2823_0[1]), .out(far_2_2823_1[1]));
    assign layer_2[783] = far_2_2823_1[0] & ~far_2_2823_1[1]; 
    wire [1:0] far_2_2824_0;    relay_conn far_2_2824_0_a(.in(layer_1[731]), .out(far_2_2824_0[0]));    relay_conn far_2_2824_0_b(.in(layer_1[827]), .out(far_2_2824_0[1]));
    wire [1:0] far_2_2824_1;    relay_conn far_2_2824_1_a(.in(far_2_2824_0[0]), .out(far_2_2824_1[0]));    relay_conn far_2_2824_1_b(.in(far_2_2824_0[1]), .out(far_2_2824_1[1]));
    wire [1:0] far_2_2824_2;    relay_conn far_2_2824_2_a(.in(far_2_2824_1[0]), .out(far_2_2824_2[0]));    relay_conn far_2_2824_2_b(.in(far_2_2824_1[1]), .out(far_2_2824_2[1]));
    assign layer_2[784] = far_2_2824_2[0] & ~far_2_2824_2[1]; 
    assign layer_2[785] = ~(layer_1[377] | layer_1[385]); 
    wire [1:0] far_2_2826_0;    relay_conn far_2_2826_0_a(.in(layer_1[721]), .out(far_2_2826_0[0]));    relay_conn far_2_2826_0_b(.in(layer_1[596]), .out(far_2_2826_0[1]));
    wire [1:0] far_2_2826_1;    relay_conn far_2_2826_1_a(.in(far_2_2826_0[0]), .out(far_2_2826_1[0]));    relay_conn far_2_2826_1_b(.in(far_2_2826_0[1]), .out(far_2_2826_1[1]));
    wire [1:0] far_2_2826_2;    relay_conn far_2_2826_2_a(.in(far_2_2826_1[0]), .out(far_2_2826_2[0]));    relay_conn far_2_2826_2_b(.in(far_2_2826_1[1]), .out(far_2_2826_2[1]));
    assign layer_2[786] = ~far_2_2826_2[1] | (far_2_2826_2[0] & far_2_2826_2[1]); 
    wire [1:0] far_2_2827_0;    relay_conn far_2_2827_0_a(.in(layer_1[688]), .out(far_2_2827_0[0]));    relay_conn far_2_2827_0_b(.in(layer_1[723]), .out(far_2_2827_0[1]));
    assign layer_2[787] = ~(far_2_2827_0[0] | far_2_2827_0[1]); 
    assign layer_2[788] = layer_1[763] & ~layer_1[765]; 
    wire [1:0] far_2_2829_0;    relay_conn far_2_2829_0_a(.in(layer_1[180]), .out(far_2_2829_0[0]));    relay_conn far_2_2829_0_b(.in(layer_1[248]), .out(far_2_2829_0[1]));
    wire [1:0] far_2_2829_1;    relay_conn far_2_2829_1_a(.in(far_2_2829_0[0]), .out(far_2_2829_1[0]));    relay_conn far_2_2829_1_b(.in(far_2_2829_0[1]), .out(far_2_2829_1[1]));
    assign layer_2[789] = ~far_2_2829_1[1] | (far_2_2829_1[0] & far_2_2829_1[1]); 
    wire [1:0] far_2_2830_0;    relay_conn far_2_2830_0_a(.in(layer_1[807]), .out(far_2_2830_0[0]));    relay_conn far_2_2830_0_b(.in(layer_1[696]), .out(far_2_2830_0[1]));
    wire [1:0] far_2_2830_1;    relay_conn far_2_2830_1_a(.in(far_2_2830_0[0]), .out(far_2_2830_1[0]));    relay_conn far_2_2830_1_b(.in(far_2_2830_0[1]), .out(far_2_2830_1[1]));
    wire [1:0] far_2_2830_2;    relay_conn far_2_2830_2_a(.in(far_2_2830_1[0]), .out(far_2_2830_2[0]));    relay_conn far_2_2830_2_b(.in(far_2_2830_1[1]), .out(far_2_2830_2[1]));
    assign layer_2[790] = far_2_2830_2[0] & far_2_2830_2[1]; 
    wire [1:0] far_2_2831_0;    relay_conn far_2_2831_0_a(.in(layer_1[815]), .out(far_2_2831_0[0]));    relay_conn far_2_2831_0_b(.in(layer_1[707]), .out(far_2_2831_0[1]));
    wire [1:0] far_2_2831_1;    relay_conn far_2_2831_1_a(.in(far_2_2831_0[0]), .out(far_2_2831_1[0]));    relay_conn far_2_2831_1_b(.in(far_2_2831_0[1]), .out(far_2_2831_1[1]));
    wire [1:0] far_2_2831_2;    relay_conn far_2_2831_2_a(.in(far_2_2831_1[0]), .out(far_2_2831_2[0]));    relay_conn far_2_2831_2_b(.in(far_2_2831_1[1]), .out(far_2_2831_2[1]));
    assign layer_2[791] = far_2_2831_2[0] & ~far_2_2831_2[1]; 
    wire [1:0] far_2_2832_0;    relay_conn far_2_2832_0_a(.in(layer_1[217]), .out(far_2_2832_0[0]));    relay_conn far_2_2832_0_b(.in(layer_1[270]), .out(far_2_2832_0[1]));
    assign layer_2[792] = far_2_2832_0[0] | far_2_2832_0[1]; 
    assign layer_2[793] = ~(layer_1[501] & layer_1[517]); 
    wire [1:0] far_2_2834_0;    relay_conn far_2_2834_0_a(.in(layer_1[875]), .out(far_2_2834_0[0]));    relay_conn far_2_2834_0_b(.in(layer_1[771]), .out(far_2_2834_0[1]));
    wire [1:0] far_2_2834_1;    relay_conn far_2_2834_1_a(.in(far_2_2834_0[0]), .out(far_2_2834_1[0]));    relay_conn far_2_2834_1_b(.in(far_2_2834_0[1]), .out(far_2_2834_1[1]));
    wire [1:0] far_2_2834_2;    relay_conn far_2_2834_2_a(.in(far_2_2834_1[0]), .out(far_2_2834_2[0]));    relay_conn far_2_2834_2_b(.in(far_2_2834_1[1]), .out(far_2_2834_2[1]));
    assign layer_2[794] = ~far_2_2834_2[0] | (far_2_2834_2[0] & far_2_2834_2[1]); 
    wire [1:0] far_2_2835_0;    relay_conn far_2_2835_0_a(.in(layer_1[213]), .out(far_2_2835_0[0]));    relay_conn far_2_2835_0_b(.in(layer_1[273]), .out(far_2_2835_0[1]));
    assign layer_2[795] = far_2_2835_0[0] & ~far_2_2835_0[1]; 
    assign layer_2[796] = ~(layer_1[257] | layer_1[228]); 
    wire [1:0] far_2_2837_0;    relay_conn far_2_2837_0_a(.in(layer_1[988]), .out(far_2_2837_0[0]));    relay_conn far_2_2837_0_b(.in(layer_1[951]), .out(far_2_2837_0[1]));
    assign layer_2[797] = ~far_2_2837_0[0] | (far_2_2837_0[0] & far_2_2837_0[1]); 
    wire [1:0] far_2_2838_0;    relay_conn far_2_2838_0_a(.in(layer_1[67]), .out(far_2_2838_0[0]));    relay_conn far_2_2838_0_b(.in(layer_1[101]), .out(far_2_2838_0[1]));
    assign layer_2[798] = far_2_2838_0[0] & far_2_2838_0[1]; 
    wire [1:0] far_2_2839_0;    relay_conn far_2_2839_0_a(.in(layer_1[430]), .out(far_2_2839_0[0]));    relay_conn far_2_2839_0_b(.in(layer_1[335]), .out(far_2_2839_0[1]));
    wire [1:0] far_2_2839_1;    relay_conn far_2_2839_1_a(.in(far_2_2839_0[0]), .out(far_2_2839_1[0]));    relay_conn far_2_2839_1_b(.in(far_2_2839_0[1]), .out(far_2_2839_1[1]));
    assign layer_2[799] = far_2_2839_1[1]; 
    wire [1:0] far_2_2840_0;    relay_conn far_2_2840_0_a(.in(layer_1[932]), .out(far_2_2840_0[0]));    relay_conn far_2_2840_0_b(.in(layer_1[1000]), .out(far_2_2840_0[1]));
    wire [1:0] far_2_2840_1;    relay_conn far_2_2840_1_a(.in(far_2_2840_0[0]), .out(far_2_2840_1[0]));    relay_conn far_2_2840_1_b(.in(far_2_2840_0[1]), .out(far_2_2840_1[1]));
    assign layer_2[800] = ~(far_2_2840_1[0] ^ far_2_2840_1[1]); 
    wire [1:0] far_2_2841_0;    relay_conn far_2_2841_0_a(.in(layer_1[555]), .out(far_2_2841_0[0]));    relay_conn far_2_2841_0_b(.in(layer_1[428]), .out(far_2_2841_0[1]));
    wire [1:0] far_2_2841_1;    relay_conn far_2_2841_1_a(.in(far_2_2841_0[0]), .out(far_2_2841_1[0]));    relay_conn far_2_2841_1_b(.in(far_2_2841_0[1]), .out(far_2_2841_1[1]));
    wire [1:0] far_2_2841_2;    relay_conn far_2_2841_2_a(.in(far_2_2841_1[0]), .out(far_2_2841_2[0]));    relay_conn far_2_2841_2_b(.in(far_2_2841_1[1]), .out(far_2_2841_2[1]));
    assign layer_2[801] = ~(far_2_2841_2[0] & far_2_2841_2[1]); 
    assign layer_2[802] = ~(layer_1[139] & layer_1[169]); 
    wire [1:0] far_2_2843_0;    relay_conn far_2_2843_0_a(.in(layer_1[379]), .out(far_2_2843_0[0]));    relay_conn far_2_2843_0_b(.in(layer_1[346]), .out(far_2_2843_0[1]));
    assign layer_2[803] = far_2_2843_0[0] & far_2_2843_0[1]; 
    assign layer_2[804] = layer_1[303]; 
    wire [1:0] far_2_2845_0;    relay_conn far_2_2845_0_a(.in(layer_1[533]), .out(far_2_2845_0[0]));    relay_conn far_2_2845_0_b(.in(layer_1[477]), .out(far_2_2845_0[1]));
    assign layer_2[805] = ~far_2_2845_0[1]; 
    assign layer_2[806] = layer_1[497] & ~layer_1[514]; 
    wire [1:0] far_2_2847_0;    relay_conn far_2_2847_0_a(.in(layer_1[8]), .out(far_2_2847_0[0]));    relay_conn far_2_2847_0_b(.in(layer_1[127]), .out(far_2_2847_0[1]));
    wire [1:0] far_2_2847_1;    relay_conn far_2_2847_1_a(.in(far_2_2847_0[0]), .out(far_2_2847_1[0]));    relay_conn far_2_2847_1_b(.in(far_2_2847_0[1]), .out(far_2_2847_1[1]));
    wire [1:0] far_2_2847_2;    relay_conn far_2_2847_2_a(.in(far_2_2847_1[0]), .out(far_2_2847_2[0]));    relay_conn far_2_2847_2_b(.in(far_2_2847_1[1]), .out(far_2_2847_2[1]));
    assign layer_2[807] = far_2_2847_2[0] & ~far_2_2847_2[1]; 
    assign layer_2[808] = layer_1[1007] ^ layer_1[1008]; 
    wire [1:0] far_2_2849_0;    relay_conn far_2_2849_0_a(.in(layer_1[663]), .out(far_2_2849_0[0]));    relay_conn far_2_2849_0_b(.in(layer_1[743]), .out(far_2_2849_0[1]));
    wire [1:0] far_2_2849_1;    relay_conn far_2_2849_1_a(.in(far_2_2849_0[0]), .out(far_2_2849_1[0]));    relay_conn far_2_2849_1_b(.in(far_2_2849_0[1]), .out(far_2_2849_1[1]));
    assign layer_2[809] = ~far_2_2849_1[1] | (far_2_2849_1[0] & far_2_2849_1[1]); 
    assign layer_2[810] = ~layer_1[756] | (layer_1[757] & layer_1[756]); 
    wire [1:0] far_2_2851_0;    relay_conn far_2_2851_0_a(.in(layer_1[312]), .out(far_2_2851_0[0]));    relay_conn far_2_2851_0_b(.in(layer_1[234]), .out(far_2_2851_0[1]));
    wire [1:0] far_2_2851_1;    relay_conn far_2_2851_1_a(.in(far_2_2851_0[0]), .out(far_2_2851_1[0]));    relay_conn far_2_2851_1_b(.in(far_2_2851_0[1]), .out(far_2_2851_1[1]));
    assign layer_2[811] = ~far_2_2851_1[1]; 
    wire [1:0] far_2_2852_0;    relay_conn far_2_2852_0_a(.in(layer_1[177]), .out(far_2_2852_0[0]));    relay_conn far_2_2852_0_b(.in(layer_1[270]), .out(far_2_2852_0[1]));
    wire [1:0] far_2_2852_1;    relay_conn far_2_2852_1_a(.in(far_2_2852_0[0]), .out(far_2_2852_1[0]));    relay_conn far_2_2852_1_b(.in(far_2_2852_0[1]), .out(far_2_2852_1[1]));
    assign layer_2[812] = far_2_2852_1[0] & far_2_2852_1[1]; 
    wire [1:0] far_2_2853_0;    relay_conn far_2_2853_0_a(.in(layer_1[694]), .out(far_2_2853_0[0]));    relay_conn far_2_2853_0_b(.in(layer_1[586]), .out(far_2_2853_0[1]));
    wire [1:0] far_2_2853_1;    relay_conn far_2_2853_1_a(.in(far_2_2853_0[0]), .out(far_2_2853_1[0]));    relay_conn far_2_2853_1_b(.in(far_2_2853_0[1]), .out(far_2_2853_1[1]));
    wire [1:0] far_2_2853_2;    relay_conn far_2_2853_2_a(.in(far_2_2853_1[0]), .out(far_2_2853_2[0]));    relay_conn far_2_2853_2_b(.in(far_2_2853_1[1]), .out(far_2_2853_2[1]));
    assign layer_2[813] = ~(far_2_2853_2[0] | far_2_2853_2[1]); 
    assign layer_2[814] = ~layer_1[546] | (layer_1[543] & layer_1[546]); 
    assign layer_2[815] = ~(layer_1[795] ^ layer_1[814]); 
    assign layer_2[816] = ~(layer_1[270] & layer_1[291]); 
    wire [1:0] far_2_2857_0;    relay_conn far_2_2857_0_a(.in(layer_1[152]), .out(far_2_2857_0[0]));    relay_conn far_2_2857_0_b(.in(layer_1[105]), .out(far_2_2857_0[1]));
    assign layer_2[817] = ~far_2_2857_0[1]; 
    wire [1:0] far_2_2858_0;    relay_conn far_2_2858_0_a(.in(layer_1[171]), .out(far_2_2858_0[0]));    relay_conn far_2_2858_0_b(.in(layer_1[259]), .out(far_2_2858_0[1]));
    wire [1:0] far_2_2858_1;    relay_conn far_2_2858_1_a(.in(far_2_2858_0[0]), .out(far_2_2858_1[0]));    relay_conn far_2_2858_1_b(.in(far_2_2858_0[1]), .out(far_2_2858_1[1]));
    assign layer_2[818] = far_2_2858_1[0] | far_2_2858_1[1]; 
    wire [1:0] far_2_2859_0;    relay_conn far_2_2859_0_a(.in(layer_1[962]), .out(far_2_2859_0[0]));    relay_conn far_2_2859_0_b(.in(layer_1[898]), .out(far_2_2859_0[1]));
    wire [1:0] far_2_2859_1;    relay_conn far_2_2859_1_a(.in(far_2_2859_0[0]), .out(far_2_2859_1[0]));    relay_conn far_2_2859_1_b(.in(far_2_2859_0[1]), .out(far_2_2859_1[1]));
    assign layer_2[819] = far_2_2859_1[0] | far_2_2859_1[1]; 
    wire [1:0] far_2_2860_0;    relay_conn far_2_2860_0_a(.in(layer_1[291]), .out(far_2_2860_0[0]));    relay_conn far_2_2860_0_b(.in(layer_1[409]), .out(far_2_2860_0[1]));
    wire [1:0] far_2_2860_1;    relay_conn far_2_2860_1_a(.in(far_2_2860_0[0]), .out(far_2_2860_1[0]));    relay_conn far_2_2860_1_b(.in(far_2_2860_0[1]), .out(far_2_2860_1[1]));
    wire [1:0] far_2_2860_2;    relay_conn far_2_2860_2_a(.in(far_2_2860_1[0]), .out(far_2_2860_2[0]));    relay_conn far_2_2860_2_b(.in(far_2_2860_1[1]), .out(far_2_2860_2[1]));
    assign layer_2[820] = far_2_2860_2[1] & ~far_2_2860_2[0]; 
    wire [1:0] far_2_2861_0;    relay_conn far_2_2861_0_a(.in(layer_1[596]), .out(far_2_2861_0[0]));    relay_conn far_2_2861_0_b(.in(layer_1[556]), .out(far_2_2861_0[1]));
    assign layer_2[821] = far_2_2861_0[0]; 
    wire [1:0] far_2_2862_0;    relay_conn far_2_2862_0_a(.in(layer_1[927]), .out(far_2_2862_0[0]));    relay_conn far_2_2862_0_b(.in(layer_1[999]), .out(far_2_2862_0[1]));
    wire [1:0] far_2_2862_1;    relay_conn far_2_2862_1_a(.in(far_2_2862_0[0]), .out(far_2_2862_1[0]));    relay_conn far_2_2862_1_b(.in(far_2_2862_0[1]), .out(far_2_2862_1[1]));
    assign layer_2[822] = ~far_2_2862_1[0]; 
    wire [1:0] far_2_2863_0;    relay_conn far_2_2863_0_a(.in(layer_1[988]), .out(far_2_2863_0[0]));    relay_conn far_2_2863_0_b(.in(layer_1[866]), .out(far_2_2863_0[1]));
    wire [1:0] far_2_2863_1;    relay_conn far_2_2863_1_a(.in(far_2_2863_0[0]), .out(far_2_2863_1[0]));    relay_conn far_2_2863_1_b(.in(far_2_2863_0[1]), .out(far_2_2863_1[1]));
    wire [1:0] far_2_2863_2;    relay_conn far_2_2863_2_a(.in(far_2_2863_1[0]), .out(far_2_2863_2[0]));    relay_conn far_2_2863_2_b(.in(far_2_2863_1[1]), .out(far_2_2863_2[1]));
    assign layer_2[823] = ~far_2_2863_2[0]; 
    wire [1:0] far_2_2864_0;    relay_conn far_2_2864_0_a(.in(layer_1[965]), .out(far_2_2864_0[0]));    relay_conn far_2_2864_0_b(.in(layer_1[922]), .out(far_2_2864_0[1]));
    assign layer_2[824] = far_2_2864_0[0] & ~far_2_2864_0[1]; 
    wire [1:0] far_2_2865_0;    relay_conn far_2_2865_0_a(.in(layer_1[28]), .out(far_2_2865_0[0]));    relay_conn far_2_2865_0_b(.in(layer_1[85]), .out(far_2_2865_0[1]));
    assign layer_2[825] = far_2_2865_0[0] & far_2_2865_0[1]; 
    wire [1:0] far_2_2866_0;    relay_conn far_2_2866_0_a(.in(layer_1[795]), .out(far_2_2866_0[0]));    relay_conn far_2_2866_0_b(.in(layer_1[747]), .out(far_2_2866_0[1]));
    assign layer_2[826] = ~far_2_2866_0[0]; 
    wire [1:0] far_2_2867_0;    relay_conn far_2_2867_0_a(.in(layer_1[561]), .out(far_2_2867_0[0]));    relay_conn far_2_2867_0_b(.in(layer_1[595]), .out(far_2_2867_0[1]));
    assign layer_2[827] = ~far_2_2867_0[1]; 
    assign layer_2[828] = ~(layer_1[627] & layer_1[605]); 
    wire [1:0] far_2_2869_0;    relay_conn far_2_2869_0_a(.in(layer_1[620]), .out(far_2_2869_0[0]));    relay_conn far_2_2869_0_b(.in(layer_1[692]), .out(far_2_2869_0[1]));
    wire [1:0] far_2_2869_1;    relay_conn far_2_2869_1_a(.in(far_2_2869_0[0]), .out(far_2_2869_1[0]));    relay_conn far_2_2869_1_b(.in(far_2_2869_0[1]), .out(far_2_2869_1[1]));
    assign layer_2[829] = ~far_2_2869_1[0] | (far_2_2869_1[0] & far_2_2869_1[1]); 
    wire [1:0] far_2_2870_0;    relay_conn far_2_2870_0_a(.in(layer_1[153]), .out(far_2_2870_0[0]));    relay_conn far_2_2870_0_b(.in(layer_1[186]), .out(far_2_2870_0[1]));
    assign layer_2[830] = ~(far_2_2870_0[0] & far_2_2870_0[1]); 
    wire [1:0] far_2_2871_0;    relay_conn far_2_2871_0_a(.in(layer_1[925]), .out(far_2_2871_0[0]));    relay_conn far_2_2871_0_b(.in(layer_1[874]), .out(far_2_2871_0[1]));
    assign layer_2[831] = far_2_2871_0[0] | far_2_2871_0[1]; 
    wire [1:0] far_2_2872_0;    relay_conn far_2_2872_0_a(.in(layer_1[494]), .out(far_2_2872_0[0]));    relay_conn far_2_2872_0_b(.in(layer_1[432]), .out(far_2_2872_0[1]));
    assign layer_2[832] = ~far_2_2872_0[0] | (far_2_2872_0[0] & far_2_2872_0[1]); 
    wire [1:0] far_2_2873_0;    relay_conn far_2_2873_0_a(.in(layer_1[828]), .out(far_2_2873_0[0]));    relay_conn far_2_2873_0_b(.in(layer_1[734]), .out(far_2_2873_0[1]));
    wire [1:0] far_2_2873_1;    relay_conn far_2_2873_1_a(.in(far_2_2873_0[0]), .out(far_2_2873_1[0]));    relay_conn far_2_2873_1_b(.in(far_2_2873_0[1]), .out(far_2_2873_1[1]));
    assign layer_2[833] = far_2_2873_1[0]; 
    assign layer_2[834] = ~layer_1[866] | (layer_1[866] & layer_1[876]); 
    wire [1:0] far_2_2875_0;    relay_conn far_2_2875_0_a(.in(layer_1[184]), .out(far_2_2875_0[0]));    relay_conn far_2_2875_0_b(.in(layer_1[242]), .out(far_2_2875_0[1]));
    assign layer_2[835] = far_2_2875_0[0] & far_2_2875_0[1]; 
    wire [1:0] far_2_2876_0;    relay_conn far_2_2876_0_a(.in(layer_1[320]), .out(far_2_2876_0[0]));    relay_conn far_2_2876_0_b(.in(layer_1[442]), .out(far_2_2876_0[1]));
    wire [1:0] far_2_2876_1;    relay_conn far_2_2876_1_a(.in(far_2_2876_0[0]), .out(far_2_2876_1[0]));    relay_conn far_2_2876_1_b(.in(far_2_2876_0[1]), .out(far_2_2876_1[1]));
    wire [1:0] far_2_2876_2;    relay_conn far_2_2876_2_a(.in(far_2_2876_1[0]), .out(far_2_2876_2[0]));    relay_conn far_2_2876_2_b(.in(far_2_2876_1[1]), .out(far_2_2876_2[1]));
    assign layer_2[836] = ~far_2_2876_2[1] | (far_2_2876_2[0] & far_2_2876_2[1]); 
    wire [1:0] far_2_2877_0;    relay_conn far_2_2877_0_a(.in(layer_1[517]), .out(far_2_2877_0[0]));    relay_conn far_2_2877_0_b(.in(layer_1[617]), .out(far_2_2877_0[1]));
    wire [1:0] far_2_2877_1;    relay_conn far_2_2877_1_a(.in(far_2_2877_0[0]), .out(far_2_2877_1[0]));    relay_conn far_2_2877_1_b(.in(far_2_2877_0[1]), .out(far_2_2877_1[1]));
    wire [1:0] far_2_2877_2;    relay_conn far_2_2877_2_a(.in(far_2_2877_1[0]), .out(far_2_2877_2[0]));    relay_conn far_2_2877_2_b(.in(far_2_2877_1[1]), .out(far_2_2877_2[1]));
    assign layer_2[837] = ~far_2_2877_2[1] | (far_2_2877_2[0] & far_2_2877_2[1]); 
    wire [1:0] far_2_2878_0;    relay_conn far_2_2878_0_a(.in(layer_1[617]), .out(far_2_2878_0[0]));    relay_conn far_2_2878_0_b(.in(layer_1[686]), .out(far_2_2878_0[1]));
    wire [1:0] far_2_2878_1;    relay_conn far_2_2878_1_a(.in(far_2_2878_0[0]), .out(far_2_2878_1[0]));    relay_conn far_2_2878_1_b(.in(far_2_2878_0[1]), .out(far_2_2878_1[1]));
    assign layer_2[838] = far_2_2878_1[0]; 
    wire [1:0] far_2_2879_0;    relay_conn far_2_2879_0_a(.in(layer_1[773]), .out(far_2_2879_0[0]));    relay_conn far_2_2879_0_b(.in(layer_1[852]), .out(far_2_2879_0[1]));
    wire [1:0] far_2_2879_1;    relay_conn far_2_2879_1_a(.in(far_2_2879_0[0]), .out(far_2_2879_1[0]));    relay_conn far_2_2879_1_b(.in(far_2_2879_0[1]), .out(far_2_2879_1[1]));
    assign layer_2[839] = ~far_2_2879_1[0]; 
    assign layer_2[840] = ~(layer_1[991] & layer_1[1018]); 
    wire [1:0] far_2_2881_0;    relay_conn far_2_2881_0_a(.in(layer_1[472]), .out(far_2_2881_0[0]));    relay_conn far_2_2881_0_b(.in(layer_1[533]), .out(far_2_2881_0[1]));
    assign layer_2[841] = ~far_2_2881_0[1] | (far_2_2881_0[0] & far_2_2881_0[1]); 
    assign layer_2[842] = layer_1[72] & ~layer_1[57]; 
    wire [1:0] far_2_2883_0;    relay_conn far_2_2883_0_a(.in(layer_1[564]), .out(far_2_2883_0[0]));    relay_conn far_2_2883_0_b(.in(layer_1[522]), .out(far_2_2883_0[1]));
    assign layer_2[843] = far_2_2883_0[0] & far_2_2883_0[1]; 
    wire [1:0] far_2_2884_0;    relay_conn far_2_2884_0_a(.in(layer_1[127]), .out(far_2_2884_0[0]));    relay_conn far_2_2884_0_b(.in(layer_1[212]), .out(far_2_2884_0[1]));
    wire [1:0] far_2_2884_1;    relay_conn far_2_2884_1_a(.in(far_2_2884_0[0]), .out(far_2_2884_1[0]));    relay_conn far_2_2884_1_b(.in(far_2_2884_0[1]), .out(far_2_2884_1[1]));
    assign layer_2[844] = ~far_2_2884_1[0]; 
    wire [1:0] far_2_2885_0;    relay_conn far_2_2885_0_a(.in(layer_1[871]), .out(far_2_2885_0[0]));    relay_conn far_2_2885_0_b(.in(layer_1[772]), .out(far_2_2885_0[1]));
    wire [1:0] far_2_2885_1;    relay_conn far_2_2885_1_a(.in(far_2_2885_0[0]), .out(far_2_2885_1[0]));    relay_conn far_2_2885_1_b(.in(far_2_2885_0[1]), .out(far_2_2885_1[1]));
    wire [1:0] far_2_2885_2;    relay_conn far_2_2885_2_a(.in(far_2_2885_1[0]), .out(far_2_2885_2[0]));    relay_conn far_2_2885_2_b(.in(far_2_2885_1[1]), .out(far_2_2885_2[1]));
    assign layer_2[845] = far_2_2885_2[0]; 
    assign layer_2[846] = layer_1[765] & layer_1[742]; 
    wire [1:0] far_2_2887_0;    relay_conn far_2_2887_0_a(.in(layer_1[158]), .out(far_2_2887_0[0]));    relay_conn far_2_2887_0_b(.in(layer_1[280]), .out(far_2_2887_0[1]));
    wire [1:0] far_2_2887_1;    relay_conn far_2_2887_1_a(.in(far_2_2887_0[0]), .out(far_2_2887_1[0]));    relay_conn far_2_2887_1_b(.in(far_2_2887_0[1]), .out(far_2_2887_1[1]));
    wire [1:0] far_2_2887_2;    relay_conn far_2_2887_2_a(.in(far_2_2887_1[0]), .out(far_2_2887_2[0]));    relay_conn far_2_2887_2_b(.in(far_2_2887_1[1]), .out(far_2_2887_2[1]));
    assign layer_2[847] = ~far_2_2887_2[0]; 
    wire [1:0] far_2_2888_0;    relay_conn far_2_2888_0_a(.in(layer_1[876]), .out(far_2_2888_0[0]));    relay_conn far_2_2888_0_b(.in(layer_1[935]), .out(far_2_2888_0[1]));
    assign layer_2[848] = far_2_2888_0[0]; 
    wire [1:0] far_2_2889_0;    relay_conn far_2_2889_0_a(.in(layer_1[346]), .out(far_2_2889_0[0]));    relay_conn far_2_2889_0_b(.in(layer_1[284]), .out(far_2_2889_0[1]));
    assign layer_2[849] = far_2_2889_0[0] & ~far_2_2889_0[1]; 
    assign layer_2[850] = ~(layer_1[696] | layer_1[675]); 
    assign layer_2[851] = ~(layer_1[426] ^ layer_1[439]); 
    wire [1:0] far_2_2892_0;    relay_conn far_2_2892_0_a(.in(layer_1[404]), .out(far_2_2892_0[0]));    relay_conn far_2_2892_0_b(.in(layer_1[336]), .out(far_2_2892_0[1]));
    wire [1:0] far_2_2892_1;    relay_conn far_2_2892_1_a(.in(far_2_2892_0[0]), .out(far_2_2892_1[0]));    relay_conn far_2_2892_1_b(.in(far_2_2892_0[1]), .out(far_2_2892_1[1]));
    assign layer_2[852] = far_2_2892_1[1] & ~far_2_2892_1[0]; 
    wire [1:0] far_2_2893_0;    relay_conn far_2_2893_0_a(.in(layer_1[303]), .out(far_2_2893_0[0]));    relay_conn far_2_2893_0_b(.in(layer_1[401]), .out(far_2_2893_0[1]));
    wire [1:0] far_2_2893_1;    relay_conn far_2_2893_1_a(.in(far_2_2893_0[0]), .out(far_2_2893_1[0]));    relay_conn far_2_2893_1_b(.in(far_2_2893_0[1]), .out(far_2_2893_1[1]));
    wire [1:0] far_2_2893_2;    relay_conn far_2_2893_2_a(.in(far_2_2893_1[0]), .out(far_2_2893_2[0]));    relay_conn far_2_2893_2_b(.in(far_2_2893_1[1]), .out(far_2_2893_2[1]));
    assign layer_2[853] = far_2_2893_2[0] & ~far_2_2893_2[1]; 
    assign layer_2[854] = ~layer_1[123]; 
    wire [1:0] far_2_2895_0;    relay_conn far_2_2895_0_a(.in(layer_1[196]), .out(far_2_2895_0[0]));    relay_conn far_2_2895_0_b(.in(layer_1[296]), .out(far_2_2895_0[1]));
    wire [1:0] far_2_2895_1;    relay_conn far_2_2895_1_a(.in(far_2_2895_0[0]), .out(far_2_2895_1[0]));    relay_conn far_2_2895_1_b(.in(far_2_2895_0[1]), .out(far_2_2895_1[1]));
    wire [1:0] far_2_2895_2;    relay_conn far_2_2895_2_a(.in(far_2_2895_1[0]), .out(far_2_2895_2[0]));    relay_conn far_2_2895_2_b(.in(far_2_2895_1[1]), .out(far_2_2895_2[1]));
    assign layer_2[855] = far_2_2895_2[0] | far_2_2895_2[1]; 
    assign layer_2[856] = ~(layer_1[768] & layer_1[795]); 
    wire [1:0] far_2_2897_0;    relay_conn far_2_2897_0_a(.in(layer_1[200]), .out(far_2_2897_0[0]));    relay_conn far_2_2897_0_b(.in(layer_1[235]), .out(far_2_2897_0[1]));
    assign layer_2[857] = far_2_2897_0[0] & far_2_2897_0[1]; 
    wire [1:0] far_2_2898_0;    relay_conn far_2_2898_0_a(.in(layer_1[781]), .out(far_2_2898_0[0]));    relay_conn far_2_2898_0_b(.in(layer_1[743]), .out(far_2_2898_0[1]));
    assign layer_2[858] = far_2_2898_0[0] & ~far_2_2898_0[1]; 
    wire [1:0] far_2_2899_0;    relay_conn far_2_2899_0_a(.in(layer_1[118]), .out(far_2_2899_0[0]));    relay_conn far_2_2899_0_b(.in(layer_1[171]), .out(far_2_2899_0[1]));
    assign layer_2[859] = ~(far_2_2899_0[0] | far_2_2899_0[1]); 
    wire [1:0] far_2_2900_0;    relay_conn far_2_2900_0_a(.in(layer_1[327]), .out(far_2_2900_0[0]));    relay_conn far_2_2900_0_b(.in(layer_1[261]), .out(far_2_2900_0[1]));
    wire [1:0] far_2_2900_1;    relay_conn far_2_2900_1_a(.in(far_2_2900_0[0]), .out(far_2_2900_1[0]));    relay_conn far_2_2900_1_b(.in(far_2_2900_0[1]), .out(far_2_2900_1[1]));
    assign layer_2[860] = far_2_2900_1[0] & far_2_2900_1[1]; 
    wire [1:0] far_2_2901_0;    relay_conn far_2_2901_0_a(.in(layer_1[288]), .out(far_2_2901_0[0]));    relay_conn far_2_2901_0_b(.in(layer_1[212]), .out(far_2_2901_0[1]));
    wire [1:0] far_2_2901_1;    relay_conn far_2_2901_1_a(.in(far_2_2901_0[0]), .out(far_2_2901_1[0]));    relay_conn far_2_2901_1_b(.in(far_2_2901_0[1]), .out(far_2_2901_1[1]));
    assign layer_2[861] = ~far_2_2901_1[1] | (far_2_2901_1[0] & far_2_2901_1[1]); 
    wire [1:0] far_2_2902_0;    relay_conn far_2_2902_0_a(.in(layer_1[273]), .out(far_2_2902_0[0]));    relay_conn far_2_2902_0_b(.in(layer_1[401]), .out(far_2_2902_0[1]));
    wire [1:0] far_2_2902_1;    relay_conn far_2_2902_1_a(.in(far_2_2902_0[0]), .out(far_2_2902_1[0]));    relay_conn far_2_2902_1_b(.in(far_2_2902_0[1]), .out(far_2_2902_1[1]));
    wire [1:0] far_2_2902_2;    relay_conn far_2_2902_2_a(.in(far_2_2902_1[0]), .out(far_2_2902_2[0]));    relay_conn far_2_2902_2_b(.in(far_2_2902_1[1]), .out(far_2_2902_2[1]));
    wire [1:0] far_2_2902_3;    relay_conn far_2_2902_3_a(.in(far_2_2902_2[0]), .out(far_2_2902_3[0]));    relay_conn far_2_2902_3_b(.in(far_2_2902_2[1]), .out(far_2_2902_3[1]));
    assign layer_2[862] = ~(far_2_2902_3[0] & far_2_2902_3[1]); 
    wire [1:0] far_2_2903_0;    relay_conn far_2_2903_0_a(.in(layer_1[106]), .out(far_2_2903_0[0]));    relay_conn far_2_2903_0_b(.in(layer_1[65]), .out(far_2_2903_0[1]));
    assign layer_2[863] = ~far_2_2903_0[1] | (far_2_2903_0[0] & far_2_2903_0[1]); 
    assign layer_2[864] = layer_1[962] & ~layer_1[964]; 
    assign layer_2[865] = layer_1[967] & layer_1[946]; 
    wire [1:0] far_2_2906_0;    relay_conn far_2_2906_0_a(.in(layer_1[213]), .out(far_2_2906_0[0]));    relay_conn far_2_2906_0_b(.in(layer_1[326]), .out(far_2_2906_0[1]));
    wire [1:0] far_2_2906_1;    relay_conn far_2_2906_1_a(.in(far_2_2906_0[0]), .out(far_2_2906_1[0]));    relay_conn far_2_2906_1_b(.in(far_2_2906_0[1]), .out(far_2_2906_1[1]));
    wire [1:0] far_2_2906_2;    relay_conn far_2_2906_2_a(.in(far_2_2906_1[0]), .out(far_2_2906_2[0]));    relay_conn far_2_2906_2_b(.in(far_2_2906_1[1]), .out(far_2_2906_2[1]));
    assign layer_2[866] = ~far_2_2906_2[1]; 
    wire [1:0] far_2_2907_0;    relay_conn far_2_2907_0_a(.in(layer_1[367]), .out(far_2_2907_0[0]));    relay_conn far_2_2907_0_b(.in(layer_1[308]), .out(far_2_2907_0[1]));
    assign layer_2[867] = far_2_2907_0[0] & far_2_2907_0[1]; 
    wire [1:0] far_2_2908_0;    relay_conn far_2_2908_0_a(.in(layer_1[281]), .out(far_2_2908_0[0]));    relay_conn far_2_2908_0_b(.in(layer_1[314]), .out(far_2_2908_0[1]));
    assign layer_2[868] = far_2_2908_0[0] | far_2_2908_0[1]; 
    assign layer_2[869] = layer_1[173] ^ layer_1[171]; 
    wire [1:0] far_2_2910_0;    relay_conn far_2_2910_0_a(.in(layer_1[127]), .out(far_2_2910_0[0]));    relay_conn far_2_2910_0_b(.in(layer_1[169]), .out(far_2_2910_0[1]));
    assign layer_2[870] = ~far_2_2910_0[1] | (far_2_2910_0[0] & far_2_2910_0[1]); 
    assign layer_2[871] = ~(layer_1[52] & layer_1[58]); 
    wire [1:0] far_2_2912_0;    relay_conn far_2_2912_0_a(.in(layer_1[879]), .out(far_2_2912_0[0]));    relay_conn far_2_2912_0_b(.in(layer_1[781]), .out(far_2_2912_0[1]));
    wire [1:0] far_2_2912_1;    relay_conn far_2_2912_1_a(.in(far_2_2912_0[0]), .out(far_2_2912_1[0]));    relay_conn far_2_2912_1_b(.in(far_2_2912_0[1]), .out(far_2_2912_1[1]));
    wire [1:0] far_2_2912_2;    relay_conn far_2_2912_2_a(.in(far_2_2912_1[0]), .out(far_2_2912_2[0]));    relay_conn far_2_2912_2_b(.in(far_2_2912_1[1]), .out(far_2_2912_2[1]));
    assign layer_2[872] = far_2_2912_2[0] & far_2_2912_2[1]; 
    wire [1:0] far_2_2913_0;    relay_conn far_2_2913_0_a(.in(layer_1[442]), .out(far_2_2913_0[0]));    relay_conn far_2_2913_0_b(.in(layer_1[553]), .out(far_2_2913_0[1]));
    wire [1:0] far_2_2913_1;    relay_conn far_2_2913_1_a(.in(far_2_2913_0[0]), .out(far_2_2913_1[0]));    relay_conn far_2_2913_1_b(.in(far_2_2913_0[1]), .out(far_2_2913_1[1]));
    wire [1:0] far_2_2913_2;    relay_conn far_2_2913_2_a(.in(far_2_2913_1[0]), .out(far_2_2913_2[0]));    relay_conn far_2_2913_2_b(.in(far_2_2913_1[1]), .out(far_2_2913_2[1]));
    assign layer_2[873] = far_2_2913_2[0]; 
    wire [1:0] far_2_2914_0;    relay_conn far_2_2914_0_a(.in(layer_1[55]), .out(far_2_2914_0[0]));    relay_conn far_2_2914_0_b(.in(layer_1[115]), .out(far_2_2914_0[1]));
    assign layer_2[874] = ~far_2_2914_0[1]; 
    assign layer_2[875] = layer_1[533]; 
    wire [1:0] far_2_2916_0;    relay_conn far_2_2916_0_a(.in(layer_1[716]), .out(far_2_2916_0[0]));    relay_conn far_2_2916_0_b(.in(layer_1[682]), .out(far_2_2916_0[1]));
    assign layer_2[876] = ~(far_2_2916_0[0] & far_2_2916_0[1]); 
    wire [1:0] far_2_2917_0;    relay_conn far_2_2917_0_a(.in(layer_1[562]), .out(far_2_2917_0[0]));    relay_conn far_2_2917_0_b(.in(layer_1[486]), .out(far_2_2917_0[1]));
    wire [1:0] far_2_2917_1;    relay_conn far_2_2917_1_a(.in(far_2_2917_0[0]), .out(far_2_2917_1[0]));    relay_conn far_2_2917_1_b(.in(far_2_2917_0[1]), .out(far_2_2917_1[1]));
    assign layer_2[877] = ~far_2_2917_1[1] | (far_2_2917_1[0] & far_2_2917_1[1]); 
    assign layer_2[878] = layer_1[955] & ~layer_1[926]; 
    wire [1:0] far_2_2919_0;    relay_conn far_2_2919_0_a(.in(layer_1[156]), .out(far_2_2919_0[0]));    relay_conn far_2_2919_0_b(.in(layer_1[46]), .out(far_2_2919_0[1]));
    wire [1:0] far_2_2919_1;    relay_conn far_2_2919_1_a(.in(far_2_2919_0[0]), .out(far_2_2919_1[0]));    relay_conn far_2_2919_1_b(.in(far_2_2919_0[1]), .out(far_2_2919_1[1]));
    wire [1:0] far_2_2919_2;    relay_conn far_2_2919_2_a(.in(far_2_2919_1[0]), .out(far_2_2919_2[0]));    relay_conn far_2_2919_2_b(.in(far_2_2919_1[1]), .out(far_2_2919_2[1]));
    assign layer_2[879] = far_2_2919_2[0] & far_2_2919_2[1]; 
    wire [1:0] far_2_2920_0;    relay_conn far_2_2920_0_a(.in(layer_1[604]), .out(far_2_2920_0[0]));    relay_conn far_2_2920_0_b(.in(layer_1[670]), .out(far_2_2920_0[1]));
    wire [1:0] far_2_2920_1;    relay_conn far_2_2920_1_a(.in(far_2_2920_0[0]), .out(far_2_2920_1[0]));    relay_conn far_2_2920_1_b(.in(far_2_2920_0[1]), .out(far_2_2920_1[1]));
    assign layer_2[880] = far_2_2920_1[0] & ~far_2_2920_1[1]; 
    wire [1:0] far_2_2921_0;    relay_conn far_2_2921_0_a(.in(layer_1[626]), .out(far_2_2921_0[0]));    relay_conn far_2_2921_0_b(.in(layer_1[562]), .out(far_2_2921_0[1]));
    wire [1:0] far_2_2921_1;    relay_conn far_2_2921_1_a(.in(far_2_2921_0[0]), .out(far_2_2921_1[0]));    relay_conn far_2_2921_1_b(.in(far_2_2921_0[1]), .out(far_2_2921_1[1]));
    assign layer_2[881] = far_2_2921_1[0] & far_2_2921_1[1]; 
    wire [1:0] far_2_2922_0;    relay_conn far_2_2922_0_a(.in(layer_1[1018]), .out(far_2_2922_0[0]));    relay_conn far_2_2922_0_b(.in(layer_1[909]), .out(far_2_2922_0[1]));
    wire [1:0] far_2_2922_1;    relay_conn far_2_2922_1_a(.in(far_2_2922_0[0]), .out(far_2_2922_1[0]));    relay_conn far_2_2922_1_b(.in(far_2_2922_0[1]), .out(far_2_2922_1[1]));
    wire [1:0] far_2_2922_2;    relay_conn far_2_2922_2_a(.in(far_2_2922_1[0]), .out(far_2_2922_2[0]));    relay_conn far_2_2922_2_b(.in(far_2_2922_1[1]), .out(far_2_2922_2[1]));
    assign layer_2[882] = ~far_2_2922_2[0]; 
    assign layer_2[883] = ~(layer_1[561] & layer_1[559]); 
    wire [1:0] far_2_2924_0;    relay_conn far_2_2924_0_a(.in(layer_1[385]), .out(far_2_2924_0[0]));    relay_conn far_2_2924_0_b(.in(layer_1[296]), .out(far_2_2924_0[1]));
    wire [1:0] far_2_2924_1;    relay_conn far_2_2924_1_a(.in(far_2_2924_0[0]), .out(far_2_2924_1[0]));    relay_conn far_2_2924_1_b(.in(far_2_2924_0[1]), .out(far_2_2924_1[1]));
    assign layer_2[884] = far_2_2924_1[0]; 
    wire [1:0] far_2_2925_0;    relay_conn far_2_2925_0_a(.in(layer_1[557]), .out(far_2_2925_0[0]));    relay_conn far_2_2925_0_b(.in(layer_1[596]), .out(far_2_2925_0[1]));
    assign layer_2[885] = ~(far_2_2925_0[0] | far_2_2925_0[1]); 
    wire [1:0] far_2_2926_0;    relay_conn far_2_2926_0_a(.in(layer_1[825]), .out(far_2_2926_0[0]));    relay_conn far_2_2926_0_b(.in(layer_1[769]), .out(far_2_2926_0[1]));
    assign layer_2[886] = ~(far_2_2926_0[0] | far_2_2926_0[1]); 
    wire [1:0] far_2_2927_0;    relay_conn far_2_2927_0_a(.in(layer_1[391]), .out(far_2_2927_0[0]));    relay_conn far_2_2927_0_b(.in(layer_1[352]), .out(far_2_2927_0[1]));
    assign layer_2[887] = ~far_2_2927_0[1] | (far_2_2927_0[0] & far_2_2927_0[1]); 
    wire [1:0] far_2_2928_0;    relay_conn far_2_2928_0_a(.in(layer_1[793]), .out(far_2_2928_0[0]));    relay_conn far_2_2928_0_b(.in(layer_1[747]), .out(far_2_2928_0[1]));
    assign layer_2[888] = far_2_2928_0[1] & ~far_2_2928_0[0]; 
    wire [1:0] far_2_2929_0;    relay_conn far_2_2929_0_a(.in(layer_1[288]), .out(far_2_2929_0[0]));    relay_conn far_2_2929_0_b(.in(layer_1[163]), .out(far_2_2929_0[1]));
    wire [1:0] far_2_2929_1;    relay_conn far_2_2929_1_a(.in(far_2_2929_0[0]), .out(far_2_2929_1[0]));    relay_conn far_2_2929_1_b(.in(far_2_2929_0[1]), .out(far_2_2929_1[1]));
    wire [1:0] far_2_2929_2;    relay_conn far_2_2929_2_a(.in(far_2_2929_1[0]), .out(far_2_2929_2[0]));    relay_conn far_2_2929_2_b(.in(far_2_2929_1[1]), .out(far_2_2929_2[1]));
    assign layer_2[889] = far_2_2929_2[1] & ~far_2_2929_2[0]; 
    wire [1:0] far_2_2930_0;    relay_conn far_2_2930_0_a(.in(layer_1[846]), .out(far_2_2930_0[0]));    relay_conn far_2_2930_0_b(.in(layer_1[896]), .out(far_2_2930_0[1]));
    assign layer_2[890] = ~far_2_2930_0[0]; 
    wire [1:0] far_2_2931_0;    relay_conn far_2_2931_0_a(.in(layer_1[232]), .out(far_2_2931_0[0]));    relay_conn far_2_2931_0_b(.in(layer_1[196]), .out(far_2_2931_0[1]));
    assign layer_2[891] = far_2_2931_0[0]; 
    assign layer_2[892] = ~(layer_1[256] | layer_1[229]); 
    assign layer_2[893] = ~layer_1[875] | (layer_1[897] & layer_1[875]); 
    wire [1:0] far_2_2934_0;    relay_conn far_2_2934_0_a(.in(layer_1[177]), .out(far_2_2934_0[0]));    relay_conn far_2_2934_0_b(.in(layer_1[115]), .out(far_2_2934_0[1]));
    assign layer_2[894] = ~far_2_2934_0[0]; 
    assign layer_2[895] = layer_1[248]; 
    wire [1:0] far_2_2936_0;    relay_conn far_2_2936_0_a(.in(layer_1[336]), .out(far_2_2936_0[0]));    relay_conn far_2_2936_0_b(.in(layer_1[396]), .out(far_2_2936_0[1]));
    assign layer_2[896] = ~far_2_2936_0[1] | (far_2_2936_0[0] & far_2_2936_0[1]); 
    wire [1:0] far_2_2937_0;    relay_conn far_2_2937_0_a(.in(layer_1[212]), .out(far_2_2937_0[0]));    relay_conn far_2_2937_0_b(.in(layer_1[280]), .out(far_2_2937_0[1]));
    wire [1:0] far_2_2937_1;    relay_conn far_2_2937_1_a(.in(far_2_2937_0[0]), .out(far_2_2937_1[0]));    relay_conn far_2_2937_1_b(.in(far_2_2937_0[1]), .out(far_2_2937_1[1]));
    assign layer_2[897] = ~far_2_2937_1[0]; 
    assign layer_2[898] = layer_1[674] & ~layer_1[694]; 
    assign layer_2[899] = layer_1[312] & ~layer_1[320]; 
    wire [1:0] far_2_2940_0;    relay_conn far_2_2940_0_a(.in(layer_1[987]), .out(far_2_2940_0[0]));    relay_conn far_2_2940_0_b(.in(layer_1[955]), .out(far_2_2940_0[1]));
    assign layer_2[900] = ~far_2_2940_0[1] | (far_2_2940_0[0] & far_2_2940_0[1]); 
    wire [1:0] far_2_2941_0;    relay_conn far_2_2941_0_a(.in(layer_1[977]), .out(far_2_2941_0[0]));    relay_conn far_2_2941_0_b(.in(layer_1[903]), .out(far_2_2941_0[1]));
    wire [1:0] far_2_2941_1;    relay_conn far_2_2941_1_a(.in(far_2_2941_0[0]), .out(far_2_2941_1[0]));    relay_conn far_2_2941_1_b(.in(far_2_2941_0[1]), .out(far_2_2941_1[1]));
    assign layer_2[901] = ~far_2_2941_1[0] | (far_2_2941_1[0] & far_2_2941_1[1]); 
    wire [1:0] far_2_2942_0;    relay_conn far_2_2942_0_a(.in(layer_1[352]), .out(far_2_2942_0[0]));    relay_conn far_2_2942_0_b(.in(layer_1[224]), .out(far_2_2942_0[1]));
    wire [1:0] far_2_2942_1;    relay_conn far_2_2942_1_a(.in(far_2_2942_0[0]), .out(far_2_2942_1[0]));    relay_conn far_2_2942_1_b(.in(far_2_2942_0[1]), .out(far_2_2942_1[1]));
    wire [1:0] far_2_2942_2;    relay_conn far_2_2942_2_a(.in(far_2_2942_1[0]), .out(far_2_2942_2[0]));    relay_conn far_2_2942_2_b(.in(far_2_2942_1[1]), .out(far_2_2942_2[1]));
    wire [1:0] far_2_2942_3;    relay_conn far_2_2942_3_a(.in(far_2_2942_2[0]), .out(far_2_2942_3[0]));    relay_conn far_2_2942_3_b(.in(far_2_2942_2[1]), .out(far_2_2942_3[1]));
    assign layer_2[902] = far_2_2942_3[0] & ~far_2_2942_3[1]; 
    wire [1:0] far_2_2943_0;    relay_conn far_2_2943_0_a(.in(layer_1[227]), .out(far_2_2943_0[0]));    relay_conn far_2_2943_0_b(.in(layer_1[115]), .out(far_2_2943_0[1]));
    wire [1:0] far_2_2943_1;    relay_conn far_2_2943_1_a(.in(far_2_2943_0[0]), .out(far_2_2943_1[0]));    relay_conn far_2_2943_1_b(.in(far_2_2943_0[1]), .out(far_2_2943_1[1]));
    wire [1:0] far_2_2943_2;    relay_conn far_2_2943_2_a(.in(far_2_2943_1[0]), .out(far_2_2943_2[0]));    relay_conn far_2_2943_2_b(.in(far_2_2943_1[1]), .out(far_2_2943_2[1]));
    assign layer_2[903] = far_2_2943_2[1]; 
    wire [1:0] far_2_2944_0;    relay_conn far_2_2944_0_a(.in(layer_1[90]), .out(far_2_2944_0[0]));    relay_conn far_2_2944_0_b(.in(layer_1[207]), .out(far_2_2944_0[1]));
    wire [1:0] far_2_2944_1;    relay_conn far_2_2944_1_a(.in(far_2_2944_0[0]), .out(far_2_2944_1[0]));    relay_conn far_2_2944_1_b(.in(far_2_2944_0[1]), .out(far_2_2944_1[1]));
    wire [1:0] far_2_2944_2;    relay_conn far_2_2944_2_a(.in(far_2_2944_1[0]), .out(far_2_2944_2[0]));    relay_conn far_2_2944_2_b(.in(far_2_2944_1[1]), .out(far_2_2944_2[1]));
    assign layer_2[904] = ~(far_2_2944_2[0] & far_2_2944_2[1]); 
    wire [1:0] far_2_2945_0;    relay_conn far_2_2945_0_a(.in(layer_1[363]), .out(far_2_2945_0[0]));    relay_conn far_2_2945_0_b(.in(layer_1[324]), .out(far_2_2945_0[1]));
    assign layer_2[905] = ~far_2_2945_0[0] | (far_2_2945_0[0] & far_2_2945_0[1]); 
    wire [1:0] far_2_2946_0;    relay_conn far_2_2946_0_a(.in(layer_1[59]), .out(far_2_2946_0[0]));    relay_conn far_2_2946_0_b(.in(layer_1[133]), .out(far_2_2946_0[1]));
    wire [1:0] far_2_2946_1;    relay_conn far_2_2946_1_a(.in(far_2_2946_0[0]), .out(far_2_2946_1[0]));    relay_conn far_2_2946_1_b(.in(far_2_2946_0[1]), .out(far_2_2946_1[1]));
    assign layer_2[906] = ~(far_2_2946_1[0] & far_2_2946_1[1]); 
    assign layer_2[907] = ~layer_1[564] | (layer_1[554] & layer_1[564]); 
    assign layer_2[908] = ~layer_1[84]; 
    wire [1:0] far_2_2949_0;    relay_conn far_2_2949_0_a(.in(layer_1[688]), .out(far_2_2949_0[0]));    relay_conn far_2_2949_0_b(.in(layer_1[804]), .out(far_2_2949_0[1]));
    wire [1:0] far_2_2949_1;    relay_conn far_2_2949_1_a(.in(far_2_2949_0[0]), .out(far_2_2949_1[0]));    relay_conn far_2_2949_1_b(.in(far_2_2949_0[1]), .out(far_2_2949_1[1]));
    wire [1:0] far_2_2949_2;    relay_conn far_2_2949_2_a(.in(far_2_2949_1[0]), .out(far_2_2949_2[0]));    relay_conn far_2_2949_2_b(.in(far_2_2949_1[1]), .out(far_2_2949_2[1]));
    assign layer_2[909] = far_2_2949_2[0] ^ far_2_2949_2[1]; 
    wire [1:0] far_2_2950_0;    relay_conn far_2_2950_0_a(.in(layer_1[57]), .out(far_2_2950_0[0]));    relay_conn far_2_2950_0_b(.in(layer_1[137]), .out(far_2_2950_0[1]));
    wire [1:0] far_2_2950_1;    relay_conn far_2_2950_1_a(.in(far_2_2950_0[0]), .out(far_2_2950_1[0]));    relay_conn far_2_2950_1_b(.in(far_2_2950_0[1]), .out(far_2_2950_1[1]));
    assign layer_2[910] = far_2_2950_1[0] & far_2_2950_1[1]; 
    wire [1:0] far_2_2951_0;    relay_conn far_2_2951_0_a(.in(layer_1[781]), .out(far_2_2951_0[0]));    relay_conn far_2_2951_0_b(.in(layer_1[709]), .out(far_2_2951_0[1]));
    wire [1:0] far_2_2951_1;    relay_conn far_2_2951_1_a(.in(far_2_2951_0[0]), .out(far_2_2951_1[0]));    relay_conn far_2_2951_1_b(.in(far_2_2951_0[1]), .out(far_2_2951_1[1]));
    assign layer_2[911] = ~far_2_2951_1[0] | (far_2_2951_1[0] & far_2_2951_1[1]); 
    wire [1:0] far_2_2952_0;    relay_conn far_2_2952_0_a(.in(layer_1[599]), .out(far_2_2952_0[0]));    relay_conn far_2_2952_0_b(.in(layer_1[717]), .out(far_2_2952_0[1]));
    wire [1:0] far_2_2952_1;    relay_conn far_2_2952_1_a(.in(far_2_2952_0[0]), .out(far_2_2952_1[0]));    relay_conn far_2_2952_1_b(.in(far_2_2952_0[1]), .out(far_2_2952_1[1]));
    wire [1:0] far_2_2952_2;    relay_conn far_2_2952_2_a(.in(far_2_2952_1[0]), .out(far_2_2952_2[0]));    relay_conn far_2_2952_2_b(.in(far_2_2952_1[1]), .out(far_2_2952_2[1]));
    assign layer_2[912] = far_2_2952_2[0] & far_2_2952_2[1]; 
    wire [1:0] far_2_2953_0;    relay_conn far_2_2953_0_a(.in(layer_1[593]), .out(far_2_2953_0[0]));    relay_conn far_2_2953_0_b(.in(layer_1[648]), .out(far_2_2953_0[1]));
    assign layer_2[913] = far_2_2953_0[0] | far_2_2953_0[1]; 
    assign layer_2[914] = layer_1[851] | layer_1[867]; 
    wire [1:0] far_2_2955_0;    relay_conn far_2_2955_0_a(.in(layer_1[623]), .out(far_2_2955_0[0]));    relay_conn far_2_2955_0_b(.in(layer_1[577]), .out(far_2_2955_0[1]));
    assign layer_2[915] = far_2_2955_0[1]; 
    wire [1:0] far_2_2956_0;    relay_conn far_2_2956_0_a(.in(layer_1[740]), .out(far_2_2956_0[0]));    relay_conn far_2_2956_0_b(.in(layer_1[796]), .out(far_2_2956_0[1]));
    assign layer_2[916] = ~(far_2_2956_0[0] & far_2_2956_0[1]); 
    wire [1:0] far_2_2957_0;    relay_conn far_2_2957_0_a(.in(layer_1[316]), .out(far_2_2957_0[0]));    relay_conn far_2_2957_0_b(.in(layer_1[357]), .out(far_2_2957_0[1]));
    assign layer_2[917] = ~(far_2_2957_0[0] ^ far_2_2957_0[1]); 
    wire [1:0] far_2_2958_0;    relay_conn far_2_2958_0_a(.in(layer_1[180]), .out(far_2_2958_0[0]));    relay_conn far_2_2958_0_b(.in(layer_1[73]), .out(far_2_2958_0[1]));
    wire [1:0] far_2_2958_1;    relay_conn far_2_2958_1_a(.in(far_2_2958_0[0]), .out(far_2_2958_1[0]));    relay_conn far_2_2958_1_b(.in(far_2_2958_0[1]), .out(far_2_2958_1[1]));
    wire [1:0] far_2_2958_2;    relay_conn far_2_2958_2_a(.in(far_2_2958_1[0]), .out(far_2_2958_2[0]));    relay_conn far_2_2958_2_b(.in(far_2_2958_1[1]), .out(far_2_2958_2[1]));
    assign layer_2[918] = far_2_2958_2[1] & ~far_2_2958_2[0]; 
    wire [1:0] far_2_2959_0;    relay_conn far_2_2959_0_a(.in(layer_1[676]), .out(far_2_2959_0[0]));    relay_conn far_2_2959_0_b(.in(layer_1[615]), .out(far_2_2959_0[1]));
    assign layer_2[919] = far_2_2959_0[0] & far_2_2959_0[1]; 
    wire [1:0] far_2_2960_0;    relay_conn far_2_2960_0_a(.in(layer_1[669]), .out(far_2_2960_0[0]));    relay_conn far_2_2960_0_b(.in(layer_1[619]), .out(far_2_2960_0[1]));
    assign layer_2[920] = ~far_2_2960_0[1] | (far_2_2960_0[0] & far_2_2960_0[1]); 
    wire [1:0] far_2_2961_0;    relay_conn far_2_2961_0_a(.in(layer_1[1]), .out(far_2_2961_0[0]));    relay_conn far_2_2961_0_b(.in(layer_1[125]), .out(far_2_2961_0[1]));
    wire [1:0] far_2_2961_1;    relay_conn far_2_2961_1_a(.in(far_2_2961_0[0]), .out(far_2_2961_1[0]));    relay_conn far_2_2961_1_b(.in(far_2_2961_0[1]), .out(far_2_2961_1[1]));
    wire [1:0] far_2_2961_2;    relay_conn far_2_2961_2_a(.in(far_2_2961_1[0]), .out(far_2_2961_2[0]));    relay_conn far_2_2961_2_b(.in(far_2_2961_1[1]), .out(far_2_2961_2[1]));
    assign layer_2[921] = ~(far_2_2961_2[0] & far_2_2961_2[1]); 
    wire [1:0] far_2_2962_0;    relay_conn far_2_2962_0_a(.in(layer_1[158]), .out(far_2_2962_0[0]));    relay_conn far_2_2962_0_b(.in(layer_1[232]), .out(far_2_2962_0[1]));
    wire [1:0] far_2_2962_1;    relay_conn far_2_2962_1_a(.in(far_2_2962_0[0]), .out(far_2_2962_1[0]));    relay_conn far_2_2962_1_b(.in(far_2_2962_0[1]), .out(far_2_2962_1[1]));
    assign layer_2[922] = ~(far_2_2962_1[0] | far_2_2962_1[1]); 
    wire [1:0] far_2_2963_0;    relay_conn far_2_2963_0_a(.in(layer_1[884]), .out(far_2_2963_0[0]));    relay_conn far_2_2963_0_b(.in(layer_1[987]), .out(far_2_2963_0[1]));
    wire [1:0] far_2_2963_1;    relay_conn far_2_2963_1_a(.in(far_2_2963_0[0]), .out(far_2_2963_1[0]));    relay_conn far_2_2963_1_b(.in(far_2_2963_0[1]), .out(far_2_2963_1[1]));
    wire [1:0] far_2_2963_2;    relay_conn far_2_2963_2_a(.in(far_2_2963_1[0]), .out(far_2_2963_2[0]));    relay_conn far_2_2963_2_b(.in(far_2_2963_1[1]), .out(far_2_2963_2[1]));
    assign layer_2[923] = ~far_2_2963_2[0] | (far_2_2963_2[0] & far_2_2963_2[1]); 
    assign layer_2[924] = layer_1[533] ^ layer_1[516]; 
    wire [1:0] far_2_2965_0;    relay_conn far_2_2965_0_a(.in(layer_1[598]), .out(far_2_2965_0[0]));    relay_conn far_2_2965_0_b(.in(layer_1[514]), .out(far_2_2965_0[1]));
    wire [1:0] far_2_2965_1;    relay_conn far_2_2965_1_a(.in(far_2_2965_0[0]), .out(far_2_2965_1[0]));    relay_conn far_2_2965_1_b(.in(far_2_2965_0[1]), .out(far_2_2965_1[1]));
    assign layer_2[925] = ~(far_2_2965_1[0] | far_2_2965_1[1]); 
    assign layer_2[926] = layer_1[597]; 
    assign layer_2[927] = ~(layer_1[428] & layer_1[406]); 
    assign layer_2[928] = layer_1[232]; 
    assign layer_2[929] = layer_1[451] & layer_1[422]; 
    wire [1:0] far_2_2970_0;    relay_conn far_2_2970_0_a(.in(layer_1[393]), .out(far_2_2970_0[0]));    relay_conn far_2_2970_0_b(.in(layer_1[456]), .out(far_2_2970_0[1]));
    assign layer_2[930] = ~far_2_2970_0[0] | (far_2_2970_0[0] & far_2_2970_0[1]); 
    assign layer_2[931] = layer_1[518]; 
    assign layer_2[932] = ~layer_1[558] | (layer_1[558] & layer_1[561]); 
    wire [1:0] far_2_2973_0;    relay_conn far_2_2973_0_a(.in(layer_1[430]), .out(far_2_2973_0[0]));    relay_conn far_2_2973_0_b(.in(layer_1[373]), .out(far_2_2973_0[1]));
    assign layer_2[933] = far_2_2973_0[0] & far_2_2973_0[1]; 
    wire [1:0] far_2_2974_0;    relay_conn far_2_2974_0_a(.in(layer_1[317]), .out(far_2_2974_0[0]));    relay_conn far_2_2974_0_b(.in(layer_1[284]), .out(far_2_2974_0[1]));
    assign layer_2[934] = ~far_2_2974_0[0]; 
    assign layer_2[935] = ~layer_1[780] | (layer_1[794] & layer_1[780]); 
    wire [1:0] far_2_2976_0;    relay_conn far_2_2976_0_a(.in(layer_1[460]), .out(far_2_2976_0[0]));    relay_conn far_2_2976_0_b(.in(layer_1[534]), .out(far_2_2976_0[1]));
    wire [1:0] far_2_2976_1;    relay_conn far_2_2976_1_a(.in(far_2_2976_0[0]), .out(far_2_2976_1[0]));    relay_conn far_2_2976_1_b(.in(far_2_2976_0[1]), .out(far_2_2976_1[1]));
    assign layer_2[936] = far_2_2976_1[0]; 
    wire [1:0] far_2_2977_0;    relay_conn far_2_2977_0_a(.in(layer_1[396]), .out(far_2_2977_0[0]));    relay_conn far_2_2977_0_b(.in(layer_1[459]), .out(far_2_2977_0[1]));
    assign layer_2[937] = ~far_2_2977_0[0] | (far_2_2977_0[0] & far_2_2977_0[1]); 
    wire [1:0] far_2_2978_0;    relay_conn far_2_2978_0_a(.in(layer_1[408]), .out(far_2_2978_0[0]));    relay_conn far_2_2978_0_b(.in(layer_1[517]), .out(far_2_2978_0[1]));
    wire [1:0] far_2_2978_1;    relay_conn far_2_2978_1_a(.in(far_2_2978_0[0]), .out(far_2_2978_1[0]));    relay_conn far_2_2978_1_b(.in(far_2_2978_0[1]), .out(far_2_2978_1[1]));
    wire [1:0] far_2_2978_2;    relay_conn far_2_2978_2_a(.in(far_2_2978_1[0]), .out(far_2_2978_2[0]));    relay_conn far_2_2978_2_b(.in(far_2_2978_1[1]), .out(far_2_2978_2[1]));
    assign layer_2[938] = far_2_2978_2[1]; 
    wire [1:0] far_2_2979_0;    relay_conn far_2_2979_0_a(.in(layer_1[452]), .out(far_2_2979_0[0]));    relay_conn far_2_2979_0_b(.in(layer_1[358]), .out(far_2_2979_0[1]));
    wire [1:0] far_2_2979_1;    relay_conn far_2_2979_1_a(.in(far_2_2979_0[0]), .out(far_2_2979_1[0]));    relay_conn far_2_2979_1_b(.in(far_2_2979_0[1]), .out(far_2_2979_1[1]));
    assign layer_2[939] = far_2_2979_1[0] & far_2_2979_1[1]; 
    wire [1:0] far_2_2980_0;    relay_conn far_2_2980_0_a(.in(layer_1[537]), .out(far_2_2980_0[0]));    relay_conn far_2_2980_0_b(.in(layer_1[455]), .out(far_2_2980_0[1]));
    wire [1:0] far_2_2980_1;    relay_conn far_2_2980_1_a(.in(far_2_2980_0[0]), .out(far_2_2980_1[0]));    relay_conn far_2_2980_1_b(.in(far_2_2980_0[1]), .out(far_2_2980_1[1]));
    assign layer_2[940] = far_2_2980_1[0] | far_2_2980_1[1]; 
    wire [1:0] far_2_2981_0;    relay_conn far_2_2981_0_a(.in(layer_1[437]), .out(far_2_2981_0[0]));    relay_conn far_2_2981_0_b(.in(layer_1[316]), .out(far_2_2981_0[1]));
    wire [1:0] far_2_2981_1;    relay_conn far_2_2981_1_a(.in(far_2_2981_0[0]), .out(far_2_2981_1[0]));    relay_conn far_2_2981_1_b(.in(far_2_2981_0[1]), .out(far_2_2981_1[1]));
    wire [1:0] far_2_2981_2;    relay_conn far_2_2981_2_a(.in(far_2_2981_1[0]), .out(far_2_2981_2[0]));    relay_conn far_2_2981_2_b(.in(far_2_2981_1[1]), .out(far_2_2981_2[1]));
    assign layer_2[941] = far_2_2981_2[0] | far_2_2981_2[1]; 
    wire [1:0] far_2_2982_0;    relay_conn far_2_2982_0_a(.in(layer_1[167]), .out(far_2_2982_0[0]));    relay_conn far_2_2982_0_b(.in(layer_1[261]), .out(far_2_2982_0[1]));
    wire [1:0] far_2_2982_1;    relay_conn far_2_2982_1_a(.in(far_2_2982_0[0]), .out(far_2_2982_1[0]));    relay_conn far_2_2982_1_b(.in(far_2_2982_0[1]), .out(far_2_2982_1[1]));
    assign layer_2[942] = ~(far_2_2982_1[0] & far_2_2982_1[1]); 
    wire [1:0] far_2_2983_0;    relay_conn far_2_2983_0_a(.in(layer_1[663]), .out(far_2_2983_0[0]));    relay_conn far_2_2983_0_b(.in(layer_1[773]), .out(far_2_2983_0[1]));
    wire [1:0] far_2_2983_1;    relay_conn far_2_2983_1_a(.in(far_2_2983_0[0]), .out(far_2_2983_1[0]));    relay_conn far_2_2983_1_b(.in(far_2_2983_0[1]), .out(far_2_2983_1[1]));
    wire [1:0] far_2_2983_2;    relay_conn far_2_2983_2_a(.in(far_2_2983_1[0]), .out(far_2_2983_2[0]));    relay_conn far_2_2983_2_b(.in(far_2_2983_1[1]), .out(far_2_2983_2[1]));
    assign layer_2[943] = far_2_2983_2[0] ^ far_2_2983_2[1]; 
    wire [1:0] far_2_2984_0;    relay_conn far_2_2984_0_a(.in(layer_1[404]), .out(far_2_2984_0[0]));    relay_conn far_2_2984_0_b(.in(layer_1[347]), .out(far_2_2984_0[1]));
    assign layer_2[944] = ~far_2_2984_0[0]; 
    wire [1:0] far_2_2985_0;    relay_conn far_2_2985_0_a(.in(layer_1[949]), .out(far_2_2985_0[0]));    relay_conn far_2_2985_0_b(.in(layer_1[870]), .out(far_2_2985_0[1]));
    wire [1:0] far_2_2985_1;    relay_conn far_2_2985_1_a(.in(far_2_2985_0[0]), .out(far_2_2985_1[0]));    relay_conn far_2_2985_1_b(.in(far_2_2985_0[1]), .out(far_2_2985_1[1]));
    assign layer_2[945] = ~(far_2_2985_1[0] & far_2_2985_1[1]); 
    wire [1:0] far_2_2986_0;    relay_conn far_2_2986_0_a(.in(layer_1[718]), .out(far_2_2986_0[0]));    relay_conn far_2_2986_0_b(.in(layer_1[614]), .out(far_2_2986_0[1]));
    wire [1:0] far_2_2986_1;    relay_conn far_2_2986_1_a(.in(far_2_2986_0[0]), .out(far_2_2986_1[0]));    relay_conn far_2_2986_1_b(.in(far_2_2986_0[1]), .out(far_2_2986_1[1]));
    wire [1:0] far_2_2986_2;    relay_conn far_2_2986_2_a(.in(far_2_2986_1[0]), .out(far_2_2986_2[0]));    relay_conn far_2_2986_2_b(.in(far_2_2986_1[1]), .out(far_2_2986_2[1]));
    assign layer_2[946] = ~(far_2_2986_2[0] & far_2_2986_2[1]); 
    wire [1:0] far_2_2987_0;    relay_conn far_2_2987_0_a(.in(layer_1[607]), .out(far_2_2987_0[0]));    relay_conn far_2_2987_0_b(.in(layer_1[532]), .out(far_2_2987_0[1]));
    wire [1:0] far_2_2987_1;    relay_conn far_2_2987_1_a(.in(far_2_2987_0[0]), .out(far_2_2987_1[0]));    relay_conn far_2_2987_1_b(.in(far_2_2987_0[1]), .out(far_2_2987_1[1]));
    assign layer_2[947] = far_2_2987_1[0] | far_2_2987_1[1]; 
    wire [1:0] far_2_2988_0;    relay_conn far_2_2988_0_a(.in(layer_1[498]), .out(far_2_2988_0[0]));    relay_conn far_2_2988_0_b(.in(layer_1[548]), .out(far_2_2988_0[1]));
    assign layer_2[948] = ~far_2_2988_0[1]; 
    wire [1:0] far_2_2989_0;    relay_conn far_2_2989_0_a(.in(layer_1[864]), .out(far_2_2989_0[0]));    relay_conn far_2_2989_0_b(.in(layer_1[986]), .out(far_2_2989_0[1]));
    wire [1:0] far_2_2989_1;    relay_conn far_2_2989_1_a(.in(far_2_2989_0[0]), .out(far_2_2989_1[0]));    relay_conn far_2_2989_1_b(.in(far_2_2989_0[1]), .out(far_2_2989_1[1]));
    wire [1:0] far_2_2989_2;    relay_conn far_2_2989_2_a(.in(far_2_2989_1[0]), .out(far_2_2989_2[0]));    relay_conn far_2_2989_2_b(.in(far_2_2989_1[1]), .out(far_2_2989_2[1]));
    assign layer_2[949] = ~(far_2_2989_2[0] & far_2_2989_2[1]); 
    assign layer_2[950] = layer_1[527] & ~layer_1[514]; 
    wire [1:0] far_2_2991_0;    relay_conn far_2_2991_0_a(.in(layer_1[98]), .out(far_2_2991_0[0]));    relay_conn far_2_2991_0_b(.in(layer_1[25]), .out(far_2_2991_0[1]));
    wire [1:0] far_2_2991_1;    relay_conn far_2_2991_1_a(.in(far_2_2991_0[0]), .out(far_2_2991_1[0]));    relay_conn far_2_2991_1_b(.in(far_2_2991_0[1]), .out(far_2_2991_1[1]));
    assign layer_2[951] = far_2_2991_1[1]; 
    wire [1:0] far_2_2992_0;    relay_conn far_2_2992_0_a(.in(layer_1[716]), .out(far_2_2992_0[0]));    relay_conn far_2_2992_0_b(.in(layer_1[839]), .out(far_2_2992_0[1]));
    wire [1:0] far_2_2992_1;    relay_conn far_2_2992_1_a(.in(far_2_2992_0[0]), .out(far_2_2992_1[0]));    relay_conn far_2_2992_1_b(.in(far_2_2992_0[1]), .out(far_2_2992_1[1]));
    wire [1:0] far_2_2992_2;    relay_conn far_2_2992_2_a(.in(far_2_2992_1[0]), .out(far_2_2992_2[0]));    relay_conn far_2_2992_2_b(.in(far_2_2992_1[1]), .out(far_2_2992_2[1]));
    assign layer_2[952] = ~far_2_2992_2[1]; 
    wire [1:0] far_2_2993_0;    relay_conn far_2_2993_0_a(.in(layer_1[161]), .out(far_2_2993_0[0]));    relay_conn far_2_2993_0_b(.in(layer_1[221]), .out(far_2_2993_0[1]));
    assign layer_2[953] = far_2_2993_0[1]; 
    assign layer_2[954] = ~layer_1[926]; 
    wire [1:0] far_2_2995_0;    relay_conn far_2_2995_0_a(.in(layer_1[882]), .out(far_2_2995_0[0]));    relay_conn far_2_2995_0_b(.in(layer_1[797]), .out(far_2_2995_0[1]));
    wire [1:0] far_2_2995_1;    relay_conn far_2_2995_1_a(.in(far_2_2995_0[0]), .out(far_2_2995_1[0]));    relay_conn far_2_2995_1_b(.in(far_2_2995_0[1]), .out(far_2_2995_1[1]));
    assign layer_2[955] = far_2_2995_1[0]; 
    wire [1:0] far_2_2996_0;    relay_conn far_2_2996_0_a(.in(layer_1[288]), .out(far_2_2996_0[0]));    relay_conn far_2_2996_0_b(.in(layer_1[404]), .out(far_2_2996_0[1]));
    wire [1:0] far_2_2996_1;    relay_conn far_2_2996_1_a(.in(far_2_2996_0[0]), .out(far_2_2996_1[0]));    relay_conn far_2_2996_1_b(.in(far_2_2996_0[1]), .out(far_2_2996_1[1]));
    wire [1:0] far_2_2996_2;    relay_conn far_2_2996_2_a(.in(far_2_2996_1[0]), .out(far_2_2996_2[0]));    relay_conn far_2_2996_2_b(.in(far_2_2996_1[1]), .out(far_2_2996_2[1]));
    assign layer_2[956] = far_2_2996_2[1] & ~far_2_2996_2[0]; 
    assign layer_2[957] = layer_1[161] & ~layer_1[171]; 
    assign layer_2[958] = ~layer_1[776] | (layer_1[776] & layer_1[801]); 
    assign layer_2[959] = layer_1[1018] & ~layer_1[1008]; 
    assign layer_2[960] = ~layer_1[932] | (layer_1[919] & layer_1[932]); 
    assign layer_2[961] = layer_1[897]; 
    wire [1:0] far_2_3002_0;    relay_conn far_2_3002_0_a(.in(layer_1[707]), .out(far_2_3002_0[0]));    relay_conn far_2_3002_0_b(.in(layer_1[742]), .out(far_2_3002_0[1]));
    assign layer_2[962] = ~far_2_3002_0[0] | (far_2_3002_0[0] & far_2_3002_0[1]); 
    wire [1:0] far_2_3003_0;    relay_conn far_2_3003_0_a(.in(layer_1[557]), .out(far_2_3003_0[0]));    relay_conn far_2_3003_0_b(.in(layer_1[646]), .out(far_2_3003_0[1]));
    wire [1:0] far_2_3003_1;    relay_conn far_2_3003_1_a(.in(far_2_3003_0[0]), .out(far_2_3003_1[0]));    relay_conn far_2_3003_1_b(.in(far_2_3003_0[1]), .out(far_2_3003_1[1]));
    assign layer_2[963] = ~(far_2_3003_1[0] & far_2_3003_1[1]); 
    wire [1:0] far_2_3004_0;    relay_conn far_2_3004_0_a(.in(layer_1[188]), .out(far_2_3004_0[0]));    relay_conn far_2_3004_0_b(.in(layer_1[105]), .out(far_2_3004_0[1]));
    wire [1:0] far_2_3004_1;    relay_conn far_2_3004_1_a(.in(far_2_3004_0[0]), .out(far_2_3004_1[0]));    relay_conn far_2_3004_1_b(.in(far_2_3004_0[1]), .out(far_2_3004_1[1]));
    assign layer_2[964] = far_2_3004_1[0] & far_2_3004_1[1]; 
    wire [1:0] far_2_3005_0;    relay_conn far_2_3005_0_a(.in(layer_1[359]), .out(far_2_3005_0[0]));    relay_conn far_2_3005_0_b(.in(layer_1[426]), .out(far_2_3005_0[1]));
    wire [1:0] far_2_3005_1;    relay_conn far_2_3005_1_a(.in(far_2_3005_0[0]), .out(far_2_3005_1[0]));    relay_conn far_2_3005_1_b(.in(far_2_3005_0[1]), .out(far_2_3005_1[1]));
    assign layer_2[965] = ~(far_2_3005_1[0] & far_2_3005_1[1]); 
    wire [1:0] far_2_3006_0;    relay_conn far_2_3006_0_a(.in(layer_1[947]), .out(far_2_3006_0[0]));    relay_conn far_2_3006_0_b(.in(layer_1[884]), .out(far_2_3006_0[1]));
    assign layer_2[966] = ~far_2_3006_0[1] | (far_2_3006_0[0] & far_2_3006_0[1]); 
    assign layer_2[967] = layer_1[954]; 
    assign layer_2[968] = ~(layer_1[476] ^ layer_1[461]); 
    wire [1:0] far_2_3009_0;    relay_conn far_2_3009_0_a(.in(layer_1[105]), .out(far_2_3009_0[0]));    relay_conn far_2_3009_0_b(.in(layer_1[12]), .out(far_2_3009_0[1]));
    wire [1:0] far_2_3009_1;    relay_conn far_2_3009_1_a(.in(far_2_3009_0[0]), .out(far_2_3009_1[0]));    relay_conn far_2_3009_1_b(.in(far_2_3009_0[1]), .out(far_2_3009_1[1]));
    assign layer_2[969] = far_2_3009_1[0]; 
    wire [1:0] far_2_3010_0;    relay_conn far_2_3010_0_a(.in(layer_1[239]), .out(far_2_3010_0[0]));    relay_conn far_2_3010_0_b(.in(layer_1[301]), .out(far_2_3010_0[1]));
    assign layer_2[970] = ~(far_2_3010_0[0] & far_2_3010_0[1]); 
    wire [1:0] far_2_3011_0;    relay_conn far_2_3011_0_a(.in(layer_1[491]), .out(far_2_3011_0[0]));    relay_conn far_2_3011_0_b(.in(layer_1[459]), .out(far_2_3011_0[1]));
    assign layer_2[971] = ~far_2_3011_0[0]; 
    wire [1:0] far_2_3012_0;    relay_conn far_2_3012_0_a(.in(layer_1[807]), .out(far_2_3012_0[0]));    relay_conn far_2_3012_0_b(.in(layer_1[932]), .out(far_2_3012_0[1]));
    wire [1:0] far_2_3012_1;    relay_conn far_2_3012_1_a(.in(far_2_3012_0[0]), .out(far_2_3012_1[0]));    relay_conn far_2_3012_1_b(.in(far_2_3012_0[1]), .out(far_2_3012_1[1]));
    wire [1:0] far_2_3012_2;    relay_conn far_2_3012_2_a(.in(far_2_3012_1[0]), .out(far_2_3012_2[0]));    relay_conn far_2_3012_2_b(.in(far_2_3012_1[1]), .out(far_2_3012_2[1]));
    assign layer_2[972] = far_2_3012_2[1] & ~far_2_3012_2[0]; 
    wire [1:0] far_2_3013_0;    relay_conn far_2_3013_0_a(.in(layer_1[701]), .out(far_2_3013_0[0]));    relay_conn far_2_3013_0_b(.in(layer_1[820]), .out(far_2_3013_0[1]));
    wire [1:0] far_2_3013_1;    relay_conn far_2_3013_1_a(.in(far_2_3013_0[0]), .out(far_2_3013_1[0]));    relay_conn far_2_3013_1_b(.in(far_2_3013_0[1]), .out(far_2_3013_1[1]));
    wire [1:0] far_2_3013_2;    relay_conn far_2_3013_2_a(.in(far_2_3013_1[0]), .out(far_2_3013_2[0]));    relay_conn far_2_3013_2_b(.in(far_2_3013_1[1]), .out(far_2_3013_2[1]));
    assign layer_2[973] = far_2_3013_2[0] & ~far_2_3013_2[1]; 
    assign layer_2[974] = layer_1[707] & ~layer_1[703]; 
    wire [1:0] far_2_3015_0;    relay_conn far_2_3015_0_a(.in(layer_1[145]), .out(far_2_3015_0[0]));    relay_conn far_2_3015_0_b(.in(layer_1[40]), .out(far_2_3015_0[1]));
    wire [1:0] far_2_3015_1;    relay_conn far_2_3015_1_a(.in(far_2_3015_0[0]), .out(far_2_3015_1[0]));    relay_conn far_2_3015_1_b(.in(far_2_3015_0[1]), .out(far_2_3015_1[1]));
    wire [1:0] far_2_3015_2;    relay_conn far_2_3015_2_a(.in(far_2_3015_1[0]), .out(far_2_3015_2[0]));    relay_conn far_2_3015_2_b(.in(far_2_3015_1[1]), .out(far_2_3015_2[1]));
    assign layer_2[975] = far_2_3015_2[0] | far_2_3015_2[1]; 
    wire [1:0] far_2_3016_0;    relay_conn far_2_3016_0_a(.in(layer_1[891]), .out(far_2_3016_0[0]));    relay_conn far_2_3016_0_b(.in(layer_1[930]), .out(far_2_3016_0[1]));
    assign layer_2[976] = far_2_3016_0[0] & far_2_3016_0[1]; 
    wire [1:0] far_2_3017_0;    relay_conn far_2_3017_0_a(.in(layer_1[793]), .out(far_2_3017_0[0]));    relay_conn far_2_3017_0_b(.in(layer_1[743]), .out(far_2_3017_0[1]));
    assign layer_2[977] = far_2_3017_0[0] | far_2_3017_0[1]; 
    wire [1:0] far_2_3018_0;    relay_conn far_2_3018_0_a(.in(layer_1[383]), .out(far_2_3018_0[0]));    relay_conn far_2_3018_0_b(.in(layer_1[492]), .out(far_2_3018_0[1]));
    wire [1:0] far_2_3018_1;    relay_conn far_2_3018_1_a(.in(far_2_3018_0[0]), .out(far_2_3018_1[0]));    relay_conn far_2_3018_1_b(.in(far_2_3018_0[1]), .out(far_2_3018_1[1]));
    wire [1:0] far_2_3018_2;    relay_conn far_2_3018_2_a(.in(far_2_3018_1[0]), .out(far_2_3018_2[0]));    relay_conn far_2_3018_2_b(.in(far_2_3018_1[1]), .out(far_2_3018_2[1]));
    assign layer_2[978] = ~(far_2_3018_2[0] & far_2_3018_2[1]); 
    wire [1:0] far_2_3019_0;    relay_conn far_2_3019_0_a(.in(layer_1[432]), .out(far_2_3019_0[0]));    relay_conn far_2_3019_0_b(.in(layer_1[315]), .out(far_2_3019_0[1]));
    wire [1:0] far_2_3019_1;    relay_conn far_2_3019_1_a(.in(far_2_3019_0[0]), .out(far_2_3019_1[0]));    relay_conn far_2_3019_1_b(.in(far_2_3019_0[1]), .out(far_2_3019_1[1]));
    wire [1:0] far_2_3019_2;    relay_conn far_2_3019_2_a(.in(far_2_3019_1[0]), .out(far_2_3019_2[0]));    relay_conn far_2_3019_2_b(.in(far_2_3019_1[1]), .out(far_2_3019_2[1]));
    assign layer_2[979] = ~(far_2_3019_2[0] & far_2_3019_2[1]); 
    assign layer_2[980] = ~(layer_1[924] ^ layer_1[950]); 
    wire [1:0] far_2_3021_0;    relay_conn far_2_3021_0_a(.in(layer_1[928]), .out(far_2_3021_0[0]));    relay_conn far_2_3021_0_b(.in(layer_1[856]), .out(far_2_3021_0[1]));
    wire [1:0] far_2_3021_1;    relay_conn far_2_3021_1_a(.in(far_2_3021_0[0]), .out(far_2_3021_1[0]));    relay_conn far_2_3021_1_b(.in(far_2_3021_0[1]), .out(far_2_3021_1[1]));
    assign layer_2[981] = far_2_3021_1[1] & ~far_2_3021_1[0]; 
    assign layer_2[982] = layer_1[464]; 
    wire [1:0] far_2_3023_0;    relay_conn far_2_3023_0_a(.in(layer_1[878]), .out(far_2_3023_0[0]));    relay_conn far_2_3023_0_b(.in(layer_1[795]), .out(far_2_3023_0[1]));
    wire [1:0] far_2_3023_1;    relay_conn far_2_3023_1_a(.in(far_2_3023_0[0]), .out(far_2_3023_1[0]));    relay_conn far_2_3023_1_b(.in(far_2_3023_0[1]), .out(far_2_3023_1[1]));
    assign layer_2[983] = ~(far_2_3023_1[0] ^ far_2_3023_1[1]); 
    wire [1:0] far_2_3024_0;    relay_conn far_2_3024_0_a(.in(layer_1[619]), .out(far_2_3024_0[0]));    relay_conn far_2_3024_0_b(.in(layer_1[502]), .out(far_2_3024_0[1]));
    wire [1:0] far_2_3024_1;    relay_conn far_2_3024_1_a(.in(far_2_3024_0[0]), .out(far_2_3024_1[0]));    relay_conn far_2_3024_1_b(.in(far_2_3024_0[1]), .out(far_2_3024_1[1]));
    wire [1:0] far_2_3024_2;    relay_conn far_2_3024_2_a(.in(far_2_3024_1[0]), .out(far_2_3024_2[0]));    relay_conn far_2_3024_2_b(.in(far_2_3024_1[1]), .out(far_2_3024_2[1]));
    assign layer_2[984] = far_2_3024_2[0] | far_2_3024_2[1]; 
    assign layer_2[985] = layer_1[9] | layer_1[40]; 
    assign layer_2[986] = layer_1[44] | layer_1[57]; 
    wire [1:0] far_2_3027_0;    relay_conn far_2_3027_0_a(.in(layer_1[346]), .out(far_2_3027_0[0]));    relay_conn far_2_3027_0_b(.in(layer_1[458]), .out(far_2_3027_0[1]));
    wire [1:0] far_2_3027_1;    relay_conn far_2_3027_1_a(.in(far_2_3027_0[0]), .out(far_2_3027_1[0]));    relay_conn far_2_3027_1_b(.in(far_2_3027_0[1]), .out(far_2_3027_1[1]));
    wire [1:0] far_2_3027_2;    relay_conn far_2_3027_2_a(.in(far_2_3027_1[0]), .out(far_2_3027_2[0]));    relay_conn far_2_3027_2_b(.in(far_2_3027_1[1]), .out(far_2_3027_2[1]));
    assign layer_2[987] = far_2_3027_2[0] & far_2_3027_2[1]; 
    wire [1:0] far_2_3028_0;    relay_conn far_2_3028_0_a(.in(layer_1[656]), .out(far_2_3028_0[0]));    relay_conn far_2_3028_0_b(.in(layer_1[742]), .out(far_2_3028_0[1]));
    wire [1:0] far_2_3028_1;    relay_conn far_2_3028_1_a(.in(far_2_3028_0[0]), .out(far_2_3028_1[0]));    relay_conn far_2_3028_1_b(.in(far_2_3028_0[1]), .out(far_2_3028_1[1]));
    assign layer_2[988] = far_2_3028_1[1]; 
    wire [1:0] far_2_3029_0;    relay_conn far_2_3029_0_a(.in(layer_1[67]), .out(far_2_3029_0[0]));    relay_conn far_2_3029_0_b(.in(layer_1[102]), .out(far_2_3029_0[1]));
    assign layer_2[989] = ~far_2_3029_0[0]; 
    wire [1:0] far_2_3030_0;    relay_conn far_2_3030_0_a(.in(layer_1[127]), .out(far_2_3030_0[0]));    relay_conn far_2_3030_0_b(.in(layer_1[236]), .out(far_2_3030_0[1]));
    wire [1:0] far_2_3030_1;    relay_conn far_2_3030_1_a(.in(far_2_3030_0[0]), .out(far_2_3030_1[0]));    relay_conn far_2_3030_1_b(.in(far_2_3030_0[1]), .out(far_2_3030_1[1]));
    wire [1:0] far_2_3030_2;    relay_conn far_2_3030_2_a(.in(far_2_3030_1[0]), .out(far_2_3030_2[0]));    relay_conn far_2_3030_2_b(.in(far_2_3030_1[1]), .out(far_2_3030_2[1]));
    assign layer_2[990] = far_2_3030_2[0] | far_2_3030_2[1]; 
    wire [1:0] far_2_3031_0;    relay_conn far_2_3031_0_a(.in(layer_1[983]), .out(far_2_3031_0[0]));    relay_conn far_2_3031_0_b(.in(layer_1[1019]), .out(far_2_3031_0[1]));
    assign layer_2[991] = far_2_3031_0[0] & far_2_3031_0[1]; 
    wire [1:0] far_2_3032_0;    relay_conn far_2_3032_0_a(.in(layer_1[723]), .out(far_2_3032_0[0]));    relay_conn far_2_3032_0_b(.in(layer_1[798]), .out(far_2_3032_0[1]));
    wire [1:0] far_2_3032_1;    relay_conn far_2_3032_1_a(.in(far_2_3032_0[0]), .out(far_2_3032_1[0]));    relay_conn far_2_3032_1_b(.in(far_2_3032_0[1]), .out(far_2_3032_1[1]));
    assign layer_2[992] = far_2_3032_1[0] | far_2_3032_1[1]; 
    wire [1:0] far_2_3033_0;    relay_conn far_2_3033_0_a(.in(layer_1[338]), .out(far_2_3033_0[0]));    relay_conn far_2_3033_0_b(.in(layer_1[439]), .out(far_2_3033_0[1]));
    wire [1:0] far_2_3033_1;    relay_conn far_2_3033_1_a(.in(far_2_3033_0[0]), .out(far_2_3033_1[0]));    relay_conn far_2_3033_1_b(.in(far_2_3033_0[1]), .out(far_2_3033_1[1]));
    wire [1:0] far_2_3033_2;    relay_conn far_2_3033_2_a(.in(far_2_3033_1[0]), .out(far_2_3033_2[0]));    relay_conn far_2_3033_2_b(.in(far_2_3033_1[1]), .out(far_2_3033_2[1]));
    assign layer_2[993] = far_2_3033_2[1] & ~far_2_3033_2[0]; 
    wire [1:0] far_2_3034_0;    relay_conn far_2_3034_0_a(.in(layer_1[516]), .out(far_2_3034_0[0]));    relay_conn far_2_3034_0_b(.in(layer_1[446]), .out(far_2_3034_0[1]));
    wire [1:0] far_2_3034_1;    relay_conn far_2_3034_1_a(.in(far_2_3034_0[0]), .out(far_2_3034_1[0]));    relay_conn far_2_3034_1_b(.in(far_2_3034_0[1]), .out(far_2_3034_1[1]));
    assign layer_2[994] = far_2_3034_1[0]; 
    wire [1:0] far_2_3035_0;    relay_conn far_2_3035_0_a(.in(layer_1[777]), .out(far_2_3035_0[0]));    relay_conn far_2_3035_0_b(.in(layer_1[690]), .out(far_2_3035_0[1]));
    wire [1:0] far_2_3035_1;    relay_conn far_2_3035_1_a(.in(far_2_3035_0[0]), .out(far_2_3035_1[0]));    relay_conn far_2_3035_1_b(.in(far_2_3035_0[1]), .out(far_2_3035_1[1]));
    assign layer_2[995] = ~(far_2_3035_1[0] | far_2_3035_1[1]); 
    wire [1:0] far_2_3036_0;    relay_conn far_2_3036_0_a(.in(layer_1[32]), .out(far_2_3036_0[0]));    relay_conn far_2_3036_0_b(.in(layer_1[110]), .out(far_2_3036_0[1]));
    wire [1:0] far_2_3036_1;    relay_conn far_2_3036_1_a(.in(far_2_3036_0[0]), .out(far_2_3036_1[0]));    relay_conn far_2_3036_1_b(.in(far_2_3036_0[1]), .out(far_2_3036_1[1]));
    assign layer_2[996] = ~far_2_3036_1[1]; 
    wire [1:0] far_2_3037_0;    relay_conn far_2_3037_0_a(.in(layer_1[740]), .out(far_2_3037_0[0]));    relay_conn far_2_3037_0_b(.in(layer_1[866]), .out(far_2_3037_0[1]));
    wire [1:0] far_2_3037_1;    relay_conn far_2_3037_1_a(.in(far_2_3037_0[0]), .out(far_2_3037_1[0]));    relay_conn far_2_3037_1_b(.in(far_2_3037_0[1]), .out(far_2_3037_1[1]));
    wire [1:0] far_2_3037_2;    relay_conn far_2_3037_2_a(.in(far_2_3037_1[0]), .out(far_2_3037_2[0]));    relay_conn far_2_3037_2_b(.in(far_2_3037_1[1]), .out(far_2_3037_2[1]));
    assign layer_2[997] = far_2_3037_2[0] & ~far_2_3037_2[1]; 
    wire [1:0] far_2_3038_0;    relay_conn far_2_3038_0_a(.in(layer_1[669]), .out(far_2_3038_0[0]));    relay_conn far_2_3038_0_b(.in(layer_1[557]), .out(far_2_3038_0[1]));
    wire [1:0] far_2_3038_1;    relay_conn far_2_3038_1_a(.in(far_2_3038_0[0]), .out(far_2_3038_1[0]));    relay_conn far_2_3038_1_b(.in(far_2_3038_0[1]), .out(far_2_3038_1[1]));
    wire [1:0] far_2_3038_2;    relay_conn far_2_3038_2_a(.in(far_2_3038_1[0]), .out(far_2_3038_2[0]));    relay_conn far_2_3038_2_b(.in(far_2_3038_1[1]), .out(far_2_3038_2[1]));
    assign layer_2[998] = ~far_2_3038_2[0] | (far_2_3038_2[0] & far_2_3038_2[1]); 
    wire [1:0] far_2_3039_0;    relay_conn far_2_3039_0_a(.in(layer_1[930]), .out(far_2_3039_0[0]));    relay_conn far_2_3039_0_b(.in(layer_1[966]), .out(far_2_3039_0[1]));
    assign layer_2[999] = ~(far_2_3039_0[0] ^ far_2_3039_0[1]); 
    wire [1:0] far_2_3040_0;    relay_conn far_2_3040_0_a(.in(layer_1[661]), .out(far_2_3040_0[0]));    relay_conn far_2_3040_0_b(.in(layer_1[581]), .out(far_2_3040_0[1]));
    wire [1:0] far_2_3040_1;    relay_conn far_2_3040_1_a(.in(far_2_3040_0[0]), .out(far_2_3040_1[0]));    relay_conn far_2_3040_1_b(.in(far_2_3040_0[1]), .out(far_2_3040_1[1]));
    assign layer_2[1000] = ~far_2_3040_1[0] | (far_2_3040_1[0] & far_2_3040_1[1]); 
    wire [1:0] far_2_3041_0;    relay_conn far_2_3041_0_a(.in(layer_1[607]), .out(far_2_3041_0[0]));    relay_conn far_2_3041_0_b(.in(layer_1[643]), .out(far_2_3041_0[1]));
    assign layer_2[1001] = ~far_2_3041_0[1] | (far_2_3041_0[0] & far_2_3041_0[1]); 
    wire [1:0] far_2_3042_0;    relay_conn far_2_3042_0_a(.in(layer_1[251]), .out(far_2_3042_0[0]));    relay_conn far_2_3042_0_b(.in(layer_1[153]), .out(far_2_3042_0[1]));
    wire [1:0] far_2_3042_1;    relay_conn far_2_3042_1_a(.in(far_2_3042_0[0]), .out(far_2_3042_1[0]));    relay_conn far_2_3042_1_b(.in(far_2_3042_0[1]), .out(far_2_3042_1[1]));
    wire [1:0] far_2_3042_2;    relay_conn far_2_3042_2_a(.in(far_2_3042_1[0]), .out(far_2_3042_2[0]));    relay_conn far_2_3042_2_b(.in(far_2_3042_1[1]), .out(far_2_3042_2[1]));
    assign layer_2[1002] = ~(far_2_3042_2[0] | far_2_3042_2[1]); 
    wire [1:0] far_2_3043_0;    relay_conn far_2_3043_0_a(.in(layer_1[620]), .out(far_2_3043_0[0]));    relay_conn far_2_3043_0_b(.in(layer_1[695]), .out(far_2_3043_0[1]));
    wire [1:0] far_2_3043_1;    relay_conn far_2_3043_1_a(.in(far_2_3043_0[0]), .out(far_2_3043_1[0]));    relay_conn far_2_3043_1_b(.in(far_2_3043_0[1]), .out(far_2_3043_1[1]));
    assign layer_2[1003] = far_2_3043_1[0] & ~far_2_3043_1[1]; 
    assign layer_2[1004] = ~layer_1[303] | (layer_1[303] & layer_1[278]); 
    wire [1:0] far_2_3045_0;    relay_conn far_2_3045_0_a(.in(layer_1[184]), .out(far_2_3045_0[0]));    relay_conn far_2_3045_0_b(.in(layer_1[127]), .out(far_2_3045_0[1]));
    assign layer_2[1005] = far_2_3045_0[1]; 
    assign layer_2[1006] = layer_1[987]; 
    wire [1:0] far_2_3047_0;    relay_conn far_2_3047_0_a(.in(layer_1[864]), .out(far_2_3047_0[0]));    relay_conn far_2_3047_0_b(.in(layer_1[768]), .out(far_2_3047_0[1]));
    wire [1:0] far_2_3047_1;    relay_conn far_2_3047_1_a(.in(far_2_3047_0[0]), .out(far_2_3047_1[0]));    relay_conn far_2_3047_1_b(.in(far_2_3047_0[1]), .out(far_2_3047_1[1]));
    wire [1:0] far_2_3047_2;    relay_conn far_2_3047_2_a(.in(far_2_3047_1[0]), .out(far_2_3047_2[0]));    relay_conn far_2_3047_2_b(.in(far_2_3047_1[1]), .out(far_2_3047_2[1]));
    assign layer_2[1007] = far_2_3047_2[1]; 
    wire [1:0] far_2_3048_0;    relay_conn far_2_3048_0_a(.in(layer_1[87]), .out(far_2_3048_0[0]));    relay_conn far_2_3048_0_b(.in(layer_1[208]), .out(far_2_3048_0[1]));
    wire [1:0] far_2_3048_1;    relay_conn far_2_3048_1_a(.in(far_2_3048_0[0]), .out(far_2_3048_1[0]));    relay_conn far_2_3048_1_b(.in(far_2_3048_0[1]), .out(far_2_3048_1[1]));
    wire [1:0] far_2_3048_2;    relay_conn far_2_3048_2_a(.in(far_2_3048_1[0]), .out(far_2_3048_2[0]));    relay_conn far_2_3048_2_b(.in(far_2_3048_1[1]), .out(far_2_3048_2[1]));
    assign layer_2[1008] = ~(far_2_3048_2[0] & far_2_3048_2[1]); 
    assign layer_2[1009] = layer_1[926] & ~layer_1[910]; 
    wire [1:0] far_2_3050_0;    relay_conn far_2_3050_0_a(.in(layer_1[555]), .out(far_2_3050_0[0]));    relay_conn far_2_3050_0_b(.in(layer_1[455]), .out(far_2_3050_0[1]));
    wire [1:0] far_2_3050_1;    relay_conn far_2_3050_1_a(.in(far_2_3050_0[0]), .out(far_2_3050_1[0]));    relay_conn far_2_3050_1_b(.in(far_2_3050_0[1]), .out(far_2_3050_1[1]));
    wire [1:0] far_2_3050_2;    relay_conn far_2_3050_2_a(.in(far_2_3050_1[0]), .out(far_2_3050_2[0]));    relay_conn far_2_3050_2_b(.in(far_2_3050_1[1]), .out(far_2_3050_2[1]));
    assign layer_2[1010] = ~far_2_3050_2[1]; 
    wire [1:0] far_2_3051_0;    relay_conn far_2_3051_0_a(.in(layer_1[812]), .out(far_2_3051_0[0]));    relay_conn far_2_3051_0_b(.in(layer_1[737]), .out(far_2_3051_0[1]));
    wire [1:0] far_2_3051_1;    relay_conn far_2_3051_1_a(.in(far_2_3051_0[0]), .out(far_2_3051_1[0]));    relay_conn far_2_3051_1_b(.in(far_2_3051_0[1]), .out(far_2_3051_1[1]));
    assign layer_2[1011] = ~(far_2_3051_1[0] ^ far_2_3051_1[1]); 
    assign layer_2[1012] = layer_1[228] & layer_1[259]; 
    assign layer_2[1013] = ~layer_1[367]; 
    assign layer_2[1014] = ~(layer_1[104] ^ layer_1[130]); 
    assign layer_2[1015] = layer_1[616] & ~layer_1[628]; 
    wire [1:0] far_2_3056_0;    relay_conn far_2_3056_0_a(.in(layer_1[419]), .out(far_2_3056_0[0]));    relay_conn far_2_3056_0_b(.in(layer_1[293]), .out(far_2_3056_0[1]));
    wire [1:0] far_2_3056_1;    relay_conn far_2_3056_1_a(.in(far_2_3056_0[0]), .out(far_2_3056_1[0]));    relay_conn far_2_3056_1_b(.in(far_2_3056_0[1]), .out(far_2_3056_1[1]));
    wire [1:0] far_2_3056_2;    relay_conn far_2_3056_2_a(.in(far_2_3056_1[0]), .out(far_2_3056_2[0]));    relay_conn far_2_3056_2_b(.in(far_2_3056_1[1]), .out(far_2_3056_2[1]));
    assign layer_2[1016] = ~far_2_3056_2[0]; 
    wire [1:0] far_2_3057_0;    relay_conn far_2_3057_0_a(.in(layer_1[443]), .out(far_2_3057_0[0]));    relay_conn far_2_3057_0_b(.in(layer_1[323]), .out(far_2_3057_0[1]));
    wire [1:0] far_2_3057_1;    relay_conn far_2_3057_1_a(.in(far_2_3057_0[0]), .out(far_2_3057_1[0]));    relay_conn far_2_3057_1_b(.in(far_2_3057_0[1]), .out(far_2_3057_1[1]));
    wire [1:0] far_2_3057_2;    relay_conn far_2_3057_2_a(.in(far_2_3057_1[0]), .out(far_2_3057_2[0]));    relay_conn far_2_3057_2_b(.in(far_2_3057_1[1]), .out(far_2_3057_2[1]));
    assign layer_2[1017] = ~(far_2_3057_2[0] | far_2_3057_2[1]); 
    assign layer_2[1018] = layer_1[353]; 
    wire [1:0] far_2_3059_0;    relay_conn far_2_3059_0_a(.in(layer_1[12]), .out(far_2_3059_0[0]));    relay_conn far_2_3059_0_b(.in(layer_1[52]), .out(far_2_3059_0[1]));
    assign layer_2[1019] = ~far_2_3059_0[1] | (far_2_3059_0[0] & far_2_3059_0[1]); 
    // Layer 3 ============================================================
    wire [1:0] far_3_3060_0;    relay_conn far_3_3060_0_a(.in(layer_2[978]), .out(far_3_3060_0[0]));    relay_conn far_3_3060_0_b(.in(layer_2[946]), .out(far_3_3060_0[1]));
    assign layer_3[0] = far_3_3060_0[1]; 
    wire [1:0] far_3_3061_0;    relay_conn far_3_3061_0_a(.in(layer_2[580]), .out(far_3_3061_0[0]));    relay_conn far_3_3061_0_b(.in(layer_2[519]), .out(far_3_3061_0[1]));
    assign layer_3[1] = far_3_3061_0[1]; 
    wire [1:0] far_3_3062_0;    relay_conn far_3_3062_0_a(.in(layer_2[534]), .out(far_3_3062_0[0]));    relay_conn far_3_3062_0_b(.in(layer_2[482]), .out(far_3_3062_0[1]));
    assign layer_3[2] = ~far_3_3062_0[0] | (far_3_3062_0[0] & far_3_3062_0[1]); 
    wire [1:0] far_3_3063_0;    relay_conn far_3_3063_0_a(.in(layer_2[588]), .out(far_3_3063_0[0]));    relay_conn far_3_3063_0_b(.in(layer_2[468]), .out(far_3_3063_0[1]));
    wire [1:0] far_3_3063_1;    relay_conn far_3_3063_1_a(.in(far_3_3063_0[0]), .out(far_3_3063_1[0]));    relay_conn far_3_3063_1_b(.in(far_3_3063_0[1]), .out(far_3_3063_1[1]));
    wire [1:0] far_3_3063_2;    relay_conn far_3_3063_2_a(.in(far_3_3063_1[0]), .out(far_3_3063_2[0]));    relay_conn far_3_3063_2_b(.in(far_3_3063_1[1]), .out(far_3_3063_2[1]));
    assign layer_3[3] = ~(far_3_3063_2[0] | far_3_3063_2[1]); 
    wire [1:0] far_3_3064_0;    relay_conn far_3_3064_0_a(.in(layer_2[365]), .out(far_3_3064_0[0]));    relay_conn far_3_3064_0_b(.in(layer_2[247]), .out(far_3_3064_0[1]));
    wire [1:0] far_3_3064_1;    relay_conn far_3_3064_1_a(.in(far_3_3064_0[0]), .out(far_3_3064_1[0]));    relay_conn far_3_3064_1_b(.in(far_3_3064_0[1]), .out(far_3_3064_1[1]));
    wire [1:0] far_3_3064_2;    relay_conn far_3_3064_2_a(.in(far_3_3064_1[0]), .out(far_3_3064_2[0]));    relay_conn far_3_3064_2_b(.in(far_3_3064_1[1]), .out(far_3_3064_2[1]));
    assign layer_3[4] = far_3_3064_2[0] | far_3_3064_2[1]; 
    wire [1:0] far_3_3065_0;    relay_conn far_3_3065_0_a(.in(layer_2[819]), .out(far_3_3065_0[0]));    relay_conn far_3_3065_0_b(.in(layer_2[728]), .out(far_3_3065_0[1]));
    wire [1:0] far_3_3065_1;    relay_conn far_3_3065_1_a(.in(far_3_3065_0[0]), .out(far_3_3065_1[0]));    relay_conn far_3_3065_1_b(.in(far_3_3065_0[1]), .out(far_3_3065_1[1]));
    assign layer_3[5] = far_3_3065_1[1] & ~far_3_3065_1[0]; 
    wire [1:0] far_3_3066_0;    relay_conn far_3_3066_0_a(.in(layer_2[765]), .out(far_3_3066_0[0]));    relay_conn far_3_3066_0_b(.in(layer_2[664]), .out(far_3_3066_0[1]));
    wire [1:0] far_3_3066_1;    relay_conn far_3_3066_1_a(.in(far_3_3066_0[0]), .out(far_3_3066_1[0]));    relay_conn far_3_3066_1_b(.in(far_3_3066_0[1]), .out(far_3_3066_1[1]));
    wire [1:0] far_3_3066_2;    relay_conn far_3_3066_2_a(.in(far_3_3066_1[0]), .out(far_3_3066_2[0]));    relay_conn far_3_3066_2_b(.in(far_3_3066_1[1]), .out(far_3_3066_2[1]));
    assign layer_3[6] = ~far_3_3066_2[0]; 
    wire [1:0] far_3_3067_0;    relay_conn far_3_3067_0_a(.in(layer_2[33]), .out(far_3_3067_0[0]));    relay_conn far_3_3067_0_b(.in(layer_2[144]), .out(far_3_3067_0[1]));
    wire [1:0] far_3_3067_1;    relay_conn far_3_3067_1_a(.in(far_3_3067_0[0]), .out(far_3_3067_1[0]));    relay_conn far_3_3067_1_b(.in(far_3_3067_0[1]), .out(far_3_3067_1[1]));
    wire [1:0] far_3_3067_2;    relay_conn far_3_3067_2_a(.in(far_3_3067_1[0]), .out(far_3_3067_2[0]));    relay_conn far_3_3067_2_b(.in(far_3_3067_1[1]), .out(far_3_3067_2[1]));
    assign layer_3[7] = far_3_3067_2[0] & ~far_3_3067_2[1]; 
    wire [1:0] far_3_3068_0;    relay_conn far_3_3068_0_a(.in(layer_2[433]), .out(far_3_3068_0[0]));    relay_conn far_3_3068_0_b(.in(layer_2[500]), .out(far_3_3068_0[1]));
    wire [1:0] far_3_3068_1;    relay_conn far_3_3068_1_a(.in(far_3_3068_0[0]), .out(far_3_3068_1[0]));    relay_conn far_3_3068_1_b(.in(far_3_3068_0[1]), .out(far_3_3068_1[1]));
    assign layer_3[8] = far_3_3068_1[0] & far_3_3068_1[1]; 
    wire [1:0] far_3_3069_0;    relay_conn far_3_3069_0_a(.in(layer_2[303]), .out(far_3_3069_0[0]));    relay_conn far_3_3069_0_b(.in(layer_2[205]), .out(far_3_3069_0[1]));
    wire [1:0] far_3_3069_1;    relay_conn far_3_3069_1_a(.in(far_3_3069_0[0]), .out(far_3_3069_1[0]));    relay_conn far_3_3069_1_b(.in(far_3_3069_0[1]), .out(far_3_3069_1[1]));
    wire [1:0] far_3_3069_2;    relay_conn far_3_3069_2_a(.in(far_3_3069_1[0]), .out(far_3_3069_2[0]));    relay_conn far_3_3069_2_b(.in(far_3_3069_1[1]), .out(far_3_3069_2[1]));
    assign layer_3[9] = ~far_3_3069_2[0]; 
    wire [1:0] far_3_3070_0;    relay_conn far_3_3070_0_a(.in(layer_2[424]), .out(far_3_3070_0[0]));    relay_conn far_3_3070_0_b(.in(layer_2[466]), .out(far_3_3070_0[1]));
    assign layer_3[10] = far_3_3070_0[0]; 
    wire [1:0] far_3_3071_0;    relay_conn far_3_3071_0_a(.in(layer_2[462]), .out(far_3_3071_0[0]));    relay_conn far_3_3071_0_b(.in(layer_2[573]), .out(far_3_3071_0[1]));
    wire [1:0] far_3_3071_1;    relay_conn far_3_3071_1_a(.in(far_3_3071_0[0]), .out(far_3_3071_1[0]));    relay_conn far_3_3071_1_b(.in(far_3_3071_0[1]), .out(far_3_3071_1[1]));
    wire [1:0] far_3_3071_2;    relay_conn far_3_3071_2_a(.in(far_3_3071_1[0]), .out(far_3_3071_2[0]));    relay_conn far_3_3071_2_b(.in(far_3_3071_1[1]), .out(far_3_3071_2[1]));
    assign layer_3[11] = ~far_3_3071_2[1]; 
    wire [1:0] far_3_3072_0;    relay_conn far_3_3072_0_a(.in(layer_2[970]), .out(far_3_3072_0[0]));    relay_conn far_3_3072_0_b(.in(layer_2[872]), .out(far_3_3072_0[1]));
    wire [1:0] far_3_3072_1;    relay_conn far_3_3072_1_a(.in(far_3_3072_0[0]), .out(far_3_3072_1[0]));    relay_conn far_3_3072_1_b(.in(far_3_3072_0[1]), .out(far_3_3072_1[1]));
    wire [1:0] far_3_3072_2;    relay_conn far_3_3072_2_a(.in(far_3_3072_1[0]), .out(far_3_3072_2[0]));    relay_conn far_3_3072_2_b(.in(far_3_3072_1[1]), .out(far_3_3072_2[1]));
    assign layer_3[12] = far_3_3072_2[0] | far_3_3072_2[1]; 
    wire [1:0] far_3_3073_0;    relay_conn far_3_3073_0_a(.in(layer_2[352]), .out(far_3_3073_0[0]));    relay_conn far_3_3073_0_b(.in(layer_2[237]), .out(far_3_3073_0[1]));
    wire [1:0] far_3_3073_1;    relay_conn far_3_3073_1_a(.in(far_3_3073_0[0]), .out(far_3_3073_1[0]));    relay_conn far_3_3073_1_b(.in(far_3_3073_0[1]), .out(far_3_3073_1[1]));
    wire [1:0] far_3_3073_2;    relay_conn far_3_3073_2_a(.in(far_3_3073_1[0]), .out(far_3_3073_2[0]));    relay_conn far_3_3073_2_b(.in(far_3_3073_1[1]), .out(far_3_3073_2[1]));
    assign layer_3[13] = ~(far_3_3073_2[0] ^ far_3_3073_2[1]); 
    wire [1:0] far_3_3074_0;    relay_conn far_3_3074_0_a(.in(layer_2[94]), .out(far_3_3074_0[0]));    relay_conn far_3_3074_0_b(.in(layer_2[130]), .out(far_3_3074_0[1]));
    assign layer_3[14] = far_3_3074_0[1] & ~far_3_3074_0[0]; 
    wire [1:0] far_3_3075_0;    relay_conn far_3_3075_0_a(.in(layer_2[730]), .out(far_3_3075_0[0]));    relay_conn far_3_3075_0_b(.in(layer_2[821]), .out(far_3_3075_0[1]));
    wire [1:0] far_3_3075_1;    relay_conn far_3_3075_1_a(.in(far_3_3075_0[0]), .out(far_3_3075_1[0]));    relay_conn far_3_3075_1_b(.in(far_3_3075_0[1]), .out(far_3_3075_1[1]));
    assign layer_3[15] = ~far_3_3075_1[1] | (far_3_3075_1[0] & far_3_3075_1[1]); 
    wire [1:0] far_3_3076_0;    relay_conn far_3_3076_0_a(.in(layer_2[39]), .out(far_3_3076_0[0]));    relay_conn far_3_3076_0_b(.in(layer_2[3]), .out(far_3_3076_0[1]));
    assign layer_3[16] = far_3_3076_0[0] & far_3_3076_0[1]; 
    wire [1:0] far_3_3077_0;    relay_conn far_3_3077_0_a(.in(layer_2[354]), .out(far_3_3077_0[0]));    relay_conn far_3_3077_0_b(.in(layer_2[414]), .out(far_3_3077_0[1]));
    assign layer_3[17] = ~far_3_3077_0[1]; 
    wire [1:0] far_3_3078_0;    relay_conn far_3_3078_0_a(.in(layer_2[57]), .out(far_3_3078_0[0]));    relay_conn far_3_3078_0_b(.in(layer_2[4]), .out(far_3_3078_0[1]));
    assign layer_3[18] = far_3_3078_0[0] & ~far_3_3078_0[1]; 
    wire [1:0] far_3_3079_0;    relay_conn far_3_3079_0_a(.in(layer_2[307]), .out(far_3_3079_0[0]));    relay_conn far_3_3079_0_b(.in(layer_2[346]), .out(far_3_3079_0[1]));
    assign layer_3[19] = ~far_3_3079_0[1]; 
    wire [1:0] far_3_3080_0;    relay_conn far_3_3080_0_a(.in(layer_2[336]), .out(far_3_3080_0[0]));    relay_conn far_3_3080_0_b(.in(layer_2[460]), .out(far_3_3080_0[1]));
    wire [1:0] far_3_3080_1;    relay_conn far_3_3080_1_a(.in(far_3_3080_0[0]), .out(far_3_3080_1[0]));    relay_conn far_3_3080_1_b(.in(far_3_3080_0[1]), .out(far_3_3080_1[1]));
    wire [1:0] far_3_3080_2;    relay_conn far_3_3080_2_a(.in(far_3_3080_1[0]), .out(far_3_3080_2[0]));    relay_conn far_3_3080_2_b(.in(far_3_3080_1[1]), .out(far_3_3080_2[1]));
    assign layer_3[20] = far_3_3080_2[1]; 
    wire [1:0] far_3_3081_0;    relay_conn far_3_3081_0_a(.in(layer_2[708]), .out(far_3_3081_0[0]));    relay_conn far_3_3081_0_b(.in(layer_2[809]), .out(far_3_3081_0[1]));
    wire [1:0] far_3_3081_1;    relay_conn far_3_3081_1_a(.in(far_3_3081_0[0]), .out(far_3_3081_1[0]));    relay_conn far_3_3081_1_b(.in(far_3_3081_0[1]), .out(far_3_3081_1[1]));
    wire [1:0] far_3_3081_2;    relay_conn far_3_3081_2_a(.in(far_3_3081_1[0]), .out(far_3_3081_2[0]));    relay_conn far_3_3081_2_b(.in(far_3_3081_1[1]), .out(far_3_3081_2[1]));
    assign layer_3[21] = ~far_3_3081_2[0] | (far_3_3081_2[0] & far_3_3081_2[1]); 
    assign layer_3[22] = ~(layer_2[374] | layer_2[361]); 
    wire [1:0] far_3_3083_0;    relay_conn far_3_3083_0_a(.in(layer_2[599]), .out(far_3_3083_0[0]));    relay_conn far_3_3083_0_b(.in(layer_2[635]), .out(far_3_3083_0[1]));
    assign layer_3[23] = far_3_3083_0[1] & ~far_3_3083_0[0]; 
    wire [1:0] far_3_3084_0;    relay_conn far_3_3084_0_a(.in(layer_2[613]), .out(far_3_3084_0[0]));    relay_conn far_3_3084_0_b(.in(layer_2[652]), .out(far_3_3084_0[1]));
    assign layer_3[24] = far_3_3084_0[0] & far_3_3084_0[1]; 
    wire [1:0] far_3_3085_0;    relay_conn far_3_3085_0_a(.in(layer_2[942]), .out(far_3_3085_0[0]));    relay_conn far_3_3085_0_b(.in(layer_2[996]), .out(far_3_3085_0[1]));
    assign layer_3[25] = ~(far_3_3085_0[0] & far_3_3085_0[1]); 
    wire [1:0] far_3_3086_0;    relay_conn far_3_3086_0_a(.in(layer_2[823]), .out(far_3_3086_0[0]));    relay_conn far_3_3086_0_b(.in(layer_2[920]), .out(far_3_3086_0[1]));
    wire [1:0] far_3_3086_1;    relay_conn far_3_3086_1_a(.in(far_3_3086_0[0]), .out(far_3_3086_1[0]));    relay_conn far_3_3086_1_b(.in(far_3_3086_0[1]), .out(far_3_3086_1[1]));
    wire [1:0] far_3_3086_2;    relay_conn far_3_3086_2_a(.in(far_3_3086_1[0]), .out(far_3_3086_2[0]));    relay_conn far_3_3086_2_b(.in(far_3_3086_1[1]), .out(far_3_3086_2[1]));
    assign layer_3[26] = far_3_3086_2[0] & ~far_3_3086_2[1]; 
    assign layer_3[27] = layer_2[276] | layer_2[248]; 
    assign layer_3[28] = layer_2[420] & ~layer_2[431]; 
    assign layer_3[29] = layer_2[624] ^ layer_2[593]; 
    wire [1:0] far_3_3090_0;    relay_conn far_3_3090_0_a(.in(layer_2[877]), .out(far_3_3090_0[0]));    relay_conn far_3_3090_0_b(.in(layer_2[956]), .out(far_3_3090_0[1]));
    wire [1:0] far_3_3090_1;    relay_conn far_3_3090_1_a(.in(far_3_3090_0[0]), .out(far_3_3090_1[0]));    relay_conn far_3_3090_1_b(.in(far_3_3090_0[1]), .out(far_3_3090_1[1]));
    assign layer_3[30] = ~(far_3_3090_1[0] & far_3_3090_1[1]); 
    assign layer_3[31] = layer_2[812] & layer_2[781]; 
    wire [1:0] far_3_3092_0;    relay_conn far_3_3092_0_a(.in(layer_2[237]), .out(far_3_3092_0[0]));    relay_conn far_3_3092_0_b(.in(layer_2[327]), .out(far_3_3092_0[1]));
    wire [1:0] far_3_3092_1;    relay_conn far_3_3092_1_a(.in(far_3_3092_0[0]), .out(far_3_3092_1[0]));    relay_conn far_3_3092_1_b(.in(far_3_3092_0[1]), .out(far_3_3092_1[1]));
    assign layer_3[32] = far_3_3092_1[1]; 
    assign layer_3[33] = ~layer_2[421]; 
    wire [1:0] far_3_3094_0;    relay_conn far_3_3094_0_a(.in(layer_2[992]), .out(far_3_3094_0[0]));    relay_conn far_3_3094_0_b(.in(layer_2[933]), .out(far_3_3094_0[1]));
    assign layer_3[34] = ~far_3_3094_0[1]; 
    wire [1:0] far_3_3095_0;    relay_conn far_3_3095_0_a(.in(layer_2[242]), .out(far_3_3095_0[0]));    relay_conn far_3_3095_0_b(.in(layer_2[191]), .out(far_3_3095_0[1]));
    assign layer_3[35] = far_3_3095_0[1] & ~far_3_3095_0[0]; 
    wire [1:0] far_3_3096_0;    relay_conn far_3_3096_0_a(.in(layer_2[299]), .out(far_3_3096_0[0]));    relay_conn far_3_3096_0_b(.in(layer_2[179]), .out(far_3_3096_0[1]));
    wire [1:0] far_3_3096_1;    relay_conn far_3_3096_1_a(.in(far_3_3096_0[0]), .out(far_3_3096_1[0]));    relay_conn far_3_3096_1_b(.in(far_3_3096_0[1]), .out(far_3_3096_1[1]));
    wire [1:0] far_3_3096_2;    relay_conn far_3_3096_2_a(.in(far_3_3096_1[0]), .out(far_3_3096_2[0]));    relay_conn far_3_3096_2_b(.in(far_3_3096_1[1]), .out(far_3_3096_2[1]));
    assign layer_3[36] = far_3_3096_2[0] & far_3_3096_2[1]; 
    wire [1:0] far_3_3097_0;    relay_conn far_3_3097_0_a(.in(layer_2[130]), .out(far_3_3097_0[0]));    relay_conn far_3_3097_0_b(.in(layer_2[95]), .out(far_3_3097_0[1]));
    assign layer_3[37] = far_3_3097_0[0] | far_3_3097_0[1]; 
    wire [1:0] far_3_3098_0;    relay_conn far_3_3098_0_a(.in(layer_2[716]), .out(far_3_3098_0[0]));    relay_conn far_3_3098_0_b(.in(layer_2[765]), .out(far_3_3098_0[1]));
    assign layer_3[38] = far_3_3098_0[0] | far_3_3098_0[1]; 
    wire [1:0] far_3_3099_0;    relay_conn far_3_3099_0_a(.in(layer_2[383]), .out(far_3_3099_0[0]));    relay_conn far_3_3099_0_b(.in(layer_2[330]), .out(far_3_3099_0[1]));
    assign layer_3[39] = far_3_3099_0[0] | far_3_3099_0[1]; 
    wire [1:0] far_3_3100_0;    relay_conn far_3_3100_0_a(.in(layer_2[1004]), .out(far_3_3100_0[0]));    relay_conn far_3_3100_0_b(.in(layer_2[925]), .out(far_3_3100_0[1]));
    wire [1:0] far_3_3100_1;    relay_conn far_3_3100_1_a(.in(far_3_3100_0[0]), .out(far_3_3100_1[0]));    relay_conn far_3_3100_1_b(.in(far_3_3100_0[1]), .out(far_3_3100_1[1]));
    assign layer_3[40] = ~far_3_3100_1[0] | (far_3_3100_1[0] & far_3_3100_1[1]); 
    wire [1:0] far_3_3101_0;    relay_conn far_3_3101_0_a(.in(layer_2[424]), .out(far_3_3101_0[0]));    relay_conn far_3_3101_0_b(.in(layer_2[546]), .out(far_3_3101_0[1]));
    wire [1:0] far_3_3101_1;    relay_conn far_3_3101_1_a(.in(far_3_3101_0[0]), .out(far_3_3101_1[0]));    relay_conn far_3_3101_1_b(.in(far_3_3101_0[1]), .out(far_3_3101_1[1]));
    wire [1:0] far_3_3101_2;    relay_conn far_3_3101_2_a(.in(far_3_3101_1[0]), .out(far_3_3101_2[0]));    relay_conn far_3_3101_2_b(.in(far_3_3101_1[1]), .out(far_3_3101_2[1]));
    assign layer_3[41] = ~far_3_3101_2[1] | (far_3_3101_2[0] & far_3_3101_2[1]); 
    wire [1:0] far_3_3102_0;    relay_conn far_3_3102_0_a(.in(layer_2[896]), .out(far_3_3102_0[0]));    relay_conn far_3_3102_0_b(.in(layer_2[858]), .out(far_3_3102_0[1]));
    assign layer_3[42] = far_3_3102_0[0] | far_3_3102_0[1]; 
    assign layer_3[43] = ~layer_2[763]; 
    assign layer_3[44] = ~(layer_2[902] & layer_2[891]); 
    assign layer_3[45] = layer_2[878]; 
    wire [1:0] far_3_3106_0;    relay_conn far_3_3106_0_a(.in(layer_2[382]), .out(far_3_3106_0[0]));    relay_conn far_3_3106_0_b(.in(layer_2[433]), .out(far_3_3106_0[1]));
    assign layer_3[46] = far_3_3106_0[0] | far_3_3106_0[1]; 
    wire [1:0] far_3_3107_0;    relay_conn far_3_3107_0_a(.in(layer_2[126]), .out(far_3_3107_0[0]));    relay_conn far_3_3107_0_b(.in(layer_2[12]), .out(far_3_3107_0[1]));
    wire [1:0] far_3_3107_1;    relay_conn far_3_3107_1_a(.in(far_3_3107_0[0]), .out(far_3_3107_1[0]));    relay_conn far_3_3107_1_b(.in(far_3_3107_0[1]), .out(far_3_3107_1[1]));
    wire [1:0] far_3_3107_2;    relay_conn far_3_3107_2_a(.in(far_3_3107_1[0]), .out(far_3_3107_2[0]));    relay_conn far_3_3107_2_b(.in(far_3_3107_1[1]), .out(far_3_3107_2[1]));
    assign layer_3[47] = ~far_3_3107_2[1]; 
    wire [1:0] far_3_3108_0;    relay_conn far_3_3108_0_a(.in(layer_2[663]), .out(far_3_3108_0[0]));    relay_conn far_3_3108_0_b(.in(layer_2[592]), .out(far_3_3108_0[1]));
    wire [1:0] far_3_3108_1;    relay_conn far_3_3108_1_a(.in(far_3_3108_0[0]), .out(far_3_3108_1[0]));    relay_conn far_3_3108_1_b(.in(far_3_3108_0[1]), .out(far_3_3108_1[1]));
    assign layer_3[48] = far_3_3108_1[0]; 
    wire [1:0] far_3_3109_0;    relay_conn far_3_3109_0_a(.in(layer_2[175]), .out(far_3_3109_0[0]));    relay_conn far_3_3109_0_b(.in(layer_2[100]), .out(far_3_3109_0[1]));
    wire [1:0] far_3_3109_1;    relay_conn far_3_3109_1_a(.in(far_3_3109_0[0]), .out(far_3_3109_1[0]));    relay_conn far_3_3109_1_b(.in(far_3_3109_0[1]), .out(far_3_3109_1[1]));
    assign layer_3[49] = far_3_3109_1[1] & ~far_3_3109_1[0]; 
    wire [1:0] far_3_3110_0;    relay_conn far_3_3110_0_a(.in(layer_2[658]), .out(far_3_3110_0[0]));    relay_conn far_3_3110_0_b(.in(layer_2[558]), .out(far_3_3110_0[1]));
    wire [1:0] far_3_3110_1;    relay_conn far_3_3110_1_a(.in(far_3_3110_0[0]), .out(far_3_3110_1[0]));    relay_conn far_3_3110_1_b(.in(far_3_3110_0[1]), .out(far_3_3110_1[1]));
    wire [1:0] far_3_3110_2;    relay_conn far_3_3110_2_a(.in(far_3_3110_1[0]), .out(far_3_3110_2[0]));    relay_conn far_3_3110_2_b(.in(far_3_3110_1[1]), .out(far_3_3110_2[1]));
    assign layer_3[50] = far_3_3110_2[0] & far_3_3110_2[1]; 
    wire [1:0] far_3_3111_0;    relay_conn far_3_3111_0_a(.in(layer_2[508]), .out(far_3_3111_0[0]));    relay_conn far_3_3111_0_b(.in(layer_2[445]), .out(far_3_3111_0[1]));
    assign layer_3[51] = far_3_3111_0[0] | far_3_3111_0[1]; 
    wire [1:0] far_3_3112_0;    relay_conn far_3_3112_0_a(.in(layer_2[886]), .out(far_3_3112_0[0]));    relay_conn far_3_3112_0_b(.in(layer_2[949]), .out(far_3_3112_0[1]));
    assign layer_3[52] = ~far_3_3112_0[0] | (far_3_3112_0[0] & far_3_3112_0[1]); 
    assign layer_3[53] = ~layer_2[640]; 
    wire [1:0] far_3_3114_0;    relay_conn far_3_3114_0_a(.in(layer_2[444]), .out(far_3_3114_0[0]));    relay_conn far_3_3114_0_b(.in(layer_2[516]), .out(far_3_3114_0[1]));
    wire [1:0] far_3_3114_1;    relay_conn far_3_3114_1_a(.in(far_3_3114_0[0]), .out(far_3_3114_1[0]));    relay_conn far_3_3114_1_b(.in(far_3_3114_0[1]), .out(far_3_3114_1[1]));
    assign layer_3[54] = far_3_3114_1[0]; 
    wire [1:0] far_3_3115_0;    relay_conn far_3_3115_0_a(.in(layer_2[778]), .out(far_3_3115_0[0]));    relay_conn far_3_3115_0_b(.in(layer_2[678]), .out(far_3_3115_0[1]));
    wire [1:0] far_3_3115_1;    relay_conn far_3_3115_1_a(.in(far_3_3115_0[0]), .out(far_3_3115_1[0]));    relay_conn far_3_3115_1_b(.in(far_3_3115_0[1]), .out(far_3_3115_1[1]));
    wire [1:0] far_3_3115_2;    relay_conn far_3_3115_2_a(.in(far_3_3115_1[0]), .out(far_3_3115_2[0]));    relay_conn far_3_3115_2_b(.in(far_3_3115_1[1]), .out(far_3_3115_2[1]));
    assign layer_3[55] = far_3_3115_2[0] & far_3_3115_2[1]; 
    assign layer_3[56] = layer_2[825] & ~layer_2[837]; 
    wire [1:0] far_3_3117_0;    relay_conn far_3_3117_0_a(.in(layer_2[223]), .out(far_3_3117_0[0]));    relay_conn far_3_3117_0_b(.in(layer_2[299]), .out(far_3_3117_0[1]));
    wire [1:0] far_3_3117_1;    relay_conn far_3_3117_1_a(.in(far_3_3117_0[0]), .out(far_3_3117_1[0]));    relay_conn far_3_3117_1_b(.in(far_3_3117_0[1]), .out(far_3_3117_1[1]));
    assign layer_3[57] = far_3_3117_1[0] & ~far_3_3117_1[1]; 
    wire [1:0] far_3_3118_0;    relay_conn far_3_3118_0_a(.in(layer_2[422]), .out(far_3_3118_0[0]));    relay_conn far_3_3118_0_b(.in(layer_2[306]), .out(far_3_3118_0[1]));
    wire [1:0] far_3_3118_1;    relay_conn far_3_3118_1_a(.in(far_3_3118_0[0]), .out(far_3_3118_1[0]));    relay_conn far_3_3118_1_b(.in(far_3_3118_0[1]), .out(far_3_3118_1[1]));
    wire [1:0] far_3_3118_2;    relay_conn far_3_3118_2_a(.in(far_3_3118_1[0]), .out(far_3_3118_2[0]));    relay_conn far_3_3118_2_b(.in(far_3_3118_1[1]), .out(far_3_3118_2[1]));
    assign layer_3[58] = ~far_3_3118_2[0] | (far_3_3118_2[0] & far_3_3118_2[1]); 
    assign layer_3[59] = layer_2[345] & ~layer_2[364]; 
    assign layer_3[60] = layer_2[429] & ~layer_2[433]; 
    wire [1:0] far_3_3121_0;    relay_conn far_3_3121_0_a(.in(layer_2[464]), .out(far_3_3121_0[0]));    relay_conn far_3_3121_0_b(.in(layer_2[578]), .out(far_3_3121_0[1]));
    wire [1:0] far_3_3121_1;    relay_conn far_3_3121_1_a(.in(far_3_3121_0[0]), .out(far_3_3121_1[0]));    relay_conn far_3_3121_1_b(.in(far_3_3121_0[1]), .out(far_3_3121_1[1]));
    wire [1:0] far_3_3121_2;    relay_conn far_3_3121_2_a(.in(far_3_3121_1[0]), .out(far_3_3121_2[0]));    relay_conn far_3_3121_2_b(.in(far_3_3121_1[1]), .out(far_3_3121_2[1]));
    assign layer_3[61] = ~(far_3_3121_2[0] & far_3_3121_2[1]); 
    assign layer_3[62] = ~layer_2[925]; 
    wire [1:0] far_3_3123_0;    relay_conn far_3_3123_0_a(.in(layer_2[414]), .out(far_3_3123_0[0]));    relay_conn far_3_3123_0_b(.in(layer_2[288]), .out(far_3_3123_0[1]));
    wire [1:0] far_3_3123_1;    relay_conn far_3_3123_1_a(.in(far_3_3123_0[0]), .out(far_3_3123_1[0]));    relay_conn far_3_3123_1_b(.in(far_3_3123_0[1]), .out(far_3_3123_1[1]));
    wire [1:0] far_3_3123_2;    relay_conn far_3_3123_2_a(.in(far_3_3123_1[0]), .out(far_3_3123_2[0]));    relay_conn far_3_3123_2_b(.in(far_3_3123_1[1]), .out(far_3_3123_2[1]));
    assign layer_3[63] = ~far_3_3123_2[0]; 
    assign layer_3[64] = ~layer_2[452]; 
    assign layer_3[65] = ~(layer_2[784] | layer_2[790]); 
    wire [1:0] far_3_3126_0;    relay_conn far_3_3126_0_a(.in(layer_2[646]), .out(far_3_3126_0[0]));    relay_conn far_3_3126_0_b(.in(layer_2[562]), .out(far_3_3126_0[1]));
    wire [1:0] far_3_3126_1;    relay_conn far_3_3126_1_a(.in(far_3_3126_0[0]), .out(far_3_3126_1[0]));    relay_conn far_3_3126_1_b(.in(far_3_3126_0[1]), .out(far_3_3126_1[1]));
    assign layer_3[66] = ~far_3_3126_1[0]; 
    wire [1:0] far_3_3127_0;    relay_conn far_3_3127_0_a(.in(layer_2[965]), .out(far_3_3127_0[0]));    relay_conn far_3_3127_0_b(.in(layer_2[843]), .out(far_3_3127_0[1]));
    wire [1:0] far_3_3127_1;    relay_conn far_3_3127_1_a(.in(far_3_3127_0[0]), .out(far_3_3127_1[0]));    relay_conn far_3_3127_1_b(.in(far_3_3127_0[1]), .out(far_3_3127_1[1]));
    wire [1:0] far_3_3127_2;    relay_conn far_3_3127_2_a(.in(far_3_3127_1[0]), .out(far_3_3127_2[0]));    relay_conn far_3_3127_2_b(.in(far_3_3127_1[1]), .out(far_3_3127_2[1]));
    assign layer_3[67] = ~far_3_3127_2[1] | (far_3_3127_2[0] & far_3_3127_2[1]); 
    wire [1:0] far_3_3128_0;    relay_conn far_3_3128_0_a(.in(layer_2[992]), .out(far_3_3128_0[0]));    relay_conn far_3_3128_0_b(.in(layer_2[949]), .out(far_3_3128_0[1]));
    assign layer_3[68] = ~far_3_3128_0[1]; 
    assign layer_3[69] = layer_2[865] ^ layer_2[839]; 
    assign layer_3[70] = ~(layer_2[138] & layer_2[151]); 
    wire [1:0] far_3_3131_0;    relay_conn far_3_3131_0_a(.in(layer_2[385]), .out(far_3_3131_0[0]));    relay_conn far_3_3131_0_b(.in(layer_2[330]), .out(far_3_3131_0[1]));
    assign layer_3[71] = far_3_3131_0[0] & far_3_3131_0[1]; 
    wire [1:0] far_3_3132_0;    relay_conn far_3_3132_0_a(.in(layer_2[832]), .out(far_3_3132_0[0]));    relay_conn far_3_3132_0_b(.in(layer_2[905]), .out(far_3_3132_0[1]));
    wire [1:0] far_3_3132_1;    relay_conn far_3_3132_1_a(.in(far_3_3132_0[0]), .out(far_3_3132_1[0]));    relay_conn far_3_3132_1_b(.in(far_3_3132_0[1]), .out(far_3_3132_1[1]));
    assign layer_3[72] = ~far_3_3132_1[0] | (far_3_3132_1[0] & far_3_3132_1[1]); 
    wire [1:0] far_3_3133_0;    relay_conn far_3_3133_0_a(.in(layer_2[519]), .out(far_3_3133_0[0]));    relay_conn far_3_3133_0_b(.in(layer_2[590]), .out(far_3_3133_0[1]));
    wire [1:0] far_3_3133_1;    relay_conn far_3_3133_1_a(.in(far_3_3133_0[0]), .out(far_3_3133_1[0]));    relay_conn far_3_3133_1_b(.in(far_3_3133_0[1]), .out(far_3_3133_1[1]));
    assign layer_3[73] = far_3_3133_1[0] & ~far_3_3133_1[1]; 
    wire [1:0] far_3_3134_0;    relay_conn far_3_3134_0_a(.in(layer_2[212]), .out(far_3_3134_0[0]));    relay_conn far_3_3134_0_b(.in(layer_2[292]), .out(far_3_3134_0[1]));
    wire [1:0] far_3_3134_1;    relay_conn far_3_3134_1_a(.in(far_3_3134_0[0]), .out(far_3_3134_1[0]));    relay_conn far_3_3134_1_b(.in(far_3_3134_0[1]), .out(far_3_3134_1[1]));
    assign layer_3[74] = ~far_3_3134_1[0]; 
    wire [1:0] far_3_3135_0;    relay_conn far_3_3135_0_a(.in(layer_2[92]), .out(far_3_3135_0[0]));    relay_conn far_3_3135_0_b(.in(layer_2[170]), .out(far_3_3135_0[1]));
    wire [1:0] far_3_3135_1;    relay_conn far_3_3135_1_a(.in(far_3_3135_0[0]), .out(far_3_3135_1[0]));    relay_conn far_3_3135_1_b(.in(far_3_3135_0[1]), .out(far_3_3135_1[1]));
    assign layer_3[75] = far_3_3135_1[0] & far_3_3135_1[1]; 
    wire [1:0] far_3_3136_0;    relay_conn far_3_3136_0_a(.in(layer_2[408]), .out(far_3_3136_0[0]));    relay_conn far_3_3136_0_b(.in(layer_2[520]), .out(far_3_3136_0[1]));
    wire [1:0] far_3_3136_1;    relay_conn far_3_3136_1_a(.in(far_3_3136_0[0]), .out(far_3_3136_1[0]));    relay_conn far_3_3136_1_b(.in(far_3_3136_0[1]), .out(far_3_3136_1[1]));
    wire [1:0] far_3_3136_2;    relay_conn far_3_3136_2_a(.in(far_3_3136_1[0]), .out(far_3_3136_2[0]));    relay_conn far_3_3136_2_b(.in(far_3_3136_1[1]), .out(far_3_3136_2[1]));
    assign layer_3[76] = ~(far_3_3136_2[0] & far_3_3136_2[1]); 
    wire [1:0] far_3_3137_0;    relay_conn far_3_3137_0_a(.in(layer_2[927]), .out(far_3_3137_0[0]));    relay_conn far_3_3137_0_b(.in(layer_2[878]), .out(far_3_3137_0[1]));
    assign layer_3[77] = ~far_3_3137_0[1]; 
    assign layer_3[78] = layer_2[505] & ~layer_2[509]; 
    wire [1:0] far_3_3139_0;    relay_conn far_3_3139_0_a(.in(layer_2[379]), .out(far_3_3139_0[0]));    relay_conn far_3_3139_0_b(.in(layer_2[307]), .out(far_3_3139_0[1]));
    wire [1:0] far_3_3139_1;    relay_conn far_3_3139_1_a(.in(far_3_3139_0[0]), .out(far_3_3139_1[0]));    relay_conn far_3_3139_1_b(.in(far_3_3139_0[1]), .out(far_3_3139_1[1]));
    assign layer_3[79] = far_3_3139_1[0] ^ far_3_3139_1[1]; 
    wire [1:0] far_3_3140_0;    relay_conn far_3_3140_0_a(.in(layer_2[8]), .out(far_3_3140_0[0]));    relay_conn far_3_3140_0_b(.in(layer_2[132]), .out(far_3_3140_0[1]));
    wire [1:0] far_3_3140_1;    relay_conn far_3_3140_1_a(.in(far_3_3140_0[0]), .out(far_3_3140_1[0]));    relay_conn far_3_3140_1_b(.in(far_3_3140_0[1]), .out(far_3_3140_1[1]));
    wire [1:0] far_3_3140_2;    relay_conn far_3_3140_2_a(.in(far_3_3140_1[0]), .out(far_3_3140_2[0]));    relay_conn far_3_3140_2_b(.in(far_3_3140_1[1]), .out(far_3_3140_2[1]));
    assign layer_3[80] = far_3_3140_2[0]; 
    wire [1:0] far_3_3141_0;    relay_conn far_3_3141_0_a(.in(layer_2[112]), .out(far_3_3141_0[0]));    relay_conn far_3_3141_0_b(.in(layer_2[5]), .out(far_3_3141_0[1]));
    wire [1:0] far_3_3141_1;    relay_conn far_3_3141_1_a(.in(far_3_3141_0[0]), .out(far_3_3141_1[0]));    relay_conn far_3_3141_1_b(.in(far_3_3141_0[1]), .out(far_3_3141_1[1]));
    wire [1:0] far_3_3141_2;    relay_conn far_3_3141_2_a(.in(far_3_3141_1[0]), .out(far_3_3141_2[0]));    relay_conn far_3_3141_2_b(.in(far_3_3141_1[1]), .out(far_3_3141_2[1]));
    assign layer_3[81] = far_3_3141_2[1] & ~far_3_3141_2[0]; 
    wire [1:0] far_3_3142_0;    relay_conn far_3_3142_0_a(.in(layer_2[509]), .out(far_3_3142_0[0]));    relay_conn far_3_3142_0_b(.in(layer_2[440]), .out(far_3_3142_0[1]));
    wire [1:0] far_3_3142_1;    relay_conn far_3_3142_1_a(.in(far_3_3142_0[0]), .out(far_3_3142_1[0]));    relay_conn far_3_3142_1_b(.in(far_3_3142_0[1]), .out(far_3_3142_1[1]));
    assign layer_3[82] = ~far_3_3142_1[1] | (far_3_3142_1[0] & far_3_3142_1[1]); 
    wire [1:0] far_3_3143_0;    relay_conn far_3_3143_0_a(.in(layer_2[809]), .out(far_3_3143_0[0]));    relay_conn far_3_3143_0_b(.in(layer_2[878]), .out(far_3_3143_0[1]));
    wire [1:0] far_3_3143_1;    relay_conn far_3_3143_1_a(.in(far_3_3143_0[0]), .out(far_3_3143_1[0]));    relay_conn far_3_3143_1_b(.in(far_3_3143_0[1]), .out(far_3_3143_1[1]));
    assign layer_3[83] = ~far_3_3143_1[0] | (far_3_3143_1[0] & far_3_3143_1[1]); 
    wire [1:0] far_3_3144_0;    relay_conn far_3_3144_0_a(.in(layer_2[244]), .out(far_3_3144_0[0]));    relay_conn far_3_3144_0_b(.in(layer_2[134]), .out(far_3_3144_0[1]));
    wire [1:0] far_3_3144_1;    relay_conn far_3_3144_1_a(.in(far_3_3144_0[0]), .out(far_3_3144_1[0]));    relay_conn far_3_3144_1_b(.in(far_3_3144_0[1]), .out(far_3_3144_1[1]));
    wire [1:0] far_3_3144_2;    relay_conn far_3_3144_2_a(.in(far_3_3144_1[0]), .out(far_3_3144_2[0]));    relay_conn far_3_3144_2_b(.in(far_3_3144_1[1]), .out(far_3_3144_2[1]));
    assign layer_3[84] = ~far_3_3144_2[0]; 
    assign layer_3[85] = ~layer_2[3] | (layer_2[3] & layer_2[2]); 
    wire [1:0] far_3_3146_0;    relay_conn far_3_3146_0_a(.in(layer_2[326]), .out(far_3_3146_0[0]));    relay_conn far_3_3146_0_b(.in(layer_2[219]), .out(far_3_3146_0[1]));
    wire [1:0] far_3_3146_1;    relay_conn far_3_3146_1_a(.in(far_3_3146_0[0]), .out(far_3_3146_1[0]));    relay_conn far_3_3146_1_b(.in(far_3_3146_0[1]), .out(far_3_3146_1[1]));
    wire [1:0] far_3_3146_2;    relay_conn far_3_3146_2_a(.in(far_3_3146_1[0]), .out(far_3_3146_2[0]));    relay_conn far_3_3146_2_b(.in(far_3_3146_1[1]), .out(far_3_3146_2[1]));
    assign layer_3[86] = far_3_3146_2[0] ^ far_3_3146_2[1]; 
    assign layer_3[87] = ~layer_2[360] | (layer_2[360] & layer_2[347]); 
    wire [1:0] far_3_3148_0;    relay_conn far_3_3148_0_a(.in(layer_2[843]), .out(far_3_3148_0[0]));    relay_conn far_3_3148_0_b(.in(layer_2[781]), .out(far_3_3148_0[1]));
    assign layer_3[88] = far_3_3148_0[1] & ~far_3_3148_0[0]; 
    wire [1:0] far_3_3149_0;    relay_conn far_3_3149_0_a(.in(layer_2[348]), .out(far_3_3149_0[0]));    relay_conn far_3_3149_0_b(.in(layer_2[244]), .out(far_3_3149_0[1]));
    wire [1:0] far_3_3149_1;    relay_conn far_3_3149_1_a(.in(far_3_3149_0[0]), .out(far_3_3149_1[0]));    relay_conn far_3_3149_1_b(.in(far_3_3149_0[1]), .out(far_3_3149_1[1]));
    wire [1:0] far_3_3149_2;    relay_conn far_3_3149_2_a(.in(far_3_3149_1[0]), .out(far_3_3149_2[0]));    relay_conn far_3_3149_2_b(.in(far_3_3149_1[1]), .out(far_3_3149_2[1]));
    assign layer_3[89] = ~(far_3_3149_2[0] ^ far_3_3149_2[1]); 
    wire [1:0] far_3_3150_0;    relay_conn far_3_3150_0_a(.in(layer_2[268]), .out(far_3_3150_0[0]));    relay_conn far_3_3150_0_b(.in(layer_2[354]), .out(far_3_3150_0[1]));
    wire [1:0] far_3_3150_1;    relay_conn far_3_3150_1_a(.in(far_3_3150_0[0]), .out(far_3_3150_1[0]));    relay_conn far_3_3150_1_b(.in(far_3_3150_0[1]), .out(far_3_3150_1[1]));
    assign layer_3[90] = ~far_3_3150_1[0] | (far_3_3150_1[0] & far_3_3150_1[1]); 
    wire [1:0] far_3_3151_0;    relay_conn far_3_3151_0_a(.in(layer_2[539]), .out(far_3_3151_0[0]));    relay_conn far_3_3151_0_b(.in(layer_2[504]), .out(far_3_3151_0[1]));
    assign layer_3[91] = far_3_3151_0[1]; 
    assign layer_3[92] = ~(layer_2[175] & layer_2[151]); 
    wire [1:0] far_3_3153_0;    relay_conn far_3_3153_0_a(.in(layer_2[733]), .out(far_3_3153_0[0]));    relay_conn far_3_3153_0_b(.in(layer_2[835]), .out(far_3_3153_0[1]));
    wire [1:0] far_3_3153_1;    relay_conn far_3_3153_1_a(.in(far_3_3153_0[0]), .out(far_3_3153_1[0]));    relay_conn far_3_3153_1_b(.in(far_3_3153_0[1]), .out(far_3_3153_1[1]));
    wire [1:0] far_3_3153_2;    relay_conn far_3_3153_2_a(.in(far_3_3153_1[0]), .out(far_3_3153_2[0]));    relay_conn far_3_3153_2_b(.in(far_3_3153_1[1]), .out(far_3_3153_2[1]));
    assign layer_3[93] = ~far_3_3153_2[0]; 
    assign layer_3[94] = layer_2[48] & layer_2[58]; 
    wire [1:0] far_3_3155_0;    relay_conn far_3_3155_0_a(.in(layer_2[284]), .out(far_3_3155_0[0]));    relay_conn far_3_3155_0_b(.in(layer_2[250]), .out(far_3_3155_0[1]));
    assign layer_3[95] = ~far_3_3155_0[1] | (far_3_3155_0[0] & far_3_3155_0[1]); 
    assign layer_3[96] = layer_2[583] | layer_2[604]; 
    wire [1:0] far_3_3157_0;    relay_conn far_3_3157_0_a(.in(layer_2[252]), .out(far_3_3157_0[0]));    relay_conn far_3_3157_0_b(.in(layer_2[345]), .out(far_3_3157_0[1]));
    wire [1:0] far_3_3157_1;    relay_conn far_3_3157_1_a(.in(far_3_3157_0[0]), .out(far_3_3157_1[0]));    relay_conn far_3_3157_1_b(.in(far_3_3157_0[1]), .out(far_3_3157_1[1]));
    assign layer_3[97] = far_3_3157_1[0] & far_3_3157_1[1]; 
    wire [1:0] far_3_3158_0;    relay_conn far_3_3158_0_a(.in(layer_2[151]), .out(far_3_3158_0[0]));    relay_conn far_3_3158_0_b(.in(layer_2[216]), .out(far_3_3158_0[1]));
    wire [1:0] far_3_3158_1;    relay_conn far_3_3158_1_a(.in(far_3_3158_0[0]), .out(far_3_3158_1[0]));    relay_conn far_3_3158_1_b(.in(far_3_3158_0[1]), .out(far_3_3158_1[1]));
    assign layer_3[98] = far_3_3158_1[1]; 
    wire [1:0] far_3_3159_0;    relay_conn far_3_3159_0_a(.in(layer_2[453]), .out(far_3_3159_0[0]));    relay_conn far_3_3159_0_b(.in(layer_2[546]), .out(far_3_3159_0[1]));
    wire [1:0] far_3_3159_1;    relay_conn far_3_3159_1_a(.in(far_3_3159_0[0]), .out(far_3_3159_1[0]));    relay_conn far_3_3159_1_b(.in(far_3_3159_0[1]), .out(far_3_3159_1[1]));
    assign layer_3[99] = far_3_3159_1[1]; 
    wire [1:0] far_3_3160_0;    relay_conn far_3_3160_0_a(.in(layer_2[565]), .out(far_3_3160_0[0]));    relay_conn far_3_3160_0_b(.in(layer_2[522]), .out(far_3_3160_0[1]));
    assign layer_3[100] = ~far_3_3160_0[1] | (far_3_3160_0[0] & far_3_3160_0[1]); 
    wire [1:0] far_3_3161_0;    relay_conn far_3_3161_0_a(.in(layer_2[946]), .out(far_3_3161_0[0]));    relay_conn far_3_3161_0_b(.in(layer_2[910]), .out(far_3_3161_0[1]));
    assign layer_3[101] = far_3_3161_0[0] & far_3_3161_0[1]; 
    wire [1:0] far_3_3162_0;    relay_conn far_3_3162_0_a(.in(layer_2[208]), .out(far_3_3162_0[0]));    relay_conn far_3_3162_0_b(.in(layer_2[100]), .out(far_3_3162_0[1]));
    wire [1:0] far_3_3162_1;    relay_conn far_3_3162_1_a(.in(far_3_3162_0[0]), .out(far_3_3162_1[0]));    relay_conn far_3_3162_1_b(.in(far_3_3162_0[1]), .out(far_3_3162_1[1]));
    wire [1:0] far_3_3162_2;    relay_conn far_3_3162_2_a(.in(far_3_3162_1[0]), .out(far_3_3162_2[0]));    relay_conn far_3_3162_2_b(.in(far_3_3162_1[1]), .out(far_3_3162_2[1]));
    assign layer_3[102] = ~far_3_3162_2[1]; 
    wire [1:0] far_3_3163_0;    relay_conn far_3_3163_0_a(.in(layer_2[528]), .out(far_3_3163_0[0]));    relay_conn far_3_3163_0_b(.in(layer_2[654]), .out(far_3_3163_0[1]));
    wire [1:0] far_3_3163_1;    relay_conn far_3_3163_1_a(.in(far_3_3163_0[0]), .out(far_3_3163_1[0]));    relay_conn far_3_3163_1_b(.in(far_3_3163_0[1]), .out(far_3_3163_1[1]));
    wire [1:0] far_3_3163_2;    relay_conn far_3_3163_2_a(.in(far_3_3163_1[0]), .out(far_3_3163_2[0]));    relay_conn far_3_3163_2_b(.in(far_3_3163_1[1]), .out(far_3_3163_2[1]));
    assign layer_3[103] = ~far_3_3163_2[1] | (far_3_3163_2[0] & far_3_3163_2[1]); 
    wire [1:0] far_3_3164_0;    relay_conn far_3_3164_0_a(.in(layer_2[479]), .out(far_3_3164_0[0]));    relay_conn far_3_3164_0_b(.in(layer_2[425]), .out(far_3_3164_0[1]));
    assign layer_3[104] = ~(far_3_3164_0[0] & far_3_3164_0[1]); 
    wire [1:0] far_3_3165_0;    relay_conn far_3_3165_0_a(.in(layer_2[509]), .out(far_3_3165_0[0]));    relay_conn far_3_3165_0_b(.in(layer_2[468]), .out(far_3_3165_0[1]));
    assign layer_3[105] = ~(far_3_3165_0[0] | far_3_3165_0[1]); 
    assign layer_3[106] = layer_2[291] & ~layer_2[315]; 
    wire [1:0] far_3_3167_0;    relay_conn far_3_3167_0_a(.in(layer_2[433]), .out(far_3_3167_0[0]));    relay_conn far_3_3167_0_b(.in(layer_2[379]), .out(far_3_3167_0[1]));
    assign layer_3[107] = far_3_3167_0[1] & ~far_3_3167_0[0]; 
    assign layer_3[108] = ~(layer_2[103] & layer_2[92]); 
    wire [1:0] far_3_3169_0;    relay_conn far_3_3169_0_a(.in(layer_2[23]), .out(far_3_3169_0[0]));    relay_conn far_3_3169_0_b(.in(layer_2[84]), .out(far_3_3169_0[1]));
    assign layer_3[109] = far_3_3169_0[0] & far_3_3169_0[1]; 
    wire [1:0] far_3_3170_0;    relay_conn far_3_3170_0_a(.in(layer_2[666]), .out(far_3_3170_0[0]));    relay_conn far_3_3170_0_b(.in(layer_2[543]), .out(far_3_3170_0[1]));
    wire [1:0] far_3_3170_1;    relay_conn far_3_3170_1_a(.in(far_3_3170_0[0]), .out(far_3_3170_1[0]));    relay_conn far_3_3170_1_b(.in(far_3_3170_0[1]), .out(far_3_3170_1[1]));
    wire [1:0] far_3_3170_2;    relay_conn far_3_3170_2_a(.in(far_3_3170_1[0]), .out(far_3_3170_2[0]));    relay_conn far_3_3170_2_b(.in(far_3_3170_1[1]), .out(far_3_3170_2[1]));
    assign layer_3[110] = far_3_3170_2[0] & ~far_3_3170_2[1]; 
    wire [1:0] far_3_3171_0;    relay_conn far_3_3171_0_a(.in(layer_2[934]), .out(far_3_3171_0[0]));    relay_conn far_3_3171_0_b(.in(layer_2[867]), .out(far_3_3171_0[1]));
    wire [1:0] far_3_3171_1;    relay_conn far_3_3171_1_a(.in(far_3_3171_0[0]), .out(far_3_3171_1[0]));    relay_conn far_3_3171_1_b(.in(far_3_3171_0[1]), .out(far_3_3171_1[1]));
    assign layer_3[111] = ~far_3_3171_1[1] | (far_3_3171_1[0] & far_3_3171_1[1]); 
    assign layer_3[112] = layer_2[188] | layer_2[180]; 
    wire [1:0] far_3_3173_0;    relay_conn far_3_3173_0_a(.in(layer_2[504]), .out(far_3_3173_0[0]));    relay_conn far_3_3173_0_b(.in(layer_2[576]), .out(far_3_3173_0[1]));
    wire [1:0] far_3_3173_1;    relay_conn far_3_3173_1_a(.in(far_3_3173_0[0]), .out(far_3_3173_1[0]));    relay_conn far_3_3173_1_b(.in(far_3_3173_0[1]), .out(far_3_3173_1[1]));
    assign layer_3[113] = ~far_3_3173_1[0] | (far_3_3173_1[0] & far_3_3173_1[1]); 
    assign layer_3[114] = ~(layer_2[361] | layer_2[389]); 
    wire [1:0] far_3_3175_0;    relay_conn far_3_3175_0_a(.in(layer_2[843]), .out(far_3_3175_0[0]));    relay_conn far_3_3175_0_b(.in(layer_2[891]), .out(far_3_3175_0[1]));
    assign layer_3[115] = ~far_3_3175_0[0]; 
    wire [1:0] far_3_3176_0;    relay_conn far_3_3176_0_a(.in(layer_2[811]), .out(far_3_3176_0[0]));    relay_conn far_3_3176_0_b(.in(layer_2[875]), .out(far_3_3176_0[1]));
    wire [1:0] far_3_3176_1;    relay_conn far_3_3176_1_a(.in(far_3_3176_0[0]), .out(far_3_3176_1[0]));    relay_conn far_3_3176_1_b(.in(far_3_3176_0[1]), .out(far_3_3176_1[1]));
    assign layer_3[116] = far_3_3176_1[0] & far_3_3176_1[1]; 
    wire [1:0] far_3_3177_0;    relay_conn far_3_3177_0_a(.in(layer_2[154]), .out(far_3_3177_0[0]));    relay_conn far_3_3177_0_b(.in(layer_2[240]), .out(far_3_3177_0[1]));
    wire [1:0] far_3_3177_1;    relay_conn far_3_3177_1_a(.in(far_3_3177_0[0]), .out(far_3_3177_1[0]));    relay_conn far_3_3177_1_b(.in(far_3_3177_0[1]), .out(far_3_3177_1[1]));
    assign layer_3[117] = ~far_3_3177_1[0] | (far_3_3177_1[0] & far_3_3177_1[1]); 
    wire [1:0] far_3_3178_0;    relay_conn far_3_3178_0_a(.in(layer_2[194]), .out(far_3_3178_0[0]));    relay_conn far_3_3178_0_b(.in(layer_2[93]), .out(far_3_3178_0[1]));
    wire [1:0] far_3_3178_1;    relay_conn far_3_3178_1_a(.in(far_3_3178_0[0]), .out(far_3_3178_1[0]));    relay_conn far_3_3178_1_b(.in(far_3_3178_0[1]), .out(far_3_3178_1[1]));
    wire [1:0] far_3_3178_2;    relay_conn far_3_3178_2_a(.in(far_3_3178_1[0]), .out(far_3_3178_2[0]));    relay_conn far_3_3178_2_b(.in(far_3_3178_1[1]), .out(far_3_3178_2[1]));
    assign layer_3[118] = far_3_3178_2[1]; 
    assign layer_3[119] = ~layer_2[495]; 
    wire [1:0] far_3_3180_0;    relay_conn far_3_3180_0_a(.in(layer_2[645]), .out(far_3_3180_0[0]));    relay_conn far_3_3180_0_b(.in(layer_2[678]), .out(far_3_3180_0[1]));
    assign layer_3[120] = far_3_3180_0[1]; 
    wire [1:0] far_3_3181_0;    relay_conn far_3_3181_0_a(.in(layer_2[827]), .out(far_3_3181_0[0]));    relay_conn far_3_3181_0_b(.in(layer_2[774]), .out(far_3_3181_0[1]));
    assign layer_3[121] = ~far_3_3181_0[1] | (far_3_3181_0[0] & far_3_3181_0[1]); 
    wire [1:0] far_3_3182_0;    relay_conn far_3_3182_0_a(.in(layer_2[915]), .out(far_3_3182_0[0]));    relay_conn far_3_3182_0_b(.in(layer_2[811]), .out(far_3_3182_0[1]));
    wire [1:0] far_3_3182_1;    relay_conn far_3_3182_1_a(.in(far_3_3182_0[0]), .out(far_3_3182_1[0]));    relay_conn far_3_3182_1_b(.in(far_3_3182_0[1]), .out(far_3_3182_1[1]));
    wire [1:0] far_3_3182_2;    relay_conn far_3_3182_2_a(.in(far_3_3182_1[0]), .out(far_3_3182_2[0]));    relay_conn far_3_3182_2_b(.in(far_3_3182_1[1]), .out(far_3_3182_2[1]));
    assign layer_3[122] = far_3_3182_2[0] | far_3_3182_2[1]; 
    wire [1:0] far_3_3183_0;    relay_conn far_3_3183_0_a(.in(layer_2[433]), .out(far_3_3183_0[0]));    relay_conn far_3_3183_0_b(.in(layer_2[491]), .out(far_3_3183_0[1]));
    assign layer_3[123] = ~far_3_3183_0[1] | (far_3_3183_0[0] & far_3_3183_0[1]); 
    wire [1:0] far_3_3184_0;    relay_conn far_3_3184_0_a(.in(layer_2[50]), .out(far_3_3184_0[0]));    relay_conn far_3_3184_0_b(.in(layer_2[118]), .out(far_3_3184_0[1]));
    wire [1:0] far_3_3184_1;    relay_conn far_3_3184_1_a(.in(far_3_3184_0[0]), .out(far_3_3184_1[0]));    relay_conn far_3_3184_1_b(.in(far_3_3184_0[1]), .out(far_3_3184_1[1]));
    assign layer_3[124] = far_3_3184_1[1] & ~far_3_3184_1[0]; 
    wire [1:0] far_3_3185_0;    relay_conn far_3_3185_0_a(.in(layer_2[354]), .out(far_3_3185_0[0]));    relay_conn far_3_3185_0_b(.in(layer_2[304]), .out(far_3_3185_0[1]));
    assign layer_3[125] = ~far_3_3185_0[1]; 
    assign layer_3[126] = ~(layer_2[265] | layer_2[281]); 
    wire [1:0] far_3_3187_0;    relay_conn far_3_3187_0_a(.in(layer_2[378]), .out(far_3_3187_0[0]));    relay_conn far_3_3187_0_b(.in(layer_2[496]), .out(far_3_3187_0[1]));
    wire [1:0] far_3_3187_1;    relay_conn far_3_3187_1_a(.in(far_3_3187_0[0]), .out(far_3_3187_1[0]));    relay_conn far_3_3187_1_b(.in(far_3_3187_0[1]), .out(far_3_3187_1[1]));
    wire [1:0] far_3_3187_2;    relay_conn far_3_3187_2_a(.in(far_3_3187_1[0]), .out(far_3_3187_2[0]));    relay_conn far_3_3187_2_b(.in(far_3_3187_1[1]), .out(far_3_3187_2[1]));
    assign layer_3[127] = ~(far_3_3187_2[0] & far_3_3187_2[1]); 
    wire [1:0] far_3_3188_0;    relay_conn far_3_3188_0_a(.in(layer_2[701]), .out(far_3_3188_0[0]));    relay_conn far_3_3188_0_b(.in(layer_2[633]), .out(far_3_3188_0[1]));
    wire [1:0] far_3_3188_1;    relay_conn far_3_3188_1_a(.in(far_3_3188_0[0]), .out(far_3_3188_1[0]));    relay_conn far_3_3188_1_b(.in(far_3_3188_0[1]), .out(far_3_3188_1[1]));
    assign layer_3[128] = ~far_3_3188_1[0]; 
    wire [1:0] far_3_3189_0;    relay_conn far_3_3189_0_a(.in(layer_2[785]), .out(far_3_3189_0[0]));    relay_conn far_3_3189_0_b(.in(layer_2[741]), .out(far_3_3189_0[1]));
    assign layer_3[129] = far_3_3189_0[1]; 
    wire [1:0] far_3_3190_0;    relay_conn far_3_3190_0_a(.in(layer_2[208]), .out(far_3_3190_0[0]));    relay_conn far_3_3190_0_b(.in(layer_2[261]), .out(far_3_3190_0[1]));
    assign layer_3[130] = ~(far_3_3190_0[0] | far_3_3190_0[1]); 
    wire [1:0] far_3_3191_0;    relay_conn far_3_3191_0_a(.in(layer_2[471]), .out(far_3_3191_0[0]));    relay_conn far_3_3191_0_b(.in(layer_2[349]), .out(far_3_3191_0[1]));
    wire [1:0] far_3_3191_1;    relay_conn far_3_3191_1_a(.in(far_3_3191_0[0]), .out(far_3_3191_1[0]));    relay_conn far_3_3191_1_b(.in(far_3_3191_0[1]), .out(far_3_3191_1[1]));
    wire [1:0] far_3_3191_2;    relay_conn far_3_3191_2_a(.in(far_3_3191_1[0]), .out(far_3_3191_2[0]));    relay_conn far_3_3191_2_b(.in(far_3_3191_1[1]), .out(far_3_3191_2[1]));
    assign layer_3[131] = ~(far_3_3191_2[0] & far_3_3191_2[1]); 
    assign layer_3[132] = ~(layer_2[361] ^ layer_2[370]); 
    wire [1:0] far_3_3193_0;    relay_conn far_3_3193_0_a(.in(layer_2[487]), .out(far_3_3193_0[0]));    relay_conn far_3_3193_0_b(.in(layer_2[565]), .out(far_3_3193_0[1]));
    wire [1:0] far_3_3193_1;    relay_conn far_3_3193_1_a(.in(far_3_3193_0[0]), .out(far_3_3193_1[0]));    relay_conn far_3_3193_1_b(.in(far_3_3193_0[1]), .out(far_3_3193_1[1]));
    assign layer_3[133] = ~far_3_3193_1[0]; 
    assign layer_3[134] = ~(layer_2[304] & layer_2[324]); 
    wire [1:0] far_3_3195_0;    relay_conn far_3_3195_0_a(.in(layer_2[718]), .out(far_3_3195_0[0]));    relay_conn far_3_3195_0_b(.in(layer_2[843]), .out(far_3_3195_0[1]));
    wire [1:0] far_3_3195_1;    relay_conn far_3_3195_1_a(.in(far_3_3195_0[0]), .out(far_3_3195_1[0]));    relay_conn far_3_3195_1_b(.in(far_3_3195_0[1]), .out(far_3_3195_1[1]));
    wire [1:0] far_3_3195_2;    relay_conn far_3_3195_2_a(.in(far_3_3195_1[0]), .out(far_3_3195_2[0]));    relay_conn far_3_3195_2_b(.in(far_3_3195_1[1]), .out(far_3_3195_2[1]));
    assign layer_3[135] = far_3_3195_2[0]; 
    wire [1:0] far_3_3196_0;    relay_conn far_3_3196_0_a(.in(layer_2[815]), .out(far_3_3196_0[0]));    relay_conn far_3_3196_0_b(.in(layer_2[778]), .out(far_3_3196_0[1]));
    assign layer_3[136] = far_3_3196_0[1]; 
    wire [1:0] far_3_3197_0;    relay_conn far_3_3197_0_a(.in(layer_2[369]), .out(far_3_3197_0[0]));    relay_conn far_3_3197_0_b(.in(layer_2[471]), .out(far_3_3197_0[1]));
    wire [1:0] far_3_3197_1;    relay_conn far_3_3197_1_a(.in(far_3_3197_0[0]), .out(far_3_3197_1[0]));    relay_conn far_3_3197_1_b(.in(far_3_3197_0[1]), .out(far_3_3197_1[1]));
    wire [1:0] far_3_3197_2;    relay_conn far_3_3197_2_a(.in(far_3_3197_1[0]), .out(far_3_3197_2[0]));    relay_conn far_3_3197_2_b(.in(far_3_3197_1[1]), .out(far_3_3197_2[1]));
    assign layer_3[137] = far_3_3197_2[1]; 
    assign layer_3[138] = layer_2[548] ^ layer_2[536]; 
    wire [1:0] far_3_3199_0;    relay_conn far_3_3199_0_a(.in(layer_2[260]), .out(far_3_3199_0[0]));    relay_conn far_3_3199_0_b(.in(layer_2[303]), .out(far_3_3199_0[1]));
    assign layer_3[139] = ~(far_3_3199_0[0] ^ far_3_3199_0[1]); 
    wire [1:0] far_3_3200_0;    relay_conn far_3_3200_0_a(.in(layer_2[639]), .out(far_3_3200_0[0]));    relay_conn far_3_3200_0_b(.in(layer_2[521]), .out(far_3_3200_0[1]));
    wire [1:0] far_3_3200_1;    relay_conn far_3_3200_1_a(.in(far_3_3200_0[0]), .out(far_3_3200_1[0]));    relay_conn far_3_3200_1_b(.in(far_3_3200_0[1]), .out(far_3_3200_1[1]));
    wire [1:0] far_3_3200_2;    relay_conn far_3_3200_2_a(.in(far_3_3200_1[0]), .out(far_3_3200_2[0]));    relay_conn far_3_3200_2_b(.in(far_3_3200_1[1]), .out(far_3_3200_2[1]));
    assign layer_3[140] = ~far_3_3200_2[1] | (far_3_3200_2[0] & far_3_3200_2[1]); 
    wire [1:0] far_3_3201_0;    relay_conn far_3_3201_0_a(.in(layer_2[278]), .out(far_3_3201_0[0]));    relay_conn far_3_3201_0_b(.in(layer_2[222]), .out(far_3_3201_0[1]));
    assign layer_3[141] = far_3_3201_0[0]; 
    wire [1:0] far_3_3202_0;    relay_conn far_3_3202_0_a(.in(layer_2[424]), .out(far_3_3202_0[0]));    relay_conn far_3_3202_0_b(.in(layer_2[324]), .out(far_3_3202_0[1]));
    wire [1:0] far_3_3202_1;    relay_conn far_3_3202_1_a(.in(far_3_3202_0[0]), .out(far_3_3202_1[0]));    relay_conn far_3_3202_1_b(.in(far_3_3202_0[1]), .out(far_3_3202_1[1]));
    wire [1:0] far_3_3202_2;    relay_conn far_3_3202_2_a(.in(far_3_3202_1[0]), .out(far_3_3202_2[0]));    relay_conn far_3_3202_2_b(.in(far_3_3202_1[1]), .out(far_3_3202_2[1]));
    assign layer_3[142] = far_3_3202_2[0] & far_3_3202_2[1]; 
    assign layer_3[143] = ~(layer_2[177] & layer_2[181]); 
    wire [1:0] far_3_3204_0;    relay_conn far_3_3204_0_a(.in(layer_2[177]), .out(far_3_3204_0[0]));    relay_conn far_3_3204_0_b(.in(layer_2[300]), .out(far_3_3204_0[1]));
    wire [1:0] far_3_3204_1;    relay_conn far_3_3204_1_a(.in(far_3_3204_0[0]), .out(far_3_3204_1[0]));    relay_conn far_3_3204_1_b(.in(far_3_3204_0[1]), .out(far_3_3204_1[1]));
    wire [1:0] far_3_3204_2;    relay_conn far_3_3204_2_a(.in(far_3_3204_1[0]), .out(far_3_3204_2[0]));    relay_conn far_3_3204_2_b(.in(far_3_3204_1[1]), .out(far_3_3204_2[1]));
    assign layer_3[144] = far_3_3204_2[0] & ~far_3_3204_2[1]; 
    wire [1:0] far_3_3205_0;    relay_conn far_3_3205_0_a(.in(layer_2[920]), .out(far_3_3205_0[0]));    relay_conn far_3_3205_0_b(.in(layer_2[877]), .out(far_3_3205_0[1]));
    assign layer_3[145] = ~(far_3_3205_0[0] ^ far_3_3205_0[1]); 
    assign layer_3[146] = layer_2[345]; 
    assign layer_3[147] = ~layer_2[167] | (layer_2[151] & layer_2[167]); 
    assign layer_3[148] = ~layer_2[850] | (layer_2[849] & layer_2[850]); 
    wire [1:0] far_3_3209_0;    relay_conn far_3_3209_0_a(.in(layer_2[818]), .out(far_3_3209_0[0]));    relay_conn far_3_3209_0_b(.in(layer_2[925]), .out(far_3_3209_0[1]));
    wire [1:0] far_3_3209_1;    relay_conn far_3_3209_1_a(.in(far_3_3209_0[0]), .out(far_3_3209_1[0]));    relay_conn far_3_3209_1_b(.in(far_3_3209_0[1]), .out(far_3_3209_1[1]));
    wire [1:0] far_3_3209_2;    relay_conn far_3_3209_2_a(.in(far_3_3209_1[0]), .out(far_3_3209_2[0]));    relay_conn far_3_3209_2_b(.in(far_3_3209_1[1]), .out(far_3_3209_2[1]));
    assign layer_3[149] = far_3_3209_2[1]; 
    wire [1:0] far_3_3210_0;    relay_conn far_3_3210_0_a(.in(layer_2[757]), .out(far_3_3210_0[0]));    relay_conn far_3_3210_0_b(.in(layer_2[876]), .out(far_3_3210_0[1]));
    wire [1:0] far_3_3210_1;    relay_conn far_3_3210_1_a(.in(far_3_3210_0[0]), .out(far_3_3210_1[0]));    relay_conn far_3_3210_1_b(.in(far_3_3210_0[1]), .out(far_3_3210_1[1]));
    wire [1:0] far_3_3210_2;    relay_conn far_3_3210_2_a(.in(far_3_3210_1[0]), .out(far_3_3210_2[0]));    relay_conn far_3_3210_2_b(.in(far_3_3210_1[1]), .out(far_3_3210_2[1]));
    assign layer_3[150] = ~(far_3_3210_2[0] | far_3_3210_2[1]); 
    wire [1:0] far_3_3211_0;    relay_conn far_3_3211_0_a(.in(layer_2[810]), .out(far_3_3211_0[0]));    relay_conn far_3_3211_0_b(.in(layer_2[737]), .out(far_3_3211_0[1]));
    wire [1:0] far_3_3211_1;    relay_conn far_3_3211_1_a(.in(far_3_3211_0[0]), .out(far_3_3211_1[0]));    relay_conn far_3_3211_1_b(.in(far_3_3211_0[1]), .out(far_3_3211_1[1]));
    assign layer_3[151] = ~(far_3_3211_1[0] | far_3_3211_1[1]); 
    wire [1:0] far_3_3212_0;    relay_conn far_3_3212_0_a(.in(layer_2[823]), .out(far_3_3212_0[0]));    relay_conn far_3_3212_0_b(.in(layer_2[758]), .out(far_3_3212_0[1]));
    wire [1:0] far_3_3212_1;    relay_conn far_3_3212_1_a(.in(far_3_3212_0[0]), .out(far_3_3212_1[0]));    relay_conn far_3_3212_1_b(.in(far_3_3212_0[1]), .out(far_3_3212_1[1]));
    assign layer_3[152] = far_3_3212_1[0]; 
    assign layer_3[153] = ~(layer_2[361] | layer_2[354]); 
    wire [1:0] far_3_3214_0;    relay_conn far_3_3214_0_a(.in(layer_2[385]), .out(far_3_3214_0[0]));    relay_conn far_3_3214_0_b(.in(layer_2[502]), .out(far_3_3214_0[1]));
    wire [1:0] far_3_3214_1;    relay_conn far_3_3214_1_a(.in(far_3_3214_0[0]), .out(far_3_3214_1[0]));    relay_conn far_3_3214_1_b(.in(far_3_3214_0[1]), .out(far_3_3214_1[1]));
    wire [1:0] far_3_3214_2;    relay_conn far_3_3214_2_a(.in(far_3_3214_1[0]), .out(far_3_3214_2[0]));    relay_conn far_3_3214_2_b(.in(far_3_3214_1[1]), .out(far_3_3214_2[1]));
    assign layer_3[154] = ~(far_3_3214_2[0] & far_3_3214_2[1]); 
    wire [1:0] far_3_3215_0;    relay_conn far_3_3215_0_a(.in(layer_2[868]), .out(far_3_3215_0[0]));    relay_conn far_3_3215_0_b(.in(layer_2[935]), .out(far_3_3215_0[1]));
    wire [1:0] far_3_3215_1;    relay_conn far_3_3215_1_a(.in(far_3_3215_0[0]), .out(far_3_3215_1[0]));    relay_conn far_3_3215_1_b(.in(far_3_3215_0[1]), .out(far_3_3215_1[1]));
    assign layer_3[155] = ~far_3_3215_1[1]; 
    wire [1:0] far_3_3216_0;    relay_conn far_3_3216_0_a(.in(layer_2[674]), .out(far_3_3216_0[0]));    relay_conn far_3_3216_0_b(.in(layer_2[577]), .out(far_3_3216_0[1]));
    wire [1:0] far_3_3216_1;    relay_conn far_3_3216_1_a(.in(far_3_3216_0[0]), .out(far_3_3216_1[0]));    relay_conn far_3_3216_1_b(.in(far_3_3216_0[1]), .out(far_3_3216_1[1]));
    wire [1:0] far_3_3216_2;    relay_conn far_3_3216_2_a(.in(far_3_3216_1[0]), .out(far_3_3216_2[0]));    relay_conn far_3_3216_2_b(.in(far_3_3216_1[1]), .out(far_3_3216_2[1]));
    assign layer_3[156] = ~far_3_3216_2[1] | (far_3_3216_2[0] & far_3_3216_2[1]); 
    wire [1:0] far_3_3217_0;    relay_conn far_3_3217_0_a(.in(layer_2[1012]), .out(far_3_3217_0[0]));    relay_conn far_3_3217_0_b(.in(layer_2[903]), .out(far_3_3217_0[1]));
    wire [1:0] far_3_3217_1;    relay_conn far_3_3217_1_a(.in(far_3_3217_0[0]), .out(far_3_3217_1[0]));    relay_conn far_3_3217_1_b(.in(far_3_3217_0[1]), .out(far_3_3217_1[1]));
    wire [1:0] far_3_3217_2;    relay_conn far_3_3217_2_a(.in(far_3_3217_1[0]), .out(far_3_3217_2[0]));    relay_conn far_3_3217_2_b(.in(far_3_3217_1[1]), .out(far_3_3217_2[1]));
    assign layer_3[157] = far_3_3217_2[1] & ~far_3_3217_2[0]; 
    assign layer_3[158] = layer_2[327] & ~layer_2[342]; 
    wire [1:0] far_3_3219_0;    relay_conn far_3_3219_0_a(.in(layer_2[198]), .out(far_3_3219_0[0]));    relay_conn far_3_3219_0_b(.in(layer_2[85]), .out(far_3_3219_0[1]));
    wire [1:0] far_3_3219_1;    relay_conn far_3_3219_1_a(.in(far_3_3219_0[0]), .out(far_3_3219_1[0]));    relay_conn far_3_3219_1_b(.in(far_3_3219_0[1]), .out(far_3_3219_1[1]));
    wire [1:0] far_3_3219_2;    relay_conn far_3_3219_2_a(.in(far_3_3219_1[0]), .out(far_3_3219_2[0]));    relay_conn far_3_3219_2_b(.in(far_3_3219_1[1]), .out(far_3_3219_2[1]));
    assign layer_3[159] = ~far_3_3219_2[0] | (far_3_3219_2[0] & far_3_3219_2[1]); 
    wire [1:0] far_3_3220_0;    relay_conn far_3_3220_0_a(.in(layer_2[181]), .out(far_3_3220_0[0]));    relay_conn far_3_3220_0_b(.in(layer_2[97]), .out(far_3_3220_0[1]));
    wire [1:0] far_3_3220_1;    relay_conn far_3_3220_1_a(.in(far_3_3220_0[0]), .out(far_3_3220_1[0]));    relay_conn far_3_3220_1_b(.in(far_3_3220_0[1]), .out(far_3_3220_1[1]));
    assign layer_3[160] = far_3_3220_1[1]; 
    assign layer_3[161] = layer_2[29] & layer_2[34]; 
    wire [1:0] far_3_3222_0;    relay_conn far_3_3222_0_a(.in(layer_2[305]), .out(far_3_3222_0[0]));    relay_conn far_3_3222_0_b(.in(layer_2[202]), .out(far_3_3222_0[1]));
    wire [1:0] far_3_3222_1;    relay_conn far_3_3222_1_a(.in(far_3_3222_0[0]), .out(far_3_3222_1[0]));    relay_conn far_3_3222_1_b(.in(far_3_3222_0[1]), .out(far_3_3222_1[1]));
    wire [1:0] far_3_3222_2;    relay_conn far_3_3222_2_a(.in(far_3_3222_1[0]), .out(far_3_3222_2[0]));    relay_conn far_3_3222_2_b(.in(far_3_3222_1[1]), .out(far_3_3222_2[1]));
    assign layer_3[162] = far_3_3222_2[0] & ~far_3_3222_2[1]; 
    wire [1:0] far_3_3223_0;    relay_conn far_3_3223_0_a(.in(layer_2[815]), .out(far_3_3223_0[0]));    relay_conn far_3_3223_0_b(.in(layer_2[931]), .out(far_3_3223_0[1]));
    wire [1:0] far_3_3223_1;    relay_conn far_3_3223_1_a(.in(far_3_3223_0[0]), .out(far_3_3223_1[0]));    relay_conn far_3_3223_1_b(.in(far_3_3223_0[1]), .out(far_3_3223_1[1]));
    wire [1:0] far_3_3223_2;    relay_conn far_3_3223_2_a(.in(far_3_3223_1[0]), .out(far_3_3223_2[0]));    relay_conn far_3_3223_2_b(.in(far_3_3223_1[1]), .out(far_3_3223_2[1]));
    assign layer_3[163] = ~far_3_3223_2[0]; 
    wire [1:0] far_3_3224_0;    relay_conn far_3_3224_0_a(.in(layer_2[946]), .out(far_3_3224_0[0]));    relay_conn far_3_3224_0_b(.in(layer_2[985]), .out(far_3_3224_0[1]));
    assign layer_3[164] = ~far_3_3224_0[1] | (far_3_3224_0[0] & far_3_3224_0[1]); 
    wire [1:0] far_3_3225_0;    relay_conn far_3_3225_0_a(.in(layer_2[802]), .out(far_3_3225_0[0]));    relay_conn far_3_3225_0_b(.in(layer_2[849]), .out(far_3_3225_0[1]));
    assign layer_3[165] = far_3_3225_0[0] & far_3_3225_0[1]; 
    wire [1:0] far_3_3226_0;    relay_conn far_3_3226_0_a(.in(layer_2[920]), .out(far_3_3226_0[0]));    relay_conn far_3_3226_0_b(.in(layer_2[888]), .out(far_3_3226_0[1]));
    assign layer_3[166] = ~(far_3_3226_0[0] | far_3_3226_0[1]); 
    wire [1:0] far_3_3227_0;    relay_conn far_3_3227_0_a(.in(layer_2[71]), .out(far_3_3227_0[0]));    relay_conn far_3_3227_0_b(.in(layer_2[151]), .out(far_3_3227_0[1]));
    wire [1:0] far_3_3227_1;    relay_conn far_3_3227_1_a(.in(far_3_3227_0[0]), .out(far_3_3227_1[0]));    relay_conn far_3_3227_1_b(.in(far_3_3227_0[1]), .out(far_3_3227_1[1]));
    assign layer_3[167] = ~far_3_3227_1[0]; 
    wire [1:0] far_3_3228_0;    relay_conn far_3_3228_0_a(.in(layer_2[765]), .out(far_3_3228_0[0]));    relay_conn far_3_3228_0_b(.in(layer_2[877]), .out(far_3_3228_0[1]));
    wire [1:0] far_3_3228_1;    relay_conn far_3_3228_1_a(.in(far_3_3228_0[0]), .out(far_3_3228_1[0]));    relay_conn far_3_3228_1_b(.in(far_3_3228_0[1]), .out(far_3_3228_1[1]));
    wire [1:0] far_3_3228_2;    relay_conn far_3_3228_2_a(.in(far_3_3228_1[0]), .out(far_3_3228_2[0]));    relay_conn far_3_3228_2_b(.in(far_3_3228_1[1]), .out(far_3_3228_2[1]));
    assign layer_3[168] = far_3_3228_2[0]; 
    wire [1:0] far_3_3229_0;    relay_conn far_3_3229_0_a(.in(layer_2[913]), .out(far_3_3229_0[0]));    relay_conn far_3_3229_0_b(.in(layer_2[987]), .out(far_3_3229_0[1]));
    wire [1:0] far_3_3229_1;    relay_conn far_3_3229_1_a(.in(far_3_3229_0[0]), .out(far_3_3229_1[0]));    relay_conn far_3_3229_1_b(.in(far_3_3229_0[1]), .out(far_3_3229_1[1]));
    assign layer_3[169] = far_3_3229_1[1]; 
    wire [1:0] far_3_3230_0;    relay_conn far_3_3230_0_a(.in(layer_2[235]), .out(far_3_3230_0[0]));    relay_conn far_3_3230_0_b(.in(layer_2[300]), .out(far_3_3230_0[1]));
    wire [1:0] far_3_3230_1;    relay_conn far_3_3230_1_a(.in(far_3_3230_0[0]), .out(far_3_3230_1[0]));    relay_conn far_3_3230_1_b(.in(far_3_3230_0[1]), .out(far_3_3230_1[1]));
    assign layer_3[170] = far_3_3230_1[0]; 
    wire [1:0] far_3_3231_0;    relay_conn far_3_3231_0_a(.in(layer_2[267]), .out(far_3_3231_0[0]));    relay_conn far_3_3231_0_b(.in(layer_2[184]), .out(far_3_3231_0[1]));
    wire [1:0] far_3_3231_1;    relay_conn far_3_3231_1_a(.in(far_3_3231_0[0]), .out(far_3_3231_1[0]));    relay_conn far_3_3231_1_b(.in(far_3_3231_0[1]), .out(far_3_3231_1[1]));
    assign layer_3[171] = ~(far_3_3231_1[0] & far_3_3231_1[1]); 
    wire [1:0] far_3_3232_0;    relay_conn far_3_3232_0_a(.in(layer_2[891]), .out(far_3_3232_0[0]));    relay_conn far_3_3232_0_b(.in(layer_2[946]), .out(far_3_3232_0[1]));
    assign layer_3[172] = far_3_3232_0[0] | far_3_3232_0[1]; 
    wire [1:0] far_3_3233_0;    relay_conn far_3_3233_0_a(.in(layer_2[950]), .out(far_3_3233_0[0]));    relay_conn far_3_3233_0_b(.in(layer_2[897]), .out(far_3_3233_0[1]));
    assign layer_3[173] = ~far_3_3233_0[0] | (far_3_3233_0[0] & far_3_3233_0[1]); 
    wire [1:0] far_3_3234_0;    relay_conn far_3_3234_0_a(.in(layer_2[130]), .out(far_3_3234_0[0]));    relay_conn far_3_3234_0_b(.in(layer_2[213]), .out(far_3_3234_0[1]));
    wire [1:0] far_3_3234_1;    relay_conn far_3_3234_1_a(.in(far_3_3234_0[0]), .out(far_3_3234_1[0]));    relay_conn far_3_3234_1_b(.in(far_3_3234_0[1]), .out(far_3_3234_1[1]));
    assign layer_3[174] = far_3_3234_1[0] ^ far_3_3234_1[1]; 
    wire [1:0] far_3_3235_0;    relay_conn far_3_3235_0_a(.in(layer_2[345]), .out(far_3_3235_0[0]));    relay_conn far_3_3235_0_b(.in(layer_2[377]), .out(far_3_3235_0[1]));
    assign layer_3[175] = ~far_3_3235_0[0] | (far_3_3235_0[0] & far_3_3235_0[1]); 
    wire [1:0] far_3_3236_0;    relay_conn far_3_3236_0_a(.in(layer_2[710]), .out(far_3_3236_0[0]));    relay_conn far_3_3236_0_b(.in(layer_2[836]), .out(far_3_3236_0[1]));
    wire [1:0] far_3_3236_1;    relay_conn far_3_3236_1_a(.in(far_3_3236_0[0]), .out(far_3_3236_1[0]));    relay_conn far_3_3236_1_b(.in(far_3_3236_0[1]), .out(far_3_3236_1[1]));
    wire [1:0] far_3_3236_2;    relay_conn far_3_3236_2_a(.in(far_3_3236_1[0]), .out(far_3_3236_2[0]));    relay_conn far_3_3236_2_b(.in(far_3_3236_1[1]), .out(far_3_3236_2[1]));
    assign layer_3[176] = ~(far_3_3236_2[0] | far_3_3236_2[1]); 
    wire [1:0] far_3_3237_0;    relay_conn far_3_3237_0_a(.in(layer_2[988]), .out(far_3_3237_0[0]));    relay_conn far_3_3237_0_b(.in(layer_2[920]), .out(far_3_3237_0[1]));
    wire [1:0] far_3_3237_1;    relay_conn far_3_3237_1_a(.in(far_3_3237_0[0]), .out(far_3_3237_1[0]));    relay_conn far_3_3237_1_b(.in(far_3_3237_0[1]), .out(far_3_3237_1[1]));
    assign layer_3[177] = ~(far_3_3237_1[0] | far_3_3237_1[1]); 
    wire [1:0] far_3_3238_0;    relay_conn far_3_3238_0_a(.in(layer_2[151]), .out(far_3_3238_0[0]));    relay_conn far_3_3238_0_b(.in(layer_2[32]), .out(far_3_3238_0[1]));
    wire [1:0] far_3_3238_1;    relay_conn far_3_3238_1_a(.in(far_3_3238_0[0]), .out(far_3_3238_1[0]));    relay_conn far_3_3238_1_b(.in(far_3_3238_0[1]), .out(far_3_3238_1[1]));
    wire [1:0] far_3_3238_2;    relay_conn far_3_3238_2_a(.in(far_3_3238_1[0]), .out(far_3_3238_2[0]));    relay_conn far_3_3238_2_b(.in(far_3_3238_1[1]), .out(far_3_3238_2[1]));
    assign layer_3[178] = ~far_3_3238_2[0] | (far_3_3238_2[0] & far_3_3238_2[1]); 
    wire [1:0] far_3_3239_0;    relay_conn far_3_3239_0_a(.in(layer_2[218]), .out(far_3_3239_0[0]));    relay_conn far_3_3239_0_b(.in(layer_2[304]), .out(far_3_3239_0[1]));
    wire [1:0] far_3_3239_1;    relay_conn far_3_3239_1_a(.in(far_3_3239_0[0]), .out(far_3_3239_1[0]));    relay_conn far_3_3239_1_b(.in(far_3_3239_0[1]), .out(far_3_3239_1[1]));
    assign layer_3[179] = ~far_3_3239_1[0] | (far_3_3239_1[0] & far_3_3239_1[1]); 
    wire [1:0] far_3_3240_0;    relay_conn far_3_3240_0_a(.in(layer_2[198]), .out(far_3_3240_0[0]));    relay_conn far_3_3240_0_b(.in(layer_2[129]), .out(far_3_3240_0[1]));
    wire [1:0] far_3_3240_1;    relay_conn far_3_3240_1_a(.in(far_3_3240_0[0]), .out(far_3_3240_1[0]));    relay_conn far_3_3240_1_b(.in(far_3_3240_0[1]), .out(far_3_3240_1[1]));
    assign layer_3[180] = ~(far_3_3240_1[0] ^ far_3_3240_1[1]); 
    wire [1:0] far_3_3241_0;    relay_conn far_3_3241_0_a(.in(layer_2[852]), .out(far_3_3241_0[0]));    relay_conn far_3_3241_0_b(.in(layer_2[809]), .out(far_3_3241_0[1]));
    assign layer_3[181] = far_3_3241_0[0] ^ far_3_3241_0[1]; 
    assign layer_3[182] = layer_2[533] & layer_2[521]; 
    wire [1:0] far_3_3243_0;    relay_conn far_3_3243_0_a(.in(layer_2[154]), .out(far_3_3243_0[0]));    relay_conn far_3_3243_0_b(.in(layer_2[101]), .out(far_3_3243_0[1]));
    assign layer_3[183] = far_3_3243_0[0] ^ far_3_3243_0[1]; 
    wire [1:0] far_3_3244_0;    relay_conn far_3_3244_0_a(.in(layer_2[199]), .out(far_3_3244_0[0]));    relay_conn far_3_3244_0_b(.in(layer_2[323]), .out(far_3_3244_0[1]));
    wire [1:0] far_3_3244_1;    relay_conn far_3_3244_1_a(.in(far_3_3244_0[0]), .out(far_3_3244_1[0]));    relay_conn far_3_3244_1_b(.in(far_3_3244_0[1]), .out(far_3_3244_1[1]));
    wire [1:0] far_3_3244_2;    relay_conn far_3_3244_2_a(.in(far_3_3244_1[0]), .out(far_3_3244_2[0]));    relay_conn far_3_3244_2_b(.in(far_3_3244_1[1]), .out(far_3_3244_2[1]));
    assign layer_3[184] = ~(far_3_3244_2[0] & far_3_3244_2[1]); 
    wire [1:0] far_3_3245_0;    relay_conn far_3_3245_0_a(.in(layer_2[412]), .out(far_3_3245_0[0]));    relay_conn far_3_3245_0_b(.in(layer_2[348]), .out(far_3_3245_0[1]));
    wire [1:0] far_3_3245_1;    relay_conn far_3_3245_1_a(.in(far_3_3245_0[0]), .out(far_3_3245_1[0]));    relay_conn far_3_3245_1_b(.in(far_3_3245_0[1]), .out(far_3_3245_1[1]));
    assign layer_3[185] = ~(far_3_3245_1[0] | far_3_3245_1[1]); 
    assign layer_3[186] = layer_2[708] & ~layer_2[727]; 
    wire [1:0] far_3_3247_0;    relay_conn far_3_3247_0_a(.in(layer_2[258]), .out(far_3_3247_0[0]));    relay_conn far_3_3247_0_b(.in(layer_2[354]), .out(far_3_3247_0[1]));
    wire [1:0] far_3_3247_1;    relay_conn far_3_3247_1_a(.in(far_3_3247_0[0]), .out(far_3_3247_1[0]));    relay_conn far_3_3247_1_b(.in(far_3_3247_0[1]), .out(far_3_3247_1[1]));
    wire [1:0] far_3_3247_2;    relay_conn far_3_3247_2_a(.in(far_3_3247_1[0]), .out(far_3_3247_2[0]));    relay_conn far_3_3247_2_b(.in(far_3_3247_1[1]), .out(far_3_3247_2[1]));
    assign layer_3[187] = ~far_3_3247_2[0]; 
    wire [1:0] far_3_3248_0;    relay_conn far_3_3248_0_a(.in(layer_2[726]), .out(far_3_3248_0[0]));    relay_conn far_3_3248_0_b(.in(layer_2[670]), .out(far_3_3248_0[1]));
    assign layer_3[188] = far_3_3248_0[0] ^ far_3_3248_0[1]; 
    wire [1:0] far_3_3249_0;    relay_conn far_3_3249_0_a(.in(layer_2[12]), .out(far_3_3249_0[0]));    relay_conn far_3_3249_0_b(.in(layer_2[104]), .out(far_3_3249_0[1]));
    wire [1:0] far_3_3249_1;    relay_conn far_3_3249_1_a(.in(far_3_3249_0[0]), .out(far_3_3249_1[0]));    relay_conn far_3_3249_1_b(.in(far_3_3249_0[1]), .out(far_3_3249_1[1]));
    assign layer_3[189] = ~far_3_3249_1[1]; 
    wire [1:0] far_3_3250_0;    relay_conn far_3_3250_0_a(.in(layer_2[43]), .out(far_3_3250_0[0]));    relay_conn far_3_3250_0_b(.in(layer_2[151]), .out(far_3_3250_0[1]));
    wire [1:0] far_3_3250_1;    relay_conn far_3_3250_1_a(.in(far_3_3250_0[0]), .out(far_3_3250_1[0]));    relay_conn far_3_3250_1_b(.in(far_3_3250_0[1]), .out(far_3_3250_1[1]));
    wire [1:0] far_3_3250_2;    relay_conn far_3_3250_2_a(.in(far_3_3250_1[0]), .out(far_3_3250_2[0]));    relay_conn far_3_3250_2_b(.in(far_3_3250_1[1]), .out(far_3_3250_2[1]));
    assign layer_3[190] = ~(far_3_3250_2[0] & far_3_3250_2[1]); 
    wire [1:0] far_3_3251_0;    relay_conn far_3_3251_0_a(.in(layer_2[208]), .out(far_3_3251_0[0]));    relay_conn far_3_3251_0_b(.in(layer_2[130]), .out(far_3_3251_0[1]));
    wire [1:0] far_3_3251_1;    relay_conn far_3_3251_1_a(.in(far_3_3251_0[0]), .out(far_3_3251_1[0]));    relay_conn far_3_3251_1_b(.in(far_3_3251_0[1]), .out(far_3_3251_1[1]));
    assign layer_3[191] = far_3_3251_1[0] & far_3_3251_1[1]; 
    assign layer_3[192] = layer_2[768] & ~layer_2[748]; 
    assign layer_3[193] = ~(layer_2[22] | layer_2[50]); 
    wire [1:0] far_3_3254_0;    relay_conn far_3_3254_0_a(.in(layer_2[101]), .out(far_3_3254_0[0]));    relay_conn far_3_3254_0_b(.in(layer_2[6]), .out(far_3_3254_0[1]));
    wire [1:0] far_3_3254_1;    relay_conn far_3_3254_1_a(.in(far_3_3254_0[0]), .out(far_3_3254_1[0]));    relay_conn far_3_3254_1_b(.in(far_3_3254_0[1]), .out(far_3_3254_1[1]));
    assign layer_3[194] = far_3_3254_1[0] & far_3_3254_1[1]; 
    wire [1:0] far_3_3255_0;    relay_conn far_3_3255_0_a(.in(layer_2[416]), .out(far_3_3255_0[0]));    relay_conn far_3_3255_0_b(.in(layer_2[508]), .out(far_3_3255_0[1]));
    wire [1:0] far_3_3255_1;    relay_conn far_3_3255_1_a(.in(far_3_3255_0[0]), .out(far_3_3255_1[0]));    relay_conn far_3_3255_1_b(.in(far_3_3255_0[1]), .out(far_3_3255_1[1]));
    assign layer_3[195] = far_3_3255_1[0]; 
    assign layer_3[196] = layer_2[785] & ~layer_2[757]; 
    wire [1:0] far_3_3257_0;    relay_conn far_3_3257_0_a(.in(layer_2[664]), .out(far_3_3257_0[0]));    relay_conn far_3_3257_0_b(.in(layer_2[604]), .out(far_3_3257_0[1]));
    assign layer_3[197] = ~far_3_3257_0[0]; 
    wire [1:0] far_3_3258_0;    relay_conn far_3_3258_0_a(.in(layer_2[146]), .out(far_3_3258_0[0]));    relay_conn far_3_3258_0_b(.in(layer_2[181]), .out(far_3_3258_0[1]));
    assign layer_3[198] = far_3_3258_0[0] & ~far_3_3258_0[1]; 
    wire [1:0] far_3_3259_0;    relay_conn far_3_3259_0_a(.in(layer_2[354]), .out(far_3_3259_0[0]));    relay_conn far_3_3259_0_b(.in(layer_2[463]), .out(far_3_3259_0[1]));
    wire [1:0] far_3_3259_1;    relay_conn far_3_3259_1_a(.in(far_3_3259_0[0]), .out(far_3_3259_1[0]));    relay_conn far_3_3259_1_b(.in(far_3_3259_0[1]), .out(far_3_3259_1[1]));
    wire [1:0] far_3_3259_2;    relay_conn far_3_3259_2_a(.in(far_3_3259_1[0]), .out(far_3_3259_2[0]));    relay_conn far_3_3259_2_b(.in(far_3_3259_1[1]), .out(far_3_3259_2[1]));
    assign layer_3[199] = ~far_3_3259_2[1] | (far_3_3259_2[0] & far_3_3259_2[1]); 
    wire [1:0] far_3_3260_0;    relay_conn far_3_3260_0_a(.in(layer_2[221]), .out(far_3_3260_0[0]));    relay_conn far_3_3260_0_b(.in(layer_2[107]), .out(far_3_3260_0[1]));
    wire [1:0] far_3_3260_1;    relay_conn far_3_3260_1_a(.in(far_3_3260_0[0]), .out(far_3_3260_1[0]));    relay_conn far_3_3260_1_b(.in(far_3_3260_0[1]), .out(far_3_3260_1[1]));
    wire [1:0] far_3_3260_2;    relay_conn far_3_3260_2_a(.in(far_3_3260_1[0]), .out(far_3_3260_2[0]));    relay_conn far_3_3260_2_b(.in(far_3_3260_1[1]), .out(far_3_3260_2[1]));
    assign layer_3[200] = ~far_3_3260_2[1]; 
    wire [1:0] far_3_3261_0;    relay_conn far_3_3261_0_a(.in(layer_2[709]), .out(far_3_3261_0[0]));    relay_conn far_3_3261_0_b(.in(layer_2[769]), .out(far_3_3261_0[1]));
    assign layer_3[201] = far_3_3261_0[1]; 
    assign layer_3[202] = ~(layer_2[758] & layer_2[745]); 
    wire [1:0] far_3_3263_0;    relay_conn far_3_3263_0_a(.in(layer_2[75]), .out(far_3_3263_0[0]));    relay_conn far_3_3263_0_b(.in(layer_2[181]), .out(far_3_3263_0[1]));
    wire [1:0] far_3_3263_1;    relay_conn far_3_3263_1_a(.in(far_3_3263_0[0]), .out(far_3_3263_1[0]));    relay_conn far_3_3263_1_b(.in(far_3_3263_0[1]), .out(far_3_3263_1[1]));
    wire [1:0] far_3_3263_2;    relay_conn far_3_3263_2_a(.in(far_3_3263_1[0]), .out(far_3_3263_2[0]));    relay_conn far_3_3263_2_b(.in(far_3_3263_1[1]), .out(far_3_3263_2[1]));
    assign layer_3[203] = far_3_3263_2[0] & ~far_3_3263_2[1]; 
    assign layer_3[204] = ~layer_2[1005]; 
    wire [1:0] far_3_3265_0;    relay_conn far_3_3265_0_a(.in(layer_2[366]), .out(far_3_3265_0[0]));    relay_conn far_3_3265_0_b(.in(layer_2[489]), .out(far_3_3265_0[1]));
    wire [1:0] far_3_3265_1;    relay_conn far_3_3265_1_a(.in(far_3_3265_0[0]), .out(far_3_3265_1[0]));    relay_conn far_3_3265_1_b(.in(far_3_3265_0[1]), .out(far_3_3265_1[1]));
    wire [1:0] far_3_3265_2;    relay_conn far_3_3265_2_a(.in(far_3_3265_1[0]), .out(far_3_3265_2[0]));    relay_conn far_3_3265_2_b(.in(far_3_3265_1[1]), .out(far_3_3265_2[1]));
    assign layer_3[205] = far_3_3265_2[0] & far_3_3265_2[1]; 
    wire [1:0] far_3_3266_0;    relay_conn far_3_3266_0_a(.in(layer_2[412]), .out(far_3_3266_0[0]));    relay_conn far_3_3266_0_b(.in(layer_2[496]), .out(far_3_3266_0[1]));
    wire [1:0] far_3_3266_1;    relay_conn far_3_3266_1_a(.in(far_3_3266_0[0]), .out(far_3_3266_1[0]));    relay_conn far_3_3266_1_b(.in(far_3_3266_0[1]), .out(far_3_3266_1[1]));
    assign layer_3[206] = ~(far_3_3266_1[0] | far_3_3266_1[1]); 
    wire [1:0] far_3_3267_0;    relay_conn far_3_3267_0_a(.in(layer_2[999]), .out(far_3_3267_0[0]));    relay_conn far_3_3267_0_b(.in(layer_2[949]), .out(far_3_3267_0[1]));
    assign layer_3[207] = ~far_3_3267_0[1] | (far_3_3267_0[0] & far_3_3267_0[1]); 
    assign layer_3[208] = layer_2[500]; 
    wire [1:0] far_3_3269_0;    relay_conn far_3_3269_0_a(.in(layer_2[927]), .out(far_3_3269_0[0]));    relay_conn far_3_3269_0_b(.in(layer_2[1012]), .out(far_3_3269_0[1]));
    wire [1:0] far_3_3269_1;    relay_conn far_3_3269_1_a(.in(far_3_3269_0[0]), .out(far_3_3269_1[0]));    relay_conn far_3_3269_1_b(.in(far_3_3269_0[1]), .out(far_3_3269_1[1]));
    assign layer_3[209] = far_3_3269_1[0] ^ far_3_3269_1[1]; 
    wire [1:0] far_3_3270_0;    relay_conn far_3_3270_0_a(.in(layer_2[791]), .out(far_3_3270_0[0]));    relay_conn far_3_3270_0_b(.in(layer_2[748]), .out(far_3_3270_0[1]));
    assign layer_3[210] = far_3_3270_0[1]; 
    wire [1:0] far_3_3271_0;    relay_conn far_3_3271_0_a(.in(layer_2[350]), .out(far_3_3271_0[0]));    relay_conn far_3_3271_0_b(.in(layer_2[250]), .out(far_3_3271_0[1]));
    wire [1:0] far_3_3271_1;    relay_conn far_3_3271_1_a(.in(far_3_3271_0[0]), .out(far_3_3271_1[0]));    relay_conn far_3_3271_1_b(.in(far_3_3271_0[1]), .out(far_3_3271_1[1]));
    wire [1:0] far_3_3271_2;    relay_conn far_3_3271_2_a(.in(far_3_3271_1[0]), .out(far_3_3271_2[0]));    relay_conn far_3_3271_2_b(.in(far_3_3271_1[1]), .out(far_3_3271_2[1]));
    assign layer_3[211] = far_3_3271_2[0]; 
    assign layer_3[212] = layer_2[835] & ~layer_2[852]; 
    assign layer_3[213] = ~(layer_2[662] ^ layer_2[649]); 
    wire [1:0] far_3_3274_0;    relay_conn far_3_3274_0_a(.in(layer_2[330]), .out(far_3_3274_0[0]));    relay_conn far_3_3274_0_b(.in(layer_2[207]), .out(far_3_3274_0[1]));
    wire [1:0] far_3_3274_1;    relay_conn far_3_3274_1_a(.in(far_3_3274_0[0]), .out(far_3_3274_1[0]));    relay_conn far_3_3274_1_b(.in(far_3_3274_0[1]), .out(far_3_3274_1[1]));
    wire [1:0] far_3_3274_2;    relay_conn far_3_3274_2_a(.in(far_3_3274_1[0]), .out(far_3_3274_2[0]));    relay_conn far_3_3274_2_b(.in(far_3_3274_1[1]), .out(far_3_3274_2[1]));
    assign layer_3[214] = far_3_3274_2[0]; 
    wire [1:0] far_3_3275_0;    relay_conn far_3_3275_0_a(.in(layer_2[986]), .out(far_3_3275_0[0]));    relay_conn far_3_3275_0_b(.in(layer_2[903]), .out(far_3_3275_0[1]));
    wire [1:0] far_3_3275_1;    relay_conn far_3_3275_1_a(.in(far_3_3275_0[0]), .out(far_3_3275_1[0]));    relay_conn far_3_3275_1_b(.in(far_3_3275_0[1]), .out(far_3_3275_1[1]));
    assign layer_3[215] = far_3_3275_1[0] & ~far_3_3275_1[1]; 
    wire [1:0] far_3_3276_0;    relay_conn far_3_3276_0_a(.in(layer_2[136]), .out(far_3_3276_0[0]));    relay_conn far_3_3276_0_b(.in(layer_2[27]), .out(far_3_3276_0[1]));
    wire [1:0] far_3_3276_1;    relay_conn far_3_3276_1_a(.in(far_3_3276_0[0]), .out(far_3_3276_1[0]));    relay_conn far_3_3276_1_b(.in(far_3_3276_0[1]), .out(far_3_3276_1[1]));
    wire [1:0] far_3_3276_2;    relay_conn far_3_3276_2_a(.in(far_3_3276_1[0]), .out(far_3_3276_2[0]));    relay_conn far_3_3276_2_b(.in(far_3_3276_1[1]), .out(far_3_3276_2[1]));
    assign layer_3[216] = ~(far_3_3276_2[0] ^ far_3_3276_2[1]); 
    wire [1:0] far_3_3277_0;    relay_conn far_3_3277_0_a(.in(layer_2[1008]), .out(far_3_3277_0[0]));    relay_conn far_3_3277_0_b(.in(layer_2[926]), .out(far_3_3277_0[1]));
    wire [1:0] far_3_3277_1;    relay_conn far_3_3277_1_a(.in(far_3_3277_0[0]), .out(far_3_3277_1[0]));    relay_conn far_3_3277_1_b(.in(far_3_3277_0[1]), .out(far_3_3277_1[1]));
    assign layer_3[217] = ~(far_3_3277_1[0] | far_3_3277_1[1]); 
    wire [1:0] far_3_3278_0;    relay_conn far_3_3278_0_a(.in(layer_2[841]), .out(far_3_3278_0[0]));    relay_conn far_3_3278_0_b(.in(layer_2[891]), .out(far_3_3278_0[1]));
    assign layer_3[218] = far_3_3278_0[0]; 
    assign layer_3[219] = ~(layer_2[336] ^ layer_2[341]); 
    wire [1:0] far_3_3280_0;    relay_conn far_3_3280_0_a(.in(layer_2[949]), .out(far_3_3280_0[0]));    relay_conn far_3_3280_0_b(.in(layer_2[891]), .out(far_3_3280_0[1]));
    assign layer_3[220] = ~far_3_3280_0[0] | (far_3_3280_0[0] & far_3_3280_0[1]); 
    wire [1:0] far_3_3281_0;    relay_conn far_3_3281_0_a(.in(layer_2[3]), .out(far_3_3281_0[0]));    relay_conn far_3_3281_0_b(.in(layer_2[65]), .out(far_3_3281_0[1]));
    assign layer_3[221] = ~far_3_3281_0[1]; 
    assign layer_3[222] = layer_2[65] | layer_2[82]; 
    wire [1:0] far_3_3283_0;    relay_conn far_3_3283_0_a(.in(layer_2[227]), .out(far_3_3283_0[0]));    relay_conn far_3_3283_0_b(.in(layer_2[334]), .out(far_3_3283_0[1]));
    wire [1:0] far_3_3283_1;    relay_conn far_3_3283_1_a(.in(far_3_3283_0[0]), .out(far_3_3283_1[0]));    relay_conn far_3_3283_1_b(.in(far_3_3283_0[1]), .out(far_3_3283_1[1]));
    wire [1:0] far_3_3283_2;    relay_conn far_3_3283_2_a(.in(far_3_3283_1[0]), .out(far_3_3283_2[0]));    relay_conn far_3_3283_2_b(.in(far_3_3283_1[1]), .out(far_3_3283_2[1]));
    assign layer_3[223] = ~(far_3_3283_2[0] ^ far_3_3283_2[1]); 
    wire [1:0] far_3_3284_0;    relay_conn far_3_3284_0_a(.in(layer_2[156]), .out(far_3_3284_0[0]));    relay_conn far_3_3284_0_b(.in(layer_2[271]), .out(far_3_3284_0[1]));
    wire [1:0] far_3_3284_1;    relay_conn far_3_3284_1_a(.in(far_3_3284_0[0]), .out(far_3_3284_1[0]));    relay_conn far_3_3284_1_b(.in(far_3_3284_0[1]), .out(far_3_3284_1[1]));
    wire [1:0] far_3_3284_2;    relay_conn far_3_3284_2_a(.in(far_3_3284_1[0]), .out(far_3_3284_2[0]));    relay_conn far_3_3284_2_b(.in(far_3_3284_1[1]), .out(far_3_3284_2[1]));
    assign layer_3[224] = ~(far_3_3284_2[0] ^ far_3_3284_2[1]); 
    wire [1:0] far_3_3285_0;    relay_conn far_3_3285_0_a(.in(layer_2[954]), .out(far_3_3285_0[0]));    relay_conn far_3_3285_0_b(.in(layer_2[1010]), .out(far_3_3285_0[1]));
    assign layer_3[225] = far_3_3285_0[0]; 
    assign layer_3[226] = layer_2[44] & ~layer_2[75]; 
    wire [1:0] far_3_3287_0;    relay_conn far_3_3287_0_a(.in(layer_2[24]), .out(far_3_3287_0[0]));    relay_conn far_3_3287_0_b(.in(layer_2[103]), .out(far_3_3287_0[1]));
    wire [1:0] far_3_3287_1;    relay_conn far_3_3287_1_a(.in(far_3_3287_0[0]), .out(far_3_3287_1[0]));    relay_conn far_3_3287_1_b(.in(far_3_3287_0[1]), .out(far_3_3287_1[1]));
    assign layer_3[227] = ~(far_3_3287_1[0] & far_3_3287_1[1]); 
    wire [1:0] far_3_3288_0;    relay_conn far_3_3288_0_a(.in(layer_2[534]), .out(far_3_3288_0[0]));    relay_conn far_3_3288_0_b(.in(layer_2[421]), .out(far_3_3288_0[1]));
    wire [1:0] far_3_3288_1;    relay_conn far_3_3288_1_a(.in(far_3_3288_0[0]), .out(far_3_3288_1[0]));    relay_conn far_3_3288_1_b(.in(far_3_3288_0[1]), .out(far_3_3288_1[1]));
    wire [1:0] far_3_3288_2;    relay_conn far_3_3288_2_a(.in(far_3_3288_1[0]), .out(far_3_3288_2[0]));    relay_conn far_3_3288_2_b(.in(far_3_3288_1[1]), .out(far_3_3288_2[1]));
    assign layer_3[228] = ~far_3_3288_2[1]; 
    wire [1:0] far_3_3289_0;    relay_conn far_3_3289_0_a(.in(layer_2[914]), .out(far_3_3289_0[0]));    relay_conn far_3_3289_0_b(.in(layer_2[878]), .out(far_3_3289_0[1]));
    assign layer_3[229] = ~far_3_3289_0[1]; 
    assign layer_3[230] = ~(layer_2[781] | layer_2[766]); 
    wire [1:0] far_3_3291_0;    relay_conn far_3_3291_0_a(.in(layer_2[811]), .out(far_3_3291_0[0]));    relay_conn far_3_3291_0_b(.in(layer_2[742]), .out(far_3_3291_0[1]));
    wire [1:0] far_3_3291_1;    relay_conn far_3_3291_1_a(.in(far_3_3291_0[0]), .out(far_3_3291_1[0]));    relay_conn far_3_3291_1_b(.in(far_3_3291_0[1]), .out(far_3_3291_1[1]));
    assign layer_3[231] = ~far_3_3291_1[1] | (far_3_3291_1[0] & far_3_3291_1[1]); 
    assign layer_3[232] = layer_2[233]; 
    wire [1:0] far_3_3293_0;    relay_conn far_3_3293_0_a(.in(layer_2[1004]), .out(far_3_3293_0[0]));    relay_conn far_3_3293_0_b(.in(layer_2[888]), .out(far_3_3293_0[1]));
    wire [1:0] far_3_3293_1;    relay_conn far_3_3293_1_a(.in(far_3_3293_0[0]), .out(far_3_3293_1[0]));    relay_conn far_3_3293_1_b(.in(far_3_3293_0[1]), .out(far_3_3293_1[1]));
    wire [1:0] far_3_3293_2;    relay_conn far_3_3293_2_a(.in(far_3_3293_1[0]), .out(far_3_3293_2[0]));    relay_conn far_3_3293_2_b(.in(far_3_3293_1[1]), .out(far_3_3293_2[1]));
    assign layer_3[233] = ~(far_3_3293_2[0] ^ far_3_3293_2[1]); 
    assign layer_3[234] = layer_2[606]; 
    wire [1:0] far_3_3295_0;    relay_conn far_3_3295_0_a(.in(layer_2[365]), .out(far_3_3295_0[0]));    relay_conn far_3_3295_0_b(.in(layer_2[471]), .out(far_3_3295_0[1]));
    wire [1:0] far_3_3295_1;    relay_conn far_3_3295_1_a(.in(far_3_3295_0[0]), .out(far_3_3295_1[0]));    relay_conn far_3_3295_1_b(.in(far_3_3295_0[1]), .out(far_3_3295_1[1]));
    wire [1:0] far_3_3295_2;    relay_conn far_3_3295_2_a(.in(far_3_3295_1[0]), .out(far_3_3295_2[0]));    relay_conn far_3_3295_2_b(.in(far_3_3295_1[1]), .out(far_3_3295_2[1]));
    assign layer_3[235] = far_3_3295_2[1] & ~far_3_3295_2[0]; 
    assign layer_3[236] = ~(layer_2[472] | layer_2[473]); 
    wire [1:0] far_3_3297_0;    relay_conn far_3_3297_0_a(.in(layer_2[306]), .out(far_3_3297_0[0]));    relay_conn far_3_3297_0_b(.in(layer_2[385]), .out(far_3_3297_0[1]));
    wire [1:0] far_3_3297_1;    relay_conn far_3_3297_1_a(.in(far_3_3297_0[0]), .out(far_3_3297_1[0]));    relay_conn far_3_3297_1_b(.in(far_3_3297_0[1]), .out(far_3_3297_1[1]));
    assign layer_3[237] = ~(far_3_3297_1[0] | far_3_3297_1[1]); 
    assign layer_3[238] = layer_2[547]; 
    wire [1:0] far_3_3299_0;    relay_conn far_3_3299_0_a(.in(layer_2[36]), .out(far_3_3299_0[0]));    relay_conn far_3_3299_0_b(.in(layer_2[87]), .out(far_3_3299_0[1]));
    assign layer_3[239] = far_3_3299_0[0] | far_3_3299_0[1]; 
    wire [1:0] far_3_3300_0;    relay_conn far_3_3300_0_a(.in(layer_2[785]), .out(far_3_3300_0[0]));    relay_conn far_3_3300_0_b(.in(layer_2[896]), .out(far_3_3300_0[1]));
    wire [1:0] far_3_3300_1;    relay_conn far_3_3300_1_a(.in(far_3_3300_0[0]), .out(far_3_3300_1[0]));    relay_conn far_3_3300_1_b(.in(far_3_3300_0[1]), .out(far_3_3300_1[1]));
    wire [1:0] far_3_3300_2;    relay_conn far_3_3300_2_a(.in(far_3_3300_1[0]), .out(far_3_3300_2[0]));    relay_conn far_3_3300_2_b(.in(far_3_3300_1[1]), .out(far_3_3300_2[1]));
    assign layer_3[240] = ~far_3_3300_2[0]; 
    wire [1:0] far_3_3301_0;    relay_conn far_3_3301_0_a(.in(layer_2[899]), .out(far_3_3301_0[0]));    relay_conn far_3_3301_0_b(.in(layer_2[953]), .out(far_3_3301_0[1]));
    assign layer_3[241] = far_3_3301_0[1]; 
    wire [1:0] far_3_3302_0;    relay_conn far_3_3302_0_a(.in(layer_2[433]), .out(far_3_3302_0[0]));    relay_conn far_3_3302_0_b(.in(layer_2[560]), .out(far_3_3302_0[1]));
    wire [1:0] far_3_3302_1;    relay_conn far_3_3302_1_a(.in(far_3_3302_0[0]), .out(far_3_3302_1[0]));    relay_conn far_3_3302_1_b(.in(far_3_3302_0[1]), .out(far_3_3302_1[1]));
    wire [1:0] far_3_3302_2;    relay_conn far_3_3302_2_a(.in(far_3_3302_1[0]), .out(far_3_3302_2[0]));    relay_conn far_3_3302_2_b(.in(far_3_3302_1[1]), .out(far_3_3302_2[1]));
    assign layer_3[242] = ~far_3_3302_2[1] | (far_3_3302_2[0] & far_3_3302_2[1]); 
    wire [1:0] far_3_3303_0;    relay_conn far_3_3303_0_a(.in(layer_2[140]), .out(far_3_3303_0[0]));    relay_conn far_3_3303_0_b(.in(layer_2[195]), .out(far_3_3303_0[1]));
    assign layer_3[243] = ~(far_3_3303_0[0] ^ far_3_3303_0[1]); 
    wire [1:0] far_3_3304_0;    relay_conn far_3_3304_0_a(.in(layer_2[681]), .out(far_3_3304_0[0]));    relay_conn far_3_3304_0_b(.in(layer_2[770]), .out(far_3_3304_0[1]));
    wire [1:0] far_3_3304_1;    relay_conn far_3_3304_1_a(.in(far_3_3304_0[0]), .out(far_3_3304_1[0]));    relay_conn far_3_3304_1_b(.in(far_3_3304_0[1]), .out(far_3_3304_1[1]));
    assign layer_3[244] = ~far_3_3304_1[0]; 
    assign layer_3[245] = ~(layer_2[362] | layer_2[341]); 
    assign layer_3[246] = layer_2[422]; 
    wire [1:0] far_3_3307_0;    relay_conn far_3_3307_0_a(.in(layer_2[674]), .out(far_3_3307_0[0]));    relay_conn far_3_3307_0_b(.in(layer_2[714]), .out(far_3_3307_0[1]));
    assign layer_3[247] = far_3_3307_0[0] & far_3_3307_0[1]; 
    wire [1:0] far_3_3308_0;    relay_conn far_3_3308_0_a(.in(layer_2[171]), .out(far_3_3308_0[0]));    relay_conn far_3_3308_0_b(.in(layer_2[211]), .out(far_3_3308_0[1]));
    assign layer_3[248] = far_3_3308_0[0] & ~far_3_3308_0[1]; 
    wire [1:0] far_3_3309_0;    relay_conn far_3_3309_0_a(.in(layer_2[32]), .out(far_3_3309_0[0]));    relay_conn far_3_3309_0_b(.in(layer_2[148]), .out(far_3_3309_0[1]));
    wire [1:0] far_3_3309_1;    relay_conn far_3_3309_1_a(.in(far_3_3309_0[0]), .out(far_3_3309_1[0]));    relay_conn far_3_3309_1_b(.in(far_3_3309_0[1]), .out(far_3_3309_1[1]));
    wire [1:0] far_3_3309_2;    relay_conn far_3_3309_2_a(.in(far_3_3309_1[0]), .out(far_3_3309_2[0]));    relay_conn far_3_3309_2_b(.in(far_3_3309_1[1]), .out(far_3_3309_2[1]));
    assign layer_3[249] = far_3_3309_2[0] & ~far_3_3309_2[1]; 
    wire [1:0] far_3_3310_0;    relay_conn far_3_3310_0_a(.in(layer_2[829]), .out(far_3_3310_0[0]));    relay_conn far_3_3310_0_b(.in(layer_2[726]), .out(far_3_3310_0[1]));
    wire [1:0] far_3_3310_1;    relay_conn far_3_3310_1_a(.in(far_3_3310_0[0]), .out(far_3_3310_1[0]));    relay_conn far_3_3310_1_b(.in(far_3_3310_0[1]), .out(far_3_3310_1[1]));
    wire [1:0] far_3_3310_2;    relay_conn far_3_3310_2_a(.in(far_3_3310_1[0]), .out(far_3_3310_2[0]));    relay_conn far_3_3310_2_b(.in(far_3_3310_1[1]), .out(far_3_3310_2[1]));
    assign layer_3[250] = ~far_3_3310_2[1] | (far_3_3310_2[0] & far_3_3310_2[1]); 
    assign layer_3[251] = layer_2[221] | layer_2[250]; 
    assign layer_3[252] = layer_2[859] & layer_2[842]; 
    assign layer_3[253] = layer_2[464] & layer_2[440]; 
    wire [1:0] far_3_3314_0;    relay_conn far_3_3314_0_a(.in(layer_2[663]), .out(far_3_3314_0[0]));    relay_conn far_3_3314_0_b(.in(layer_2[753]), .out(far_3_3314_0[1]));
    wire [1:0] far_3_3314_1;    relay_conn far_3_3314_1_a(.in(far_3_3314_0[0]), .out(far_3_3314_1[0]));    relay_conn far_3_3314_1_b(.in(far_3_3314_0[1]), .out(far_3_3314_1[1]));
    assign layer_3[254] = far_3_3314_1[0] ^ far_3_3314_1[1]; 
    wire [1:0] far_3_3315_0;    relay_conn far_3_3315_0_a(.in(layer_2[553]), .out(far_3_3315_0[0]));    relay_conn far_3_3315_0_b(.in(layer_2[590]), .out(far_3_3315_0[1]));
    assign layer_3[255] = far_3_3315_0[0] | far_3_3315_0[1]; 
    wire [1:0] far_3_3316_0;    relay_conn far_3_3316_0_a(.in(layer_2[500]), .out(far_3_3316_0[0]));    relay_conn far_3_3316_0_b(.in(layer_2[468]), .out(far_3_3316_0[1]));
    assign layer_3[256] = far_3_3316_0[1] & ~far_3_3316_0[0]; 
    assign layer_3[257] = layer_2[714] & ~layer_2[731]; 
    wire [1:0] far_3_3318_0;    relay_conn far_3_3318_0_a(.in(layer_2[51]), .out(far_3_3318_0[0]));    relay_conn far_3_3318_0_b(.in(layer_2[109]), .out(far_3_3318_0[1]));
    assign layer_3[258] = ~far_3_3318_0[0] | (far_3_3318_0[0] & far_3_3318_0[1]); 
    assign layer_3[259] = ~(layer_2[57] | layer_2[82]); 
    wire [1:0] far_3_3320_0;    relay_conn far_3_3320_0_a(.in(layer_2[487]), .out(far_3_3320_0[0]));    relay_conn far_3_3320_0_b(.in(layer_2[400]), .out(far_3_3320_0[1]));
    wire [1:0] far_3_3320_1;    relay_conn far_3_3320_1_a(.in(far_3_3320_0[0]), .out(far_3_3320_1[0]));    relay_conn far_3_3320_1_b(.in(far_3_3320_0[1]), .out(far_3_3320_1[1]));
    assign layer_3[260] = ~(far_3_3320_1[0] & far_3_3320_1[1]); 
    wire [1:0] far_3_3321_0;    relay_conn far_3_3321_0_a(.in(layer_2[824]), .out(far_3_3321_0[0]));    relay_conn far_3_3321_0_b(.in(layer_2[949]), .out(far_3_3321_0[1]));
    wire [1:0] far_3_3321_1;    relay_conn far_3_3321_1_a(.in(far_3_3321_0[0]), .out(far_3_3321_1[0]));    relay_conn far_3_3321_1_b(.in(far_3_3321_0[1]), .out(far_3_3321_1[1]));
    wire [1:0] far_3_3321_2;    relay_conn far_3_3321_2_a(.in(far_3_3321_1[0]), .out(far_3_3321_2[0]));    relay_conn far_3_3321_2_b(.in(far_3_3321_1[1]), .out(far_3_3321_2[1]));
    assign layer_3[261] = far_3_3321_2[0] & ~far_3_3321_2[1]; 
    wire [1:0] far_3_3322_0;    relay_conn far_3_3322_0_a(.in(layer_2[419]), .out(far_3_3322_0[0]));    relay_conn far_3_3322_0_b(.in(layer_2[301]), .out(far_3_3322_0[1]));
    wire [1:0] far_3_3322_1;    relay_conn far_3_3322_1_a(.in(far_3_3322_0[0]), .out(far_3_3322_1[0]));    relay_conn far_3_3322_1_b(.in(far_3_3322_0[1]), .out(far_3_3322_1[1]));
    wire [1:0] far_3_3322_2;    relay_conn far_3_3322_2_a(.in(far_3_3322_1[0]), .out(far_3_3322_2[0]));    relay_conn far_3_3322_2_b(.in(far_3_3322_1[1]), .out(far_3_3322_2[1]));
    assign layer_3[262] = far_3_3322_2[0] & ~far_3_3322_2[1]; 
    wire [1:0] far_3_3323_0;    relay_conn far_3_3323_0_a(.in(layer_2[227]), .out(far_3_3323_0[0]));    relay_conn far_3_3323_0_b(.in(layer_2[352]), .out(far_3_3323_0[1]));
    wire [1:0] far_3_3323_1;    relay_conn far_3_3323_1_a(.in(far_3_3323_0[0]), .out(far_3_3323_1[0]));    relay_conn far_3_3323_1_b(.in(far_3_3323_0[1]), .out(far_3_3323_1[1]));
    wire [1:0] far_3_3323_2;    relay_conn far_3_3323_2_a(.in(far_3_3323_1[0]), .out(far_3_3323_2[0]));    relay_conn far_3_3323_2_b(.in(far_3_3323_1[1]), .out(far_3_3323_2[1]));
    assign layer_3[263] = far_3_3323_2[1]; 
    wire [1:0] far_3_3324_0;    relay_conn far_3_3324_0_a(.in(layer_2[844]), .out(far_3_3324_0[0]));    relay_conn far_3_3324_0_b(.in(layer_2[797]), .out(far_3_3324_0[1]));
    assign layer_3[264] = ~far_3_3324_0[0]; 
    assign layer_3[265] = layer_2[126] & ~layer_2[151]; 
    wire [1:0] far_3_3326_0;    relay_conn far_3_3326_0_a(.in(layer_2[304]), .out(far_3_3326_0[0]));    relay_conn far_3_3326_0_b(.in(layer_2[201]), .out(far_3_3326_0[1]));
    wire [1:0] far_3_3326_1;    relay_conn far_3_3326_1_a(.in(far_3_3326_0[0]), .out(far_3_3326_1[0]));    relay_conn far_3_3326_1_b(.in(far_3_3326_0[1]), .out(far_3_3326_1[1]));
    wire [1:0] far_3_3326_2;    relay_conn far_3_3326_2_a(.in(far_3_3326_1[0]), .out(far_3_3326_2[0]));    relay_conn far_3_3326_2_b(.in(far_3_3326_1[1]), .out(far_3_3326_2[1]));
    assign layer_3[266] = far_3_3326_2[1]; 
    wire [1:0] far_3_3327_0;    relay_conn far_3_3327_0_a(.in(layer_2[191]), .out(far_3_3327_0[0]));    relay_conn far_3_3327_0_b(.in(layer_2[265]), .out(far_3_3327_0[1]));
    wire [1:0] far_3_3327_1;    relay_conn far_3_3327_1_a(.in(far_3_3327_0[0]), .out(far_3_3327_1[0]));    relay_conn far_3_3327_1_b(.in(far_3_3327_0[1]), .out(far_3_3327_1[1]));
    assign layer_3[267] = far_3_3327_1[0] & ~far_3_3327_1[1]; 
    wire [1:0] far_3_3328_0;    relay_conn far_3_3328_0_a(.in(layer_2[354]), .out(far_3_3328_0[0]));    relay_conn far_3_3328_0_b(.in(layer_2[264]), .out(far_3_3328_0[1]));
    wire [1:0] far_3_3328_1;    relay_conn far_3_3328_1_a(.in(far_3_3328_0[0]), .out(far_3_3328_1[0]));    relay_conn far_3_3328_1_b(.in(far_3_3328_0[1]), .out(far_3_3328_1[1]));
    assign layer_3[268] = ~far_3_3328_1[0]; 
    wire [1:0] far_3_3329_0;    relay_conn far_3_3329_0_a(.in(layer_2[368]), .out(far_3_3329_0[0]));    relay_conn far_3_3329_0_b(.in(layer_2[245]), .out(far_3_3329_0[1]));
    wire [1:0] far_3_3329_1;    relay_conn far_3_3329_1_a(.in(far_3_3329_0[0]), .out(far_3_3329_1[0]));    relay_conn far_3_3329_1_b(.in(far_3_3329_0[1]), .out(far_3_3329_1[1]));
    wire [1:0] far_3_3329_2;    relay_conn far_3_3329_2_a(.in(far_3_3329_1[0]), .out(far_3_3329_2[0]));    relay_conn far_3_3329_2_b(.in(far_3_3329_1[1]), .out(far_3_3329_2[1]));
    assign layer_3[269] = ~(far_3_3329_2[0] & far_3_3329_2[1]); 
    wire [1:0] far_3_3330_0;    relay_conn far_3_3330_0_a(.in(layer_2[779]), .out(far_3_3330_0[0]));    relay_conn far_3_3330_0_b(.in(layer_2[890]), .out(far_3_3330_0[1]));
    wire [1:0] far_3_3330_1;    relay_conn far_3_3330_1_a(.in(far_3_3330_0[0]), .out(far_3_3330_1[0]));    relay_conn far_3_3330_1_b(.in(far_3_3330_0[1]), .out(far_3_3330_1[1]));
    wire [1:0] far_3_3330_2;    relay_conn far_3_3330_2_a(.in(far_3_3330_1[0]), .out(far_3_3330_2[0]));    relay_conn far_3_3330_2_b(.in(far_3_3330_1[1]), .out(far_3_3330_2[1]));
    assign layer_3[270] = far_3_3330_2[0] & far_3_3330_2[1]; 
    assign layer_3[271] = ~layer_2[423] | (layer_2[404] & layer_2[423]); 
    wire [1:0] far_3_3332_0;    relay_conn far_3_3332_0_a(.in(layer_2[141]), .out(far_3_3332_0[0]));    relay_conn far_3_3332_0_b(.in(layer_2[235]), .out(far_3_3332_0[1]));
    wire [1:0] far_3_3332_1;    relay_conn far_3_3332_1_a(.in(far_3_3332_0[0]), .out(far_3_3332_1[0]));    relay_conn far_3_3332_1_b(.in(far_3_3332_0[1]), .out(far_3_3332_1[1]));
    assign layer_3[272] = far_3_3332_1[0]; 
    wire [1:0] far_3_3333_0;    relay_conn far_3_3333_0_a(.in(layer_2[956]), .out(far_3_3333_0[0]));    relay_conn far_3_3333_0_b(.in(layer_2[1002]), .out(far_3_3333_0[1]));
    assign layer_3[273] = far_3_3333_0[1]; 
    wire [1:0] far_3_3334_0;    relay_conn far_3_3334_0_a(.in(layer_2[496]), .out(far_3_3334_0[0]));    relay_conn far_3_3334_0_b(.in(layer_2[433]), .out(far_3_3334_0[1]));
    assign layer_3[274] = far_3_3334_0[0] & far_3_3334_0[1]; 
    wire [1:0] far_3_3335_0;    relay_conn far_3_3335_0_a(.in(layer_2[471]), .out(far_3_3335_0[0]));    relay_conn far_3_3335_0_b(.in(layer_2[415]), .out(far_3_3335_0[1]));
    assign layer_3[275] = far_3_3335_0[1] & ~far_3_3335_0[0]; 
    wire [1:0] far_3_3336_0;    relay_conn far_3_3336_0_a(.in(layer_2[651]), .out(far_3_3336_0[0]));    relay_conn far_3_3336_0_b(.in(layer_2[688]), .out(far_3_3336_0[1]));
    assign layer_3[276] = far_3_3336_0[1]; 
    assign layer_3[277] = layer_2[880] & ~layer_2[882]; 
    wire [1:0] far_3_3338_0;    relay_conn far_3_3338_0_a(.in(layer_2[67]), .out(far_3_3338_0[0]));    relay_conn far_3_3338_0_b(.in(layer_2[126]), .out(far_3_3338_0[1]));
    assign layer_3[278] = ~(far_3_3338_0[0] ^ far_3_3338_0[1]); 
    wire [1:0] far_3_3339_0;    relay_conn far_3_3339_0_a(.in(layer_2[682]), .out(far_3_3339_0[0]));    relay_conn far_3_3339_0_b(.in(layer_2[558]), .out(far_3_3339_0[1]));
    wire [1:0] far_3_3339_1;    relay_conn far_3_3339_1_a(.in(far_3_3339_0[0]), .out(far_3_3339_1[0]));    relay_conn far_3_3339_1_b(.in(far_3_3339_0[1]), .out(far_3_3339_1[1]));
    wire [1:0] far_3_3339_2;    relay_conn far_3_3339_2_a(.in(far_3_3339_1[0]), .out(far_3_3339_2[0]));    relay_conn far_3_3339_2_b(.in(far_3_3339_1[1]), .out(far_3_3339_2[1]));
    assign layer_3[279] = ~(far_3_3339_2[0] | far_3_3339_2[1]); 
    assign layer_3[280] = layer_2[281] | layer_2[295]; 
    wire [1:0] far_3_3341_0;    relay_conn far_3_3341_0_a(.in(layer_2[247]), .out(far_3_3341_0[0]));    relay_conn far_3_3341_0_b(.in(layer_2[126]), .out(far_3_3341_0[1]));
    wire [1:0] far_3_3341_1;    relay_conn far_3_3341_1_a(.in(far_3_3341_0[0]), .out(far_3_3341_1[0]));    relay_conn far_3_3341_1_b(.in(far_3_3341_0[1]), .out(far_3_3341_1[1]));
    wire [1:0] far_3_3341_2;    relay_conn far_3_3341_2_a(.in(far_3_3341_1[0]), .out(far_3_3341_2[0]));    relay_conn far_3_3341_2_b(.in(far_3_3341_1[1]), .out(far_3_3341_2[1]));
    assign layer_3[281] = ~(far_3_3341_2[0] & far_3_3341_2[1]); 
    wire [1:0] far_3_3342_0;    relay_conn far_3_3342_0_a(.in(layer_2[446]), .out(far_3_3342_0[0]));    relay_conn far_3_3342_0_b(.in(layer_2[509]), .out(far_3_3342_0[1]));
    assign layer_3[282] = far_3_3342_0[0] | far_3_3342_0[1]; 
    wire [1:0] far_3_3343_0;    relay_conn far_3_3343_0_a(.in(layer_2[130]), .out(far_3_3343_0[0]));    relay_conn far_3_3343_0_b(.in(layer_2[66]), .out(far_3_3343_0[1]));
    wire [1:0] far_3_3343_1;    relay_conn far_3_3343_1_a(.in(far_3_3343_0[0]), .out(far_3_3343_1[0]));    relay_conn far_3_3343_1_b(.in(far_3_3343_0[1]), .out(far_3_3343_1[1]));
    assign layer_3[283] = far_3_3343_1[0] & far_3_3343_1[1]; 
    wire [1:0] far_3_3344_0;    relay_conn far_3_3344_0_a(.in(layer_2[480]), .out(far_3_3344_0[0]));    relay_conn far_3_3344_0_b(.in(layer_2[386]), .out(far_3_3344_0[1]));
    wire [1:0] far_3_3344_1;    relay_conn far_3_3344_1_a(.in(far_3_3344_0[0]), .out(far_3_3344_1[0]));    relay_conn far_3_3344_1_b(.in(far_3_3344_0[1]), .out(far_3_3344_1[1]));
    assign layer_3[284] = ~far_3_3344_1[0] | (far_3_3344_1[0] & far_3_3344_1[1]); 
    wire [1:0] far_3_3345_0;    relay_conn far_3_3345_0_a(.in(layer_2[841]), .out(far_3_3345_0[0]));    relay_conn far_3_3345_0_b(.in(layer_2[727]), .out(far_3_3345_0[1]));
    wire [1:0] far_3_3345_1;    relay_conn far_3_3345_1_a(.in(far_3_3345_0[0]), .out(far_3_3345_1[0]));    relay_conn far_3_3345_1_b(.in(far_3_3345_0[1]), .out(far_3_3345_1[1]));
    wire [1:0] far_3_3345_2;    relay_conn far_3_3345_2_a(.in(far_3_3345_1[0]), .out(far_3_3345_2[0]));    relay_conn far_3_3345_2_b(.in(far_3_3345_1[1]), .out(far_3_3345_2[1]));
    assign layer_3[285] = far_3_3345_2[1] & ~far_3_3345_2[0]; 
    assign layer_3[286] = layer_2[483]; 
    wire [1:0] far_3_3347_0;    relay_conn far_3_3347_0_a(.in(layer_2[630]), .out(far_3_3347_0[0]));    relay_conn far_3_3347_0_b(.in(layer_2[509]), .out(far_3_3347_0[1]));
    wire [1:0] far_3_3347_1;    relay_conn far_3_3347_1_a(.in(far_3_3347_0[0]), .out(far_3_3347_1[0]));    relay_conn far_3_3347_1_b(.in(far_3_3347_0[1]), .out(far_3_3347_1[1]));
    wire [1:0] far_3_3347_2;    relay_conn far_3_3347_2_a(.in(far_3_3347_1[0]), .out(far_3_3347_2[0]));    relay_conn far_3_3347_2_b(.in(far_3_3347_1[1]), .out(far_3_3347_2[1]));
    assign layer_3[287] = ~far_3_3347_2[0] | (far_3_3347_2[0] & far_3_3347_2[1]); 
    wire [1:0] far_3_3348_0;    relay_conn far_3_3348_0_a(.in(layer_2[876]), .out(far_3_3348_0[0]));    relay_conn far_3_3348_0_b(.in(layer_2[797]), .out(far_3_3348_0[1]));
    wire [1:0] far_3_3348_1;    relay_conn far_3_3348_1_a(.in(far_3_3348_0[0]), .out(far_3_3348_1[0]));    relay_conn far_3_3348_1_b(.in(far_3_3348_0[1]), .out(far_3_3348_1[1]));
    assign layer_3[288] = far_3_3348_1[1] & ~far_3_3348_1[0]; 
    wire [1:0] far_3_3349_0;    relay_conn far_3_3349_0_a(.in(layer_2[590]), .out(far_3_3349_0[0]));    relay_conn far_3_3349_0_b(.in(layer_2[532]), .out(far_3_3349_0[1]));
    assign layer_3[289] = ~far_3_3349_0[1] | (far_3_3349_0[0] & far_3_3349_0[1]); 
    wire [1:0] far_3_3350_0;    relay_conn far_3_3350_0_a(.in(layer_2[777]), .out(far_3_3350_0[0]));    relay_conn far_3_3350_0_b(.in(layer_2[819]), .out(far_3_3350_0[1]));
    assign layer_3[290] = far_3_3350_0[0] & far_3_3350_0[1]; 
    wire [1:0] far_3_3351_0;    relay_conn far_3_3351_0_a(.in(layer_2[197]), .out(far_3_3351_0[0]));    relay_conn far_3_3351_0_b(.in(layer_2[233]), .out(far_3_3351_0[1]));
    assign layer_3[291] = far_3_3351_0[0]; 
    assign layer_3[292] = layer_2[992] ^ layer_2[989]; 
    wire [1:0] far_3_3353_0;    relay_conn far_3_3353_0_a(.in(layer_2[830]), .out(far_3_3353_0[0]));    relay_conn far_3_3353_0_b(.in(layer_2[757]), .out(far_3_3353_0[1]));
    wire [1:0] far_3_3353_1;    relay_conn far_3_3353_1_a(.in(far_3_3353_0[0]), .out(far_3_3353_1[0]));    relay_conn far_3_3353_1_b(.in(far_3_3353_0[1]), .out(far_3_3353_1[1]));
    assign layer_3[293] = far_3_3353_1[0] & far_3_3353_1[1]; 
    wire [1:0] far_3_3354_0;    relay_conn far_3_3354_0_a(.in(layer_2[85]), .out(far_3_3354_0[0]));    relay_conn far_3_3354_0_b(.in(layer_2[205]), .out(far_3_3354_0[1]));
    wire [1:0] far_3_3354_1;    relay_conn far_3_3354_1_a(.in(far_3_3354_0[0]), .out(far_3_3354_1[0]));    relay_conn far_3_3354_1_b(.in(far_3_3354_0[1]), .out(far_3_3354_1[1]));
    wire [1:0] far_3_3354_2;    relay_conn far_3_3354_2_a(.in(far_3_3354_1[0]), .out(far_3_3354_2[0]));    relay_conn far_3_3354_2_b(.in(far_3_3354_1[1]), .out(far_3_3354_2[1]));
    assign layer_3[294] = far_3_3354_2[0] | far_3_3354_2[1]; 
    wire [1:0] far_3_3355_0;    relay_conn far_3_3355_0_a(.in(layer_2[380]), .out(far_3_3355_0[0]));    relay_conn far_3_3355_0_b(.in(layer_2[463]), .out(far_3_3355_0[1]));
    wire [1:0] far_3_3355_1;    relay_conn far_3_3355_1_a(.in(far_3_3355_0[0]), .out(far_3_3355_1[0]));    relay_conn far_3_3355_1_b(.in(far_3_3355_0[1]), .out(far_3_3355_1[1]));
    assign layer_3[295] = ~(far_3_3355_1[0] & far_3_3355_1[1]); 
    wire [1:0] far_3_3356_0;    relay_conn far_3_3356_0_a(.in(layer_2[839]), .out(far_3_3356_0[0]));    relay_conn far_3_3356_0_b(.in(layer_2[949]), .out(far_3_3356_0[1]));
    wire [1:0] far_3_3356_1;    relay_conn far_3_3356_1_a(.in(far_3_3356_0[0]), .out(far_3_3356_1[0]));    relay_conn far_3_3356_1_b(.in(far_3_3356_0[1]), .out(far_3_3356_1[1]));
    wire [1:0] far_3_3356_2;    relay_conn far_3_3356_2_a(.in(far_3_3356_1[0]), .out(far_3_3356_2[0]));    relay_conn far_3_3356_2_b(.in(far_3_3356_1[1]), .out(far_3_3356_2[1]));
    assign layer_3[296] = far_3_3356_2[1] & ~far_3_3356_2[0]; 
    assign layer_3[297] = layer_2[572]; 
    assign layer_3[298] = layer_2[173] | layer_2[188]; 
    wire [1:0] far_3_3359_0;    relay_conn far_3_3359_0_a(.in(layer_2[254]), .out(far_3_3359_0[0]));    relay_conn far_3_3359_0_b(.in(layer_2[303]), .out(far_3_3359_0[1]));
    assign layer_3[299] = far_3_3359_0[0] & far_3_3359_0[1]; 
    wire [1:0] far_3_3360_0;    relay_conn far_3_3360_0_a(.in(layer_2[835]), .out(far_3_3360_0[0]));    relay_conn far_3_3360_0_b(.in(layer_2[920]), .out(far_3_3360_0[1]));
    wire [1:0] far_3_3360_1;    relay_conn far_3_3360_1_a(.in(far_3_3360_0[0]), .out(far_3_3360_1[0]));    relay_conn far_3_3360_1_b(.in(far_3_3360_0[1]), .out(far_3_3360_1[1]));
    assign layer_3[300] = far_3_3360_1[0] | far_3_3360_1[1]; 
    wire [1:0] far_3_3361_0;    relay_conn far_3_3361_0_a(.in(layer_2[950]), .out(far_3_3361_0[0]));    relay_conn far_3_3361_0_b(.in(layer_2[995]), .out(far_3_3361_0[1]));
    assign layer_3[301] = ~far_3_3361_0[1]; 
    wire [1:0] far_3_3362_0;    relay_conn far_3_3362_0_a(.in(layer_2[76]), .out(far_3_3362_0[0]));    relay_conn far_3_3362_0_b(.in(layer_2[110]), .out(far_3_3362_0[1]));
    assign layer_3[302] = ~far_3_3362_0[0]; 
    wire [1:0] far_3_3363_0;    relay_conn far_3_3363_0_a(.in(layer_2[146]), .out(far_3_3363_0[0]));    relay_conn far_3_3363_0_b(.in(layer_2[181]), .out(far_3_3363_0[1]));
    assign layer_3[303] = ~(far_3_3363_0[0] | far_3_3363_0[1]); 
    wire [1:0] far_3_3364_0;    relay_conn far_3_3364_0_a(.in(layer_2[899]), .out(far_3_3364_0[0]));    relay_conn far_3_3364_0_b(.in(layer_2[830]), .out(far_3_3364_0[1]));
    wire [1:0] far_3_3364_1;    relay_conn far_3_3364_1_a(.in(far_3_3364_0[0]), .out(far_3_3364_1[0]));    relay_conn far_3_3364_1_b(.in(far_3_3364_0[1]), .out(far_3_3364_1[1]));
    assign layer_3[304] = far_3_3364_1[1] & ~far_3_3364_1[0]; 
    wire [1:0] far_3_3365_0;    relay_conn far_3_3365_0_a(.in(layer_2[986]), .out(far_3_3365_0[0]));    relay_conn far_3_3365_0_b(.in(layer_2[859]), .out(far_3_3365_0[1]));
    wire [1:0] far_3_3365_1;    relay_conn far_3_3365_1_a(.in(far_3_3365_0[0]), .out(far_3_3365_1[0]));    relay_conn far_3_3365_1_b(.in(far_3_3365_0[1]), .out(far_3_3365_1[1]));
    wire [1:0] far_3_3365_2;    relay_conn far_3_3365_2_a(.in(far_3_3365_1[0]), .out(far_3_3365_2[0]));    relay_conn far_3_3365_2_b(.in(far_3_3365_1[1]), .out(far_3_3365_2[1]));
    assign layer_3[305] = ~far_3_3365_2[0]; 
    assign layer_3[306] = layer_2[845] & layer_2[839]; 
    wire [1:0] far_3_3367_0;    relay_conn far_3_3367_0_a(.in(layer_2[427]), .out(far_3_3367_0[0]));    relay_conn far_3_3367_0_b(.in(layer_2[345]), .out(far_3_3367_0[1]));
    wire [1:0] far_3_3367_1;    relay_conn far_3_3367_1_a(.in(far_3_3367_0[0]), .out(far_3_3367_1[0]));    relay_conn far_3_3367_1_b(.in(far_3_3367_0[1]), .out(far_3_3367_1[1]));
    assign layer_3[307] = far_3_3367_1[0] & far_3_3367_1[1]; 
    assign layer_3[308] = layer_2[733] & ~layer_2[742]; 
    wire [1:0] far_3_3369_0;    relay_conn far_3_3369_0_a(.in(layer_2[350]), .out(far_3_3369_0[0]));    relay_conn far_3_3369_0_b(.in(layer_2[307]), .out(far_3_3369_0[1]));
    assign layer_3[309] = far_3_3369_0[1] & ~far_3_3369_0[0]; 
    wire [1:0] far_3_3370_0;    relay_conn far_3_3370_0_a(.in(layer_2[835]), .out(far_3_3370_0[0]));    relay_conn far_3_3370_0_b(.in(layer_2[740]), .out(far_3_3370_0[1]));
    wire [1:0] far_3_3370_1;    relay_conn far_3_3370_1_a(.in(far_3_3370_0[0]), .out(far_3_3370_1[0]));    relay_conn far_3_3370_1_b(.in(far_3_3370_0[1]), .out(far_3_3370_1[1]));
    assign layer_3[310] = far_3_3370_1[0]; 
    wire [1:0] far_3_3371_0;    relay_conn far_3_3371_0_a(.in(layer_2[422]), .out(far_3_3371_0[0]));    relay_conn far_3_3371_0_b(.in(layer_2[376]), .out(far_3_3371_0[1]));
    assign layer_3[311] = ~(far_3_3371_0[0] ^ far_3_3371_0[1]); 
    assign layer_3[312] = layer_2[142]; 
    wire [1:0] far_3_3373_0;    relay_conn far_3_3373_0_a(.in(layer_2[379]), .out(far_3_3373_0[0]));    relay_conn far_3_3373_0_b(.in(layer_2[303]), .out(far_3_3373_0[1]));
    wire [1:0] far_3_3373_1;    relay_conn far_3_3373_1_a(.in(far_3_3373_0[0]), .out(far_3_3373_1[0]));    relay_conn far_3_3373_1_b(.in(far_3_3373_0[1]), .out(far_3_3373_1[1]));
    assign layer_3[313] = ~far_3_3373_1[1]; 
    wire [1:0] far_3_3374_0;    relay_conn far_3_3374_0_a(.in(layer_2[103]), .out(far_3_3374_0[0]));    relay_conn far_3_3374_0_b(.in(layer_2[151]), .out(far_3_3374_0[1]));
    assign layer_3[314] = far_3_3374_0[0]; 
    wire [1:0] far_3_3375_0;    relay_conn far_3_3375_0_a(.in(layer_2[626]), .out(far_3_3375_0[0]));    relay_conn far_3_3375_0_b(.in(layer_2[517]), .out(far_3_3375_0[1]));
    wire [1:0] far_3_3375_1;    relay_conn far_3_3375_1_a(.in(far_3_3375_0[0]), .out(far_3_3375_1[0]));    relay_conn far_3_3375_1_b(.in(far_3_3375_0[1]), .out(far_3_3375_1[1]));
    wire [1:0] far_3_3375_2;    relay_conn far_3_3375_2_a(.in(far_3_3375_1[0]), .out(far_3_3375_2[0]));    relay_conn far_3_3375_2_b(.in(far_3_3375_1[1]), .out(far_3_3375_2[1]));
    assign layer_3[315] = ~(far_3_3375_2[0] & far_3_3375_2[1]); 
    wire [1:0] far_3_3376_0;    relay_conn far_3_3376_0_a(.in(layer_2[156]), .out(far_3_3376_0[0]));    relay_conn far_3_3376_0_b(.in(layer_2[228]), .out(far_3_3376_0[1]));
    wire [1:0] far_3_3376_1;    relay_conn far_3_3376_1_a(.in(far_3_3376_0[0]), .out(far_3_3376_1[0]));    relay_conn far_3_3376_1_b(.in(far_3_3376_0[1]), .out(far_3_3376_1[1]));
    assign layer_3[316] = ~(far_3_3376_1[0] | far_3_3376_1[1]); 
    wire [1:0] far_3_3377_0;    relay_conn far_3_3377_0_a(.in(layer_2[201]), .out(far_3_3377_0[0]));    relay_conn far_3_3377_0_b(.in(layer_2[314]), .out(far_3_3377_0[1]));
    wire [1:0] far_3_3377_1;    relay_conn far_3_3377_1_a(.in(far_3_3377_0[0]), .out(far_3_3377_1[0]));    relay_conn far_3_3377_1_b(.in(far_3_3377_0[1]), .out(far_3_3377_1[1]));
    wire [1:0] far_3_3377_2;    relay_conn far_3_3377_2_a(.in(far_3_3377_1[0]), .out(far_3_3377_2[0]));    relay_conn far_3_3377_2_b(.in(far_3_3377_1[1]), .out(far_3_3377_2[1]));
    assign layer_3[317] = far_3_3377_2[0]; 
    wire [1:0] far_3_3378_0;    relay_conn far_3_3378_0_a(.in(layer_2[211]), .out(far_3_3378_0[0]));    relay_conn far_3_3378_0_b(.in(layer_2[325]), .out(far_3_3378_0[1]));
    wire [1:0] far_3_3378_1;    relay_conn far_3_3378_1_a(.in(far_3_3378_0[0]), .out(far_3_3378_1[0]));    relay_conn far_3_3378_1_b(.in(far_3_3378_0[1]), .out(far_3_3378_1[1]));
    wire [1:0] far_3_3378_2;    relay_conn far_3_3378_2_a(.in(far_3_3378_1[0]), .out(far_3_3378_2[0]));    relay_conn far_3_3378_2_b(.in(far_3_3378_1[1]), .out(far_3_3378_2[1]));
    assign layer_3[318] = ~far_3_3378_2[1]; 
    assign layer_3[319] = layer_2[65] | layer_2[67]; 
    wire [1:0] far_3_3380_0;    relay_conn far_3_3380_0_a(.in(layer_2[543]), .out(far_3_3380_0[0]));    relay_conn far_3_3380_0_b(.in(layer_2[505]), .out(far_3_3380_0[1]));
    assign layer_3[320] = ~far_3_3380_0[1] | (far_3_3380_0[0] & far_3_3380_0[1]); 
    wire [1:0] far_3_3381_0;    relay_conn far_3_3381_0_a(.in(layer_2[927]), .out(far_3_3381_0[0]));    relay_conn far_3_3381_0_b(.in(layer_2[992]), .out(far_3_3381_0[1]));
    wire [1:0] far_3_3381_1;    relay_conn far_3_3381_1_a(.in(far_3_3381_0[0]), .out(far_3_3381_1[0]));    relay_conn far_3_3381_1_b(.in(far_3_3381_0[1]), .out(far_3_3381_1[1]));
    assign layer_3[321] = ~far_3_3381_1[0]; 
    wire [1:0] far_3_3382_0;    relay_conn far_3_3382_0_a(.in(layer_2[755]), .out(far_3_3382_0[0]));    relay_conn far_3_3382_0_b(.in(layer_2[683]), .out(far_3_3382_0[1]));
    wire [1:0] far_3_3382_1;    relay_conn far_3_3382_1_a(.in(far_3_3382_0[0]), .out(far_3_3382_1[0]));    relay_conn far_3_3382_1_b(.in(far_3_3382_0[1]), .out(far_3_3382_1[1]));
    assign layer_3[322] = ~far_3_3382_1[1]; 
    assign layer_3[323] = ~layer_2[471] | (layer_2[471] & layer_2[445]); 
    wire [1:0] far_3_3384_0;    relay_conn far_3_3384_0_a(.in(layer_2[246]), .out(far_3_3384_0[0]));    relay_conn far_3_3384_0_b(.in(layer_2[326]), .out(far_3_3384_0[1]));
    wire [1:0] far_3_3384_1;    relay_conn far_3_3384_1_a(.in(far_3_3384_0[0]), .out(far_3_3384_1[0]));    relay_conn far_3_3384_1_b(.in(far_3_3384_0[1]), .out(far_3_3384_1[1]));
    assign layer_3[324] = far_3_3384_1[1] & ~far_3_3384_1[0]; 
    wire [1:0] far_3_3385_0;    relay_conn far_3_3385_0_a(.in(layer_2[194]), .out(far_3_3385_0[0]));    relay_conn far_3_3385_0_b(.in(layer_2[117]), .out(far_3_3385_0[1]));
    wire [1:0] far_3_3385_1;    relay_conn far_3_3385_1_a(.in(far_3_3385_0[0]), .out(far_3_3385_1[0]));    relay_conn far_3_3385_1_b(.in(far_3_3385_0[1]), .out(far_3_3385_1[1]));
    assign layer_3[325] = far_3_3385_1[0] | far_3_3385_1[1]; 
    wire [1:0] far_3_3386_0;    relay_conn far_3_3386_0_a(.in(layer_2[774]), .out(far_3_3386_0[0]));    relay_conn far_3_3386_0_b(.in(layer_2[812]), .out(far_3_3386_0[1]));
    assign layer_3[326] = far_3_3386_0[0]; 
    assign layer_3[327] = layer_2[50] & ~layer_2[43]; 
    assign layer_3[328] = ~layer_2[565]; 
    wire [1:0] far_3_3389_0;    relay_conn far_3_3389_0_a(.in(layer_2[998]), .out(far_3_3389_0[0]));    relay_conn far_3_3389_0_b(.in(layer_2[910]), .out(far_3_3389_0[1]));
    wire [1:0] far_3_3389_1;    relay_conn far_3_3389_1_a(.in(far_3_3389_0[0]), .out(far_3_3389_1[0]));    relay_conn far_3_3389_1_b(.in(far_3_3389_0[1]), .out(far_3_3389_1[1]));
    assign layer_3[329] = far_3_3389_1[0] & ~far_3_3389_1[1]; 
    wire [1:0] far_3_3390_0;    relay_conn far_3_3390_0_a(.in(layer_2[785]), .out(far_3_3390_0[0]));    relay_conn far_3_3390_0_b(.in(layer_2[910]), .out(far_3_3390_0[1]));
    wire [1:0] far_3_3390_1;    relay_conn far_3_3390_1_a(.in(far_3_3390_0[0]), .out(far_3_3390_1[0]));    relay_conn far_3_3390_1_b(.in(far_3_3390_0[1]), .out(far_3_3390_1[1]));
    wire [1:0] far_3_3390_2;    relay_conn far_3_3390_2_a(.in(far_3_3390_1[0]), .out(far_3_3390_2[0]));    relay_conn far_3_3390_2_b(.in(far_3_3390_1[1]), .out(far_3_3390_2[1]));
    assign layer_3[330] = far_3_3390_2[0] ^ far_3_3390_2[1]; 
    assign layer_3[331] = ~(layer_2[922] | layer_2[920]); 
    wire [1:0] far_3_3392_0;    relay_conn far_3_3392_0_a(.in(layer_2[327]), .out(far_3_3392_0[0]));    relay_conn far_3_3392_0_b(.in(layer_2[237]), .out(far_3_3392_0[1]));
    wire [1:0] far_3_3392_1;    relay_conn far_3_3392_1_a(.in(far_3_3392_0[0]), .out(far_3_3392_1[0]));    relay_conn far_3_3392_1_b(.in(far_3_3392_0[1]), .out(far_3_3392_1[1]));
    assign layer_3[332] = ~(far_3_3392_1[0] | far_3_3392_1[1]); 
    wire [1:0] far_3_3393_0;    relay_conn far_3_3393_0_a(.in(layer_2[636]), .out(far_3_3393_0[0]));    relay_conn far_3_3393_0_b(.in(layer_2[570]), .out(far_3_3393_0[1]));
    wire [1:0] far_3_3393_1;    relay_conn far_3_3393_1_a(.in(far_3_3393_0[0]), .out(far_3_3393_1[0]));    relay_conn far_3_3393_1_b(.in(far_3_3393_0[1]), .out(far_3_3393_1[1]));
    assign layer_3[333] = far_3_3393_1[0] & ~far_3_3393_1[1]; 
    assign layer_3[334] = ~layer_2[181]; 
    wire [1:0] far_3_3395_0;    relay_conn far_3_3395_0_a(.in(layer_2[900]), .out(far_3_3395_0[0]));    relay_conn far_3_3395_0_b(.in(layer_2[775]), .out(far_3_3395_0[1]));
    wire [1:0] far_3_3395_1;    relay_conn far_3_3395_1_a(.in(far_3_3395_0[0]), .out(far_3_3395_1[0]));    relay_conn far_3_3395_1_b(.in(far_3_3395_0[1]), .out(far_3_3395_1[1]));
    wire [1:0] far_3_3395_2;    relay_conn far_3_3395_2_a(.in(far_3_3395_1[0]), .out(far_3_3395_2[0]));    relay_conn far_3_3395_2_b(.in(far_3_3395_1[1]), .out(far_3_3395_2[1]));
    assign layer_3[335] = ~far_3_3395_2[0] | (far_3_3395_2[0] & far_3_3395_2[1]); 
    wire [1:0] far_3_3396_0;    relay_conn far_3_3396_0_a(.in(layer_2[151]), .out(far_3_3396_0[0]));    relay_conn far_3_3396_0_b(.in(layer_2[188]), .out(far_3_3396_0[1]));
    assign layer_3[336] = ~far_3_3396_0[1] | (far_3_3396_0[0] & far_3_3396_0[1]); 
    wire [1:0] far_3_3397_0;    relay_conn far_3_3397_0_a(.in(layer_2[188]), .out(far_3_3397_0[0]));    relay_conn far_3_3397_0_b(.in(layer_2[94]), .out(far_3_3397_0[1]));
    wire [1:0] far_3_3397_1;    relay_conn far_3_3397_1_a(.in(far_3_3397_0[0]), .out(far_3_3397_1[0]));    relay_conn far_3_3397_1_b(.in(far_3_3397_0[1]), .out(far_3_3397_1[1]));
    assign layer_3[337] = far_3_3397_1[1] & ~far_3_3397_1[0]; 
    wire [1:0] far_3_3398_0;    relay_conn far_3_3398_0_a(.in(layer_2[265]), .out(far_3_3398_0[0]));    relay_conn far_3_3398_0_b(.in(layer_2[228]), .out(far_3_3398_0[1]));
    assign layer_3[338] = ~far_3_3398_0[0] | (far_3_3398_0[0] & far_3_3398_0[1]); 
    wire [1:0] far_3_3399_0;    relay_conn far_3_3399_0_a(.in(layer_2[737]), .out(far_3_3399_0[0]));    relay_conn far_3_3399_0_b(.in(layer_2[695]), .out(far_3_3399_0[1]));
    assign layer_3[339] = ~(far_3_3399_0[0] ^ far_3_3399_0[1]); 
    wire [1:0] far_3_3400_0;    relay_conn far_3_3400_0_a(.in(layer_2[794]), .out(far_3_3400_0[0]));    relay_conn far_3_3400_0_b(.in(layer_2[901]), .out(far_3_3400_0[1]));
    wire [1:0] far_3_3400_1;    relay_conn far_3_3400_1_a(.in(far_3_3400_0[0]), .out(far_3_3400_1[0]));    relay_conn far_3_3400_1_b(.in(far_3_3400_0[1]), .out(far_3_3400_1[1]));
    wire [1:0] far_3_3400_2;    relay_conn far_3_3400_2_a(.in(far_3_3400_1[0]), .out(far_3_3400_2[0]));    relay_conn far_3_3400_2_b(.in(far_3_3400_1[1]), .out(far_3_3400_2[1]));
    assign layer_3[340] = far_3_3400_2[0] | far_3_3400_2[1]; 
    wire [1:0] far_3_3401_0;    relay_conn far_3_3401_0_a(.in(layer_2[371]), .out(far_3_3401_0[0]));    relay_conn far_3_3401_0_b(.in(layer_2[328]), .out(far_3_3401_0[1]));
    assign layer_3[341] = ~far_3_3401_0[0]; 
    assign layer_3[342] = layer_2[43] & ~layer_2[32]; 
    assign layer_3[343] = ~layer_2[978] | (layer_2[978] & layer_2[969]); 
    wire [1:0] far_3_3404_0;    relay_conn far_3_3404_0_a(.in(layer_2[138]), .out(far_3_3404_0[0]));    relay_conn far_3_3404_0_b(.in(layer_2[188]), .out(far_3_3404_0[1]));
    assign layer_3[344] = far_3_3404_0[0] & ~far_3_3404_0[1]; 
    wire [1:0] far_3_3405_0;    relay_conn far_3_3405_0_a(.in(layer_2[183]), .out(far_3_3405_0[0]));    relay_conn far_3_3405_0_b(.in(layer_2[142]), .out(far_3_3405_0[1]));
    assign layer_3[345] = ~(far_3_3405_0[0] | far_3_3405_0[1]); 
    wire [1:0] far_3_3406_0;    relay_conn far_3_3406_0_a(.in(layer_2[141]), .out(far_3_3406_0[0]));    relay_conn far_3_3406_0_b(.in(layer_2[177]), .out(far_3_3406_0[1]));
    assign layer_3[346] = far_3_3406_0[0] | far_3_3406_0[1]; 
    wire [1:0] far_3_3407_0;    relay_conn far_3_3407_0_a(.in(layer_2[950]), .out(far_3_3407_0[0]));    relay_conn far_3_3407_0_b(.in(layer_2[825]), .out(far_3_3407_0[1]));
    wire [1:0] far_3_3407_1;    relay_conn far_3_3407_1_a(.in(far_3_3407_0[0]), .out(far_3_3407_1[0]));    relay_conn far_3_3407_1_b(.in(far_3_3407_0[1]), .out(far_3_3407_1[1]));
    wire [1:0] far_3_3407_2;    relay_conn far_3_3407_2_a(.in(far_3_3407_1[0]), .out(far_3_3407_2[0]));    relay_conn far_3_3407_2_b(.in(far_3_3407_1[1]), .out(far_3_3407_2[1]));
    assign layer_3[347] = far_3_3407_2[0]; 
    wire [1:0] far_3_3408_0;    relay_conn far_3_3408_0_a(.in(layer_2[315]), .out(far_3_3408_0[0]));    relay_conn far_3_3408_0_b(.in(layer_2[361]), .out(far_3_3408_0[1]));
    assign layer_3[348] = far_3_3408_0[0]; 
    wire [1:0] far_3_3409_0;    relay_conn far_3_3409_0_a(.in(layer_2[438]), .out(far_3_3409_0[0]));    relay_conn far_3_3409_0_b(.in(layer_2[376]), .out(far_3_3409_0[1]));
    assign layer_3[349] = ~far_3_3409_0[1] | (far_3_3409_0[0] & far_3_3409_0[1]); 
    wire [1:0] far_3_3410_0;    relay_conn far_3_3410_0_a(.in(layer_2[742]), .out(far_3_3410_0[0]));    relay_conn far_3_3410_0_b(.in(layer_2[683]), .out(far_3_3410_0[1]));
    assign layer_3[350] = far_3_3410_0[0] | far_3_3410_0[1]; 
    assign layer_3[351] = layer_2[401] | layer_2[376]; 
    wire [1:0] far_3_3412_0;    relay_conn far_3_3412_0_a(.in(layer_2[143]), .out(far_3_3412_0[0]));    relay_conn far_3_3412_0_b(.in(layer_2[263]), .out(far_3_3412_0[1]));
    wire [1:0] far_3_3412_1;    relay_conn far_3_3412_1_a(.in(far_3_3412_0[0]), .out(far_3_3412_1[0]));    relay_conn far_3_3412_1_b(.in(far_3_3412_0[1]), .out(far_3_3412_1[1]));
    wire [1:0] far_3_3412_2;    relay_conn far_3_3412_2_a(.in(far_3_3412_1[0]), .out(far_3_3412_2[0]));    relay_conn far_3_3412_2_b(.in(far_3_3412_1[1]), .out(far_3_3412_2[1]));
    assign layer_3[352] = ~far_3_3412_2[1]; 
    wire [1:0] far_3_3413_0;    relay_conn far_3_3413_0_a(.in(layer_2[120]), .out(far_3_3413_0[0]));    relay_conn far_3_3413_0_b(.in(layer_2[237]), .out(far_3_3413_0[1]));
    wire [1:0] far_3_3413_1;    relay_conn far_3_3413_1_a(.in(far_3_3413_0[0]), .out(far_3_3413_1[0]));    relay_conn far_3_3413_1_b(.in(far_3_3413_0[1]), .out(far_3_3413_1[1]));
    wire [1:0] far_3_3413_2;    relay_conn far_3_3413_2_a(.in(far_3_3413_1[0]), .out(far_3_3413_2[0]));    relay_conn far_3_3413_2_b(.in(far_3_3413_1[1]), .out(far_3_3413_2[1]));
    assign layer_3[353] = ~far_3_3413_2[1]; 
    wire [1:0] far_3_3414_0;    relay_conn far_3_3414_0_a(.in(layer_2[1007]), .out(far_3_3414_0[0]));    relay_conn far_3_3414_0_b(.in(layer_2[926]), .out(far_3_3414_0[1]));
    wire [1:0] far_3_3414_1;    relay_conn far_3_3414_1_a(.in(far_3_3414_0[0]), .out(far_3_3414_1[0]));    relay_conn far_3_3414_1_b(.in(far_3_3414_0[1]), .out(far_3_3414_1[1]));
    assign layer_3[354] = ~far_3_3414_1[1] | (far_3_3414_1[0] & far_3_3414_1[1]); 
    assign layer_3[355] = layer_2[934] & ~layer_2[925]; 
    wire [1:0] far_3_3416_0;    relay_conn far_3_3416_0_a(.in(layer_2[620]), .out(far_3_3416_0[0]));    relay_conn far_3_3416_0_b(.in(layer_2[513]), .out(far_3_3416_0[1]));
    wire [1:0] far_3_3416_1;    relay_conn far_3_3416_1_a(.in(far_3_3416_0[0]), .out(far_3_3416_1[0]));    relay_conn far_3_3416_1_b(.in(far_3_3416_0[1]), .out(far_3_3416_1[1]));
    wire [1:0] far_3_3416_2;    relay_conn far_3_3416_2_a(.in(far_3_3416_1[0]), .out(far_3_3416_2[0]));    relay_conn far_3_3416_2_b(.in(far_3_3416_1[1]), .out(far_3_3416_2[1]));
    assign layer_3[356] = ~(far_3_3416_2[0] ^ far_3_3416_2[1]); 
    assign layer_3[357] = layer_2[768] | layer_2[758]; 
    wire [1:0] far_3_3418_0;    relay_conn far_3_3418_0_a(.in(layer_2[32]), .out(far_3_3418_0[0]));    relay_conn far_3_3418_0_b(.in(layer_2[112]), .out(far_3_3418_0[1]));
    wire [1:0] far_3_3418_1;    relay_conn far_3_3418_1_a(.in(far_3_3418_0[0]), .out(far_3_3418_1[0]));    relay_conn far_3_3418_1_b(.in(far_3_3418_0[1]), .out(far_3_3418_1[1]));
    assign layer_3[358] = far_3_3418_1[0]; 
    wire [1:0] far_3_3419_0;    relay_conn far_3_3419_0_a(.in(layer_2[52]), .out(far_3_3419_0[0]));    relay_conn far_3_3419_0_b(.in(layer_2[10]), .out(far_3_3419_0[1]));
    assign layer_3[359] = far_3_3419_0[0]; 
    wire [1:0] far_3_3420_0;    relay_conn far_3_3420_0_a(.in(layer_2[826]), .out(far_3_3420_0[0]));    relay_conn far_3_3420_0_b(.in(layer_2[949]), .out(far_3_3420_0[1]));
    wire [1:0] far_3_3420_1;    relay_conn far_3_3420_1_a(.in(far_3_3420_0[0]), .out(far_3_3420_1[0]));    relay_conn far_3_3420_1_b(.in(far_3_3420_0[1]), .out(far_3_3420_1[1]));
    wire [1:0] far_3_3420_2;    relay_conn far_3_3420_2_a(.in(far_3_3420_1[0]), .out(far_3_3420_2[0]));    relay_conn far_3_3420_2_b(.in(far_3_3420_1[1]), .out(far_3_3420_2[1]));
    assign layer_3[360] = far_3_3420_2[0] & ~far_3_3420_2[1]; 
    assign layer_3[361] = ~(layer_2[849] & layer_2[872]); 
    assign layer_3[362] = layer_2[109] & layer_2[103]; 
    wire [1:0] far_3_3423_0;    relay_conn far_3_3423_0_a(.in(layer_2[422]), .out(far_3_3423_0[0]));    relay_conn far_3_3423_0_b(.in(layer_2[487]), .out(far_3_3423_0[1]));
    wire [1:0] far_3_3423_1;    relay_conn far_3_3423_1_a(.in(far_3_3423_0[0]), .out(far_3_3423_1[0]));    relay_conn far_3_3423_1_b(.in(far_3_3423_0[1]), .out(far_3_3423_1[1]));
    assign layer_3[363] = ~far_3_3423_1[1]; 
    wire [1:0] far_3_3424_0;    relay_conn far_3_3424_0_a(.in(layer_2[706]), .out(far_3_3424_0[0]));    relay_conn far_3_3424_0_b(.in(layer_2[758]), .out(far_3_3424_0[1]));
    assign layer_3[364] = far_3_3424_0[1]; 
    wire [1:0] far_3_3425_0;    relay_conn far_3_3425_0_a(.in(layer_2[910]), .out(far_3_3425_0[0]));    relay_conn far_3_3425_0_b(.in(layer_2[956]), .out(far_3_3425_0[1]));
    assign layer_3[365] = far_3_3425_0[0]; 
    assign layer_3[366] = ~layer_2[971]; 
    assign layer_3[367] = layer_2[1005]; 
    wire [1:0] far_3_3428_0;    relay_conn far_3_3428_0_a(.in(layer_2[880]), .out(far_3_3428_0[0]));    relay_conn far_3_3428_0_b(.in(layer_2[913]), .out(far_3_3428_0[1]));
    assign layer_3[368] = far_3_3428_0[0] & far_3_3428_0[1]; 
    wire [1:0] far_3_3429_0;    relay_conn far_3_3429_0_a(.in(layer_2[32]), .out(far_3_3429_0[0]));    relay_conn far_3_3429_0_b(.in(layer_2[78]), .out(far_3_3429_0[1]));
    assign layer_3[369] = far_3_3429_0[0] | far_3_3429_0[1]; 
    wire [1:0] far_3_3430_0;    relay_conn far_3_3430_0_a(.in(layer_2[1]), .out(far_3_3430_0[0]));    relay_conn far_3_3430_0_b(.in(layer_2[86]), .out(far_3_3430_0[1]));
    wire [1:0] far_3_3430_1;    relay_conn far_3_3430_1_a(.in(far_3_3430_0[0]), .out(far_3_3430_1[0]));    relay_conn far_3_3430_1_b(.in(far_3_3430_0[1]), .out(far_3_3430_1[1]));
    assign layer_3[370] = ~far_3_3430_1[1]; 
    assign layer_3[371] = ~(layer_2[10] & layer_2[1]); 
    wire [1:0] far_3_3432_0;    relay_conn far_3_3432_0_a(.in(layer_2[845]), .out(far_3_3432_0[0]));    relay_conn far_3_3432_0_b(.in(layer_2[963]), .out(far_3_3432_0[1]));
    wire [1:0] far_3_3432_1;    relay_conn far_3_3432_1_a(.in(far_3_3432_0[0]), .out(far_3_3432_1[0]));    relay_conn far_3_3432_1_b(.in(far_3_3432_0[1]), .out(far_3_3432_1[1]));
    wire [1:0] far_3_3432_2;    relay_conn far_3_3432_2_a(.in(far_3_3432_1[0]), .out(far_3_3432_2[0]));    relay_conn far_3_3432_2_b(.in(far_3_3432_1[1]), .out(far_3_3432_2[1]));
    assign layer_3[372] = ~far_3_3432_2[0] | (far_3_3432_2[0] & far_3_3432_2[1]); 
    assign layer_3[373] = ~layer_2[138] | (layer_2[138] & layer_2[155]); 
    wire [1:0] far_3_3434_0;    relay_conn far_3_3434_0_a(.in(layer_2[106]), .out(far_3_3434_0[0]));    relay_conn far_3_3434_0_b(.in(layer_2[56]), .out(far_3_3434_0[1]));
    assign layer_3[374] = ~far_3_3434_0[1] | (far_3_3434_0[0] & far_3_3434_0[1]); 
    assign layer_3[375] = ~layer_2[971] | (layer_2[971] & layer_2[965]); 
    wire [1:0] far_3_3436_0;    relay_conn far_3_3436_0_a(.in(layer_2[298]), .out(far_3_3436_0[0]));    relay_conn far_3_3436_0_b(.in(layer_2[207]), .out(far_3_3436_0[1]));
    wire [1:0] far_3_3436_1;    relay_conn far_3_3436_1_a(.in(far_3_3436_0[0]), .out(far_3_3436_1[0]));    relay_conn far_3_3436_1_b(.in(far_3_3436_0[1]), .out(far_3_3436_1[1]));
    assign layer_3[376] = ~far_3_3436_1[0] | (far_3_3436_1[0] & far_3_3436_1[1]); 
    wire [1:0] far_3_3437_0;    relay_conn far_3_3437_0_a(.in(layer_2[547]), .out(far_3_3437_0[0]));    relay_conn far_3_3437_0_b(.in(layer_2[511]), .out(far_3_3437_0[1]));
    assign layer_3[377] = ~(far_3_3437_0[0] & far_3_3437_0[1]); 
    wire [1:0] far_3_3438_0;    relay_conn far_3_3438_0_a(.in(layer_2[845]), .out(far_3_3438_0[0]));    relay_conn far_3_3438_0_b(.in(layer_2[813]), .out(far_3_3438_0[1]));
    assign layer_3[378] = ~(far_3_3438_0[0] & far_3_3438_0[1]); 
    wire [1:0] far_3_3439_0;    relay_conn far_3_3439_0_a(.in(layer_2[287]), .out(far_3_3439_0[0]));    relay_conn far_3_3439_0_b(.in(layer_2[366]), .out(far_3_3439_0[1]));
    wire [1:0] far_3_3439_1;    relay_conn far_3_3439_1_a(.in(far_3_3439_0[0]), .out(far_3_3439_1[0]));    relay_conn far_3_3439_1_b(.in(far_3_3439_0[1]), .out(far_3_3439_1[1]));
    assign layer_3[379] = far_3_3439_1[0] ^ far_3_3439_1[1]; 
    assign layer_3[380] = ~layer_2[352] | (layer_2[362] & layer_2[352]); 
    wire [1:0] far_3_3441_0;    relay_conn far_3_3441_0_a(.in(layer_2[578]), .out(far_3_3441_0[0]));    relay_conn far_3_3441_0_b(.in(layer_2[514]), .out(far_3_3441_0[1]));
    wire [1:0] far_3_3441_1;    relay_conn far_3_3441_1_a(.in(far_3_3441_0[0]), .out(far_3_3441_1[0]));    relay_conn far_3_3441_1_b(.in(far_3_3441_0[1]), .out(far_3_3441_1[1]));
    assign layer_3[381] = ~far_3_3441_1[1]; 
    assign layer_3[382] = layer_2[335]; 
    wire [1:0] far_3_3443_0;    relay_conn far_3_3443_0_a(.in(layer_2[644]), .out(far_3_3443_0[0]));    relay_conn far_3_3443_0_b(.in(layer_2[735]), .out(far_3_3443_0[1]));
    wire [1:0] far_3_3443_1;    relay_conn far_3_3443_1_a(.in(far_3_3443_0[0]), .out(far_3_3443_1[0]));    relay_conn far_3_3443_1_b(.in(far_3_3443_0[1]), .out(far_3_3443_1[1]));
    assign layer_3[383] = far_3_3443_1[0]; 
    assign layer_3[384] = layer_2[857] | layer_2[871]; 
    wire [1:0] far_3_3445_0;    relay_conn far_3_3445_0_a(.in(layer_2[922]), .out(far_3_3445_0[0]));    relay_conn far_3_3445_0_b(.in(layer_2[1011]), .out(far_3_3445_0[1]));
    wire [1:0] far_3_3445_1;    relay_conn far_3_3445_1_a(.in(far_3_3445_0[0]), .out(far_3_3445_1[0]));    relay_conn far_3_3445_1_b(.in(far_3_3445_0[1]), .out(far_3_3445_1[1]));
    assign layer_3[385] = far_3_3445_1[0] | far_3_3445_1[1]; 
    wire [1:0] far_3_3446_0;    relay_conn far_3_3446_0_a(.in(layer_2[370]), .out(far_3_3446_0[0]));    relay_conn far_3_3446_0_b(.in(layer_2[281]), .out(far_3_3446_0[1]));
    wire [1:0] far_3_3446_1;    relay_conn far_3_3446_1_a(.in(far_3_3446_0[0]), .out(far_3_3446_1[0]));    relay_conn far_3_3446_1_b(.in(far_3_3446_0[1]), .out(far_3_3446_1[1]));
    assign layer_3[386] = ~(far_3_3446_1[0] & far_3_3446_1[1]); 
    wire [1:0] far_3_3447_0;    relay_conn far_3_3447_0_a(.in(layer_2[182]), .out(far_3_3447_0[0]));    relay_conn far_3_3447_0_b(.in(layer_2[218]), .out(far_3_3447_0[1]));
    assign layer_3[387] = ~(far_3_3447_0[0] ^ far_3_3447_0[1]); 
    assign layer_3[388] = ~layer_2[840]; 
    wire [1:0] far_3_3449_0;    relay_conn far_3_3449_0_a(.in(layer_2[366]), .out(far_3_3449_0[0]));    relay_conn far_3_3449_0_b(.in(layer_2[471]), .out(far_3_3449_0[1]));
    wire [1:0] far_3_3449_1;    relay_conn far_3_3449_1_a(.in(far_3_3449_0[0]), .out(far_3_3449_1[0]));    relay_conn far_3_3449_1_b(.in(far_3_3449_0[1]), .out(far_3_3449_1[1]));
    wire [1:0] far_3_3449_2;    relay_conn far_3_3449_2_a(.in(far_3_3449_1[0]), .out(far_3_3449_2[0]));    relay_conn far_3_3449_2_b(.in(far_3_3449_1[1]), .out(far_3_3449_2[1]));
    assign layer_3[389] = ~(far_3_3449_2[0] | far_3_3449_2[1]); 
    wire [1:0] far_3_3450_0;    relay_conn far_3_3450_0_a(.in(layer_2[520]), .out(far_3_3450_0[0]));    relay_conn far_3_3450_0_b(.in(layer_2[421]), .out(far_3_3450_0[1]));
    wire [1:0] far_3_3450_1;    relay_conn far_3_3450_1_a(.in(far_3_3450_0[0]), .out(far_3_3450_1[0]));    relay_conn far_3_3450_1_b(.in(far_3_3450_0[1]), .out(far_3_3450_1[1]));
    wire [1:0] far_3_3450_2;    relay_conn far_3_3450_2_a(.in(far_3_3450_1[0]), .out(far_3_3450_2[0]));    relay_conn far_3_3450_2_b(.in(far_3_3450_1[1]), .out(far_3_3450_2[1]));
    assign layer_3[390] = ~far_3_3450_2[0]; 
    assign layer_3[391] = layer_2[649]; 
    wire [1:0] far_3_3452_0;    relay_conn far_3_3452_0_a(.in(layer_2[510]), .out(far_3_3452_0[0]));    relay_conn far_3_3452_0_b(.in(layer_2[577]), .out(far_3_3452_0[1]));
    wire [1:0] far_3_3452_1;    relay_conn far_3_3452_1_a(.in(far_3_3452_0[0]), .out(far_3_3452_1[0]));    relay_conn far_3_3452_1_b(.in(far_3_3452_0[1]), .out(far_3_3452_1[1]));
    assign layer_3[392] = far_3_3452_1[1] & ~far_3_3452_1[0]; 
    wire [1:0] far_3_3453_0;    relay_conn far_3_3453_0_a(.in(layer_2[92]), .out(far_3_3453_0[0]));    relay_conn far_3_3453_0_b(.in(layer_2[124]), .out(far_3_3453_0[1]));
    assign layer_3[393] = ~(far_3_3453_0[0] | far_3_3453_0[1]); 
    wire [1:0] far_3_3454_0;    relay_conn far_3_3454_0_a(.in(layer_2[541]), .out(far_3_3454_0[0]));    relay_conn far_3_3454_0_b(.in(layer_2[651]), .out(far_3_3454_0[1]));
    wire [1:0] far_3_3454_1;    relay_conn far_3_3454_1_a(.in(far_3_3454_0[0]), .out(far_3_3454_1[0]));    relay_conn far_3_3454_1_b(.in(far_3_3454_0[1]), .out(far_3_3454_1[1]));
    wire [1:0] far_3_3454_2;    relay_conn far_3_3454_2_a(.in(far_3_3454_1[0]), .out(far_3_3454_2[0]));    relay_conn far_3_3454_2_b(.in(far_3_3454_1[1]), .out(far_3_3454_2[1]));
    assign layer_3[394] = ~far_3_3454_2[1] | (far_3_3454_2[0] & far_3_3454_2[1]); 
    assign layer_3[395] = layer_2[565]; 
    assign layer_3[396] = layer_2[880]; 
    wire [1:0] far_3_3457_0;    relay_conn far_3_3457_0_a(.in(layer_2[954]), .out(far_3_3457_0[0]));    relay_conn far_3_3457_0_b(.in(layer_2[859]), .out(far_3_3457_0[1]));
    wire [1:0] far_3_3457_1;    relay_conn far_3_3457_1_a(.in(far_3_3457_0[0]), .out(far_3_3457_1[0]));    relay_conn far_3_3457_1_b(.in(far_3_3457_0[1]), .out(far_3_3457_1[1]));
    assign layer_3[397] = ~far_3_3457_1[1] | (far_3_3457_1[0] & far_3_3457_1[1]); 
    assign layer_3[398] = ~layer_2[198]; 
    wire [1:0] far_3_3459_0;    relay_conn far_3_3459_0_a(.in(layer_2[48]), .out(far_3_3459_0[0]));    relay_conn far_3_3459_0_b(.in(layer_2[126]), .out(far_3_3459_0[1]));
    wire [1:0] far_3_3459_1;    relay_conn far_3_3459_1_a(.in(far_3_3459_0[0]), .out(far_3_3459_1[0]));    relay_conn far_3_3459_1_b(.in(far_3_3459_0[1]), .out(far_3_3459_1[1]));
    assign layer_3[399] = ~far_3_3459_1[1] | (far_3_3459_1[0] & far_3_3459_1[1]); 
    assign layer_3[400] = layer_2[209]; 
    wire [1:0] far_3_3461_0;    relay_conn far_3_3461_0_a(.in(layer_2[262]), .out(far_3_3461_0[0]));    relay_conn far_3_3461_0_b(.in(layer_2[357]), .out(far_3_3461_0[1]));
    wire [1:0] far_3_3461_1;    relay_conn far_3_3461_1_a(.in(far_3_3461_0[0]), .out(far_3_3461_1[0]));    relay_conn far_3_3461_1_b(.in(far_3_3461_0[1]), .out(far_3_3461_1[1]));
    assign layer_3[401] = far_3_3461_1[0]; 
    wire [1:0] far_3_3462_0;    relay_conn far_3_3462_0_a(.in(layer_2[84]), .out(far_3_3462_0[0]));    relay_conn far_3_3462_0_b(.in(layer_2[168]), .out(far_3_3462_0[1]));
    wire [1:0] far_3_3462_1;    relay_conn far_3_3462_1_a(.in(far_3_3462_0[0]), .out(far_3_3462_1[0]));    relay_conn far_3_3462_1_b(.in(far_3_3462_0[1]), .out(far_3_3462_1[1]));
    assign layer_3[402] = far_3_3462_1[0] & ~far_3_3462_1[1]; 
    assign layer_3[403] = layer_2[146] & ~layer_2[142]; 
    wire [1:0] far_3_3464_0;    relay_conn far_3_3464_0_a(.in(layer_2[254]), .out(far_3_3464_0[0]));    relay_conn far_3_3464_0_b(.in(layer_2[143]), .out(far_3_3464_0[1]));
    wire [1:0] far_3_3464_1;    relay_conn far_3_3464_1_a(.in(far_3_3464_0[0]), .out(far_3_3464_1[0]));    relay_conn far_3_3464_1_b(.in(far_3_3464_0[1]), .out(far_3_3464_1[1]));
    wire [1:0] far_3_3464_2;    relay_conn far_3_3464_2_a(.in(far_3_3464_1[0]), .out(far_3_3464_2[0]));    relay_conn far_3_3464_2_b(.in(far_3_3464_1[1]), .out(far_3_3464_2[1]));
    assign layer_3[404] = ~(far_3_3464_2[0] | far_3_3464_2[1]); 
    assign layer_3[405] = ~(layer_2[421] | layer_2[419]); 
    wire [1:0] far_3_3466_0;    relay_conn far_3_3466_0_a(.in(layer_2[338]), .out(far_3_3466_0[0]));    relay_conn far_3_3466_0_b(.in(layer_2[306]), .out(far_3_3466_0[1]));
    assign layer_3[406] = ~(far_3_3466_0[0] | far_3_3466_0[1]); 
    wire [1:0] far_3_3467_0;    relay_conn far_3_3467_0_a(.in(layer_2[951]), .out(far_3_3467_0[0]));    relay_conn far_3_3467_0_b(.in(layer_2[907]), .out(far_3_3467_0[1]));
    assign layer_3[407] = ~(far_3_3467_0[0] | far_3_3467_0[1]); 
    assign layer_3[408] = ~(layer_2[915] & layer_2[920]); 
    wire [1:0] far_3_3469_0;    relay_conn far_3_3469_0_a(.in(layer_2[164]), .out(far_3_3469_0[0]));    relay_conn far_3_3469_0_b(.in(layer_2[43]), .out(far_3_3469_0[1]));
    wire [1:0] far_3_3469_1;    relay_conn far_3_3469_1_a(.in(far_3_3469_0[0]), .out(far_3_3469_1[0]));    relay_conn far_3_3469_1_b(.in(far_3_3469_0[1]), .out(far_3_3469_1[1]));
    wire [1:0] far_3_3469_2;    relay_conn far_3_3469_2_a(.in(far_3_3469_1[0]), .out(far_3_3469_2[0]));    relay_conn far_3_3469_2_b(.in(far_3_3469_1[1]), .out(far_3_3469_2[1]));
    assign layer_3[409] = far_3_3469_2[0] & far_3_3469_2[1]; 
    wire [1:0] far_3_3470_0;    relay_conn far_3_3470_0_a(.in(layer_2[954]), .out(far_3_3470_0[0]));    relay_conn far_3_3470_0_b(.in(layer_2[870]), .out(far_3_3470_0[1]));
    wire [1:0] far_3_3470_1;    relay_conn far_3_3470_1_a(.in(far_3_3470_0[0]), .out(far_3_3470_1[0]));    relay_conn far_3_3470_1_b(.in(far_3_3470_0[1]), .out(far_3_3470_1[1]));
    assign layer_3[410] = ~far_3_3470_1[1]; 
    wire [1:0] far_3_3471_0;    relay_conn far_3_3471_0_a(.in(layer_2[370]), .out(far_3_3471_0[0]));    relay_conn far_3_3471_0_b(.in(layer_2[260]), .out(far_3_3471_0[1]));
    wire [1:0] far_3_3471_1;    relay_conn far_3_3471_1_a(.in(far_3_3471_0[0]), .out(far_3_3471_1[0]));    relay_conn far_3_3471_1_b(.in(far_3_3471_0[1]), .out(far_3_3471_1[1]));
    wire [1:0] far_3_3471_2;    relay_conn far_3_3471_2_a(.in(far_3_3471_1[0]), .out(far_3_3471_2[0]));    relay_conn far_3_3471_2_b(.in(far_3_3471_1[1]), .out(far_3_3471_2[1]));
    assign layer_3[411] = ~(far_3_3471_2[0] ^ far_3_3471_2[1]); 
    wire [1:0] far_3_3472_0;    relay_conn far_3_3472_0_a(.in(layer_2[680]), .out(far_3_3472_0[0]));    relay_conn far_3_3472_0_b(.in(layer_2[775]), .out(far_3_3472_0[1]));
    wire [1:0] far_3_3472_1;    relay_conn far_3_3472_1_a(.in(far_3_3472_0[0]), .out(far_3_3472_1[0]));    relay_conn far_3_3472_1_b(.in(far_3_3472_0[1]), .out(far_3_3472_1[1]));
    assign layer_3[412] = far_3_3472_1[1]; 
    wire [1:0] far_3_3473_0;    relay_conn far_3_3473_0_a(.in(layer_2[132]), .out(far_3_3473_0[0]));    relay_conn far_3_3473_0_b(.in(layer_2[100]), .out(far_3_3473_0[1]));
    assign layer_3[413] = far_3_3473_0[0] | far_3_3473_0[1]; 
    wire [1:0] far_3_3474_0;    relay_conn far_3_3474_0_a(.in(layer_2[412]), .out(far_3_3474_0[0]));    relay_conn far_3_3474_0_b(.in(layer_2[352]), .out(far_3_3474_0[1]));
    assign layer_3[414] = ~(far_3_3474_0[0] & far_3_3474_0[1]); 
    wire [1:0] far_3_3475_0;    relay_conn far_3_3475_0_a(.in(layer_2[361]), .out(far_3_3475_0[0]));    relay_conn far_3_3475_0_b(.in(layer_2[424]), .out(far_3_3475_0[1]));
    assign layer_3[415] = ~far_3_3475_0[1]; 
    wire [1:0] far_3_3476_0;    relay_conn far_3_3476_0_a(.in(layer_2[946]), .out(far_3_3476_0[0]));    relay_conn far_3_3476_0_b(.in(layer_2[844]), .out(far_3_3476_0[1]));
    wire [1:0] far_3_3476_1;    relay_conn far_3_3476_1_a(.in(far_3_3476_0[0]), .out(far_3_3476_1[0]));    relay_conn far_3_3476_1_b(.in(far_3_3476_0[1]), .out(far_3_3476_1[1]));
    wire [1:0] far_3_3476_2;    relay_conn far_3_3476_2_a(.in(far_3_3476_1[0]), .out(far_3_3476_2[0]));    relay_conn far_3_3476_2_b(.in(far_3_3476_1[1]), .out(far_3_3476_2[1]));
    assign layer_3[416] = ~(far_3_3476_2[0] | far_3_3476_2[1]); 
    wire [1:0] far_3_3477_0;    relay_conn far_3_3477_0_a(.in(layer_2[861]), .out(far_3_3477_0[0]));    relay_conn far_3_3477_0_b(.in(layer_2[909]), .out(far_3_3477_0[1]));
    assign layer_3[417] = ~far_3_3477_0[1] | (far_3_3477_0[0] & far_3_3477_0[1]); 
    assign layer_3[418] = layer_2[737] & ~layer_2[729]; 
    wire [1:0] far_3_3479_0;    relay_conn far_3_3479_0_a(.in(layer_2[872]), .out(far_3_3479_0[0]));    relay_conn far_3_3479_0_b(.in(layer_2[954]), .out(far_3_3479_0[1]));
    wire [1:0] far_3_3479_1;    relay_conn far_3_3479_1_a(.in(far_3_3479_0[0]), .out(far_3_3479_1[0]));    relay_conn far_3_3479_1_b(.in(far_3_3479_0[1]), .out(far_3_3479_1[1]));
    assign layer_3[419] = ~far_3_3479_1[1]; 
    wire [1:0] far_3_3480_0;    relay_conn far_3_3480_0_a(.in(layer_2[858]), .out(far_3_3480_0[0]));    relay_conn far_3_3480_0_b(.in(layer_2[762]), .out(far_3_3480_0[1]));
    wire [1:0] far_3_3480_1;    relay_conn far_3_3480_1_a(.in(far_3_3480_0[0]), .out(far_3_3480_1[0]));    relay_conn far_3_3480_1_b(.in(far_3_3480_0[1]), .out(far_3_3480_1[1]));
    wire [1:0] far_3_3480_2;    relay_conn far_3_3480_2_a(.in(far_3_3480_1[0]), .out(far_3_3480_2[0]));    relay_conn far_3_3480_2_b(.in(far_3_3480_1[1]), .out(far_3_3480_2[1]));
    assign layer_3[420] = ~far_3_3480_2[0] | (far_3_3480_2[0] & far_3_3480_2[1]); 
    assign layer_3[421] = ~(layer_2[262] & layer_2[292]); 
    wire [1:0] far_3_3482_0;    relay_conn far_3_3482_0_a(.in(layer_2[304]), .out(far_3_3482_0[0]));    relay_conn far_3_3482_0_b(.in(layer_2[195]), .out(far_3_3482_0[1]));
    wire [1:0] far_3_3482_1;    relay_conn far_3_3482_1_a(.in(far_3_3482_0[0]), .out(far_3_3482_1[0]));    relay_conn far_3_3482_1_b(.in(far_3_3482_0[1]), .out(far_3_3482_1[1]));
    wire [1:0] far_3_3482_2;    relay_conn far_3_3482_2_a(.in(far_3_3482_1[0]), .out(far_3_3482_2[0]));    relay_conn far_3_3482_2_b(.in(far_3_3482_1[1]), .out(far_3_3482_2[1]));
    assign layer_3[422] = ~(far_3_3482_2[0] | far_3_3482_2[1]); 
    wire [1:0] far_3_3483_0;    relay_conn far_3_3483_0_a(.in(layer_2[489]), .out(far_3_3483_0[0]));    relay_conn far_3_3483_0_b(.in(layer_2[583]), .out(far_3_3483_0[1]));
    wire [1:0] far_3_3483_1;    relay_conn far_3_3483_1_a(.in(far_3_3483_0[0]), .out(far_3_3483_1[0]));    relay_conn far_3_3483_1_b(.in(far_3_3483_0[1]), .out(far_3_3483_1[1]));
    assign layer_3[423] = ~(far_3_3483_1[0] | far_3_3483_1[1]); 
    wire [1:0] far_3_3484_0;    relay_conn far_3_3484_0_a(.in(layer_2[965]), .out(far_3_3484_0[0]));    relay_conn far_3_3484_0_b(.in(layer_2[876]), .out(far_3_3484_0[1]));
    wire [1:0] far_3_3484_1;    relay_conn far_3_3484_1_a(.in(far_3_3484_0[0]), .out(far_3_3484_1[0]));    relay_conn far_3_3484_1_b(.in(far_3_3484_0[1]), .out(far_3_3484_1[1]));
    assign layer_3[424] = far_3_3484_1[0] & ~far_3_3484_1[1]; 
    assign layer_3[425] = layer_2[992] & ~layer_2[1011]; 
    assign layer_3[426] = ~(layer_2[862] & layer_2[845]); 
    assign layer_3[427] = layer_2[595] & layer_2[575]; 
    wire [1:0] far_3_3488_0;    relay_conn far_3_3488_0_a(.in(layer_2[398]), .out(far_3_3488_0[0]));    relay_conn far_3_3488_0_b(.in(layer_2[499]), .out(far_3_3488_0[1]));
    wire [1:0] far_3_3488_1;    relay_conn far_3_3488_1_a(.in(far_3_3488_0[0]), .out(far_3_3488_1[0]));    relay_conn far_3_3488_1_b(.in(far_3_3488_0[1]), .out(far_3_3488_1[1]));
    wire [1:0] far_3_3488_2;    relay_conn far_3_3488_2_a(.in(far_3_3488_1[0]), .out(far_3_3488_2[0]));    relay_conn far_3_3488_2_b(.in(far_3_3488_1[1]), .out(far_3_3488_2[1]));
    assign layer_3[428] = far_3_3488_2[0] | far_3_3488_2[1]; 
    assign layer_3[429] = ~(layer_2[889] & layer_2[890]); 
    wire [1:0] far_3_3490_0;    relay_conn far_3_3490_0_a(.in(layer_2[915]), .out(far_3_3490_0[0]));    relay_conn far_3_3490_0_b(.in(layer_2[861]), .out(far_3_3490_0[1]));
    assign layer_3[430] = far_3_3490_0[1] & ~far_3_3490_0[0]; 
    assign layer_3[431] = layer_2[681] & ~layer_2[663]; 
    wire [1:0] far_3_3492_0;    relay_conn far_3_3492_0_a(.in(layer_2[855]), .out(far_3_3492_0[0]));    relay_conn far_3_3492_0_b(.in(layer_2[966]), .out(far_3_3492_0[1]));
    wire [1:0] far_3_3492_1;    relay_conn far_3_3492_1_a(.in(far_3_3492_0[0]), .out(far_3_3492_1[0]));    relay_conn far_3_3492_1_b(.in(far_3_3492_0[1]), .out(far_3_3492_1[1]));
    wire [1:0] far_3_3492_2;    relay_conn far_3_3492_2_a(.in(far_3_3492_1[0]), .out(far_3_3492_2[0]));    relay_conn far_3_3492_2_b(.in(far_3_3492_1[1]), .out(far_3_3492_2[1]));
    assign layer_3[432] = far_3_3492_2[0] | far_3_3492_2[1]; 
    wire [1:0] far_3_3493_0;    relay_conn far_3_3493_0_a(.in(layer_2[93]), .out(far_3_3493_0[0]));    relay_conn far_3_3493_0_b(.in(layer_2[48]), .out(far_3_3493_0[1]));
    assign layer_3[433] = far_3_3493_0[0]; 
    wire [1:0] far_3_3494_0;    relay_conn far_3_3494_0_a(.in(layer_2[132]), .out(far_3_3494_0[0]));    relay_conn far_3_3494_0_b(.in(layer_2[94]), .out(far_3_3494_0[1]));
    assign layer_3[434] = far_3_3494_0[0] & far_3_3494_0[1]; 
    wire [1:0] far_3_3495_0;    relay_conn far_3_3495_0_a(.in(layer_2[625]), .out(far_3_3495_0[0]));    relay_conn far_3_3495_0_b(.in(layer_2[691]), .out(far_3_3495_0[1]));
    wire [1:0] far_3_3495_1;    relay_conn far_3_3495_1_a(.in(far_3_3495_0[0]), .out(far_3_3495_1[0]));    relay_conn far_3_3495_1_b(.in(far_3_3495_0[1]), .out(far_3_3495_1[1]));
    assign layer_3[435] = ~far_3_3495_1[1]; 
    assign layer_3[436] = ~(layer_2[628] | layer_2[599]); 
    wire [1:0] far_3_3497_0;    relay_conn far_3_3497_0_a(.in(layer_2[132]), .out(far_3_3497_0[0]));    relay_conn far_3_3497_0_b(.in(layer_2[178]), .out(far_3_3497_0[1]));
    assign layer_3[437] = far_3_3497_0[0] & ~far_3_3497_0[1]; 
    wire [1:0] far_3_3498_0;    relay_conn far_3_3498_0_a(.in(layer_2[163]), .out(far_3_3498_0[0]));    relay_conn far_3_3498_0_b(.in(layer_2[265]), .out(far_3_3498_0[1]));
    wire [1:0] far_3_3498_1;    relay_conn far_3_3498_1_a(.in(far_3_3498_0[0]), .out(far_3_3498_1[0]));    relay_conn far_3_3498_1_b(.in(far_3_3498_0[1]), .out(far_3_3498_1[1]));
    wire [1:0] far_3_3498_2;    relay_conn far_3_3498_2_a(.in(far_3_3498_1[0]), .out(far_3_3498_2[0]));    relay_conn far_3_3498_2_b(.in(far_3_3498_1[1]), .out(far_3_3498_2[1]));
    assign layer_3[438] = ~(far_3_3498_2[0] & far_3_3498_2[1]); 
    wire [1:0] far_3_3499_0;    relay_conn far_3_3499_0_a(.in(layer_2[183]), .out(far_3_3499_0[0]));    relay_conn far_3_3499_0_b(.in(layer_2[300]), .out(far_3_3499_0[1]));
    wire [1:0] far_3_3499_1;    relay_conn far_3_3499_1_a(.in(far_3_3499_0[0]), .out(far_3_3499_1[0]));    relay_conn far_3_3499_1_b(.in(far_3_3499_0[1]), .out(far_3_3499_1[1]));
    wire [1:0] far_3_3499_2;    relay_conn far_3_3499_2_a(.in(far_3_3499_1[0]), .out(far_3_3499_2[0]));    relay_conn far_3_3499_2_b(.in(far_3_3499_1[1]), .out(far_3_3499_2[1]));
    assign layer_3[439] = ~far_3_3499_2[1] | (far_3_3499_2[0] & far_3_3499_2[1]); 
    assign layer_3[440] = layer_2[636]; 
    wire [1:0] far_3_3501_0;    relay_conn far_3_3501_0_a(.in(layer_2[399]), .out(far_3_3501_0[0]));    relay_conn far_3_3501_0_b(.in(layer_2[520]), .out(far_3_3501_0[1]));
    wire [1:0] far_3_3501_1;    relay_conn far_3_3501_1_a(.in(far_3_3501_0[0]), .out(far_3_3501_1[0]));    relay_conn far_3_3501_1_b(.in(far_3_3501_0[1]), .out(far_3_3501_1[1]));
    wire [1:0] far_3_3501_2;    relay_conn far_3_3501_2_a(.in(far_3_3501_1[0]), .out(far_3_3501_2[0]));    relay_conn far_3_3501_2_b(.in(far_3_3501_1[1]), .out(far_3_3501_2[1]));
    assign layer_3[441] = ~(far_3_3501_2[0] & far_3_3501_2[1]); 
    wire [1:0] far_3_3502_0;    relay_conn far_3_3502_0_a(.in(layer_2[410]), .out(far_3_3502_0[0]));    relay_conn far_3_3502_0_b(.in(layer_2[328]), .out(far_3_3502_0[1]));
    wire [1:0] far_3_3502_1;    relay_conn far_3_3502_1_a(.in(far_3_3502_0[0]), .out(far_3_3502_1[0]));    relay_conn far_3_3502_1_b(.in(far_3_3502_0[1]), .out(far_3_3502_1[1]));
    assign layer_3[442] = ~far_3_3502_1[1]; 
    wire [1:0] far_3_3503_0;    relay_conn far_3_3503_0_a(.in(layer_2[29]), .out(far_3_3503_0[0]));    relay_conn far_3_3503_0_b(.in(layer_2[94]), .out(far_3_3503_0[1]));
    wire [1:0] far_3_3503_1;    relay_conn far_3_3503_1_a(.in(far_3_3503_0[0]), .out(far_3_3503_1[0]));    relay_conn far_3_3503_1_b(.in(far_3_3503_0[1]), .out(far_3_3503_1[1]));
    assign layer_3[443] = ~far_3_3503_1[1]; 
    assign layer_3[444] = ~layer_2[92] | (layer_2[113] & layer_2[92]); 
    assign layer_3[445] = layer_2[852]; 
    assign layer_3[446] = ~layer_2[244]; 
    assign layer_3[447] = ~layer_2[790] | (layer_2[818] & layer_2[790]); 
    wire [1:0] far_3_3508_0;    relay_conn far_3_3508_0_a(.in(layer_2[749]), .out(far_3_3508_0[0]));    relay_conn far_3_3508_0_b(.in(layer_2[695]), .out(far_3_3508_0[1]));
    assign layer_3[448] = ~(far_3_3508_0[0] & far_3_3508_0[1]); 
    wire [1:0] far_3_3509_0;    relay_conn far_3_3509_0_a(.in(layer_2[716]), .out(far_3_3509_0[0]));    relay_conn far_3_3509_0_b(.in(layer_2[800]), .out(far_3_3509_0[1]));
    wire [1:0] far_3_3509_1;    relay_conn far_3_3509_1_a(.in(far_3_3509_0[0]), .out(far_3_3509_1[0]));    relay_conn far_3_3509_1_b(.in(far_3_3509_0[1]), .out(far_3_3509_1[1]));
    assign layer_3[449] = far_3_3509_1[1] & ~far_3_3509_1[0]; 
    wire [1:0] far_3_3510_0;    relay_conn far_3_3510_0_a(.in(layer_2[878]), .out(far_3_3510_0[0]));    relay_conn far_3_3510_0_b(.in(layer_2[791]), .out(far_3_3510_0[1]));
    wire [1:0] far_3_3510_1;    relay_conn far_3_3510_1_a(.in(far_3_3510_0[0]), .out(far_3_3510_1[0]));    relay_conn far_3_3510_1_b(.in(far_3_3510_0[1]), .out(far_3_3510_1[1]));
    assign layer_3[450] = far_3_3510_1[1]; 
    wire [1:0] far_3_3511_0;    relay_conn far_3_3511_0_a(.in(layer_2[418]), .out(far_3_3511_0[0]));    relay_conn far_3_3511_0_b(.in(layer_2[538]), .out(far_3_3511_0[1]));
    wire [1:0] far_3_3511_1;    relay_conn far_3_3511_1_a(.in(far_3_3511_0[0]), .out(far_3_3511_1[0]));    relay_conn far_3_3511_1_b(.in(far_3_3511_0[1]), .out(far_3_3511_1[1]));
    wire [1:0] far_3_3511_2;    relay_conn far_3_3511_2_a(.in(far_3_3511_1[0]), .out(far_3_3511_2[0]));    relay_conn far_3_3511_2_b(.in(far_3_3511_1[1]), .out(far_3_3511_2[1]));
    assign layer_3[451] = ~far_3_3511_2[1] | (far_3_3511_2[0] & far_3_3511_2[1]); 
    wire [1:0] far_3_3512_0;    relay_conn far_3_3512_0_a(.in(layer_2[144]), .out(far_3_3512_0[0]));    relay_conn far_3_3512_0_b(.in(layer_2[55]), .out(far_3_3512_0[1]));
    wire [1:0] far_3_3512_1;    relay_conn far_3_3512_1_a(.in(far_3_3512_0[0]), .out(far_3_3512_1[0]));    relay_conn far_3_3512_1_b(.in(far_3_3512_0[1]), .out(far_3_3512_1[1]));
    assign layer_3[452] = far_3_3512_1[0] & far_3_3512_1[1]; 
    wire [1:0] far_3_3513_0;    relay_conn far_3_3513_0_a(.in(layer_2[905]), .out(far_3_3513_0[0]));    relay_conn far_3_3513_0_b(.in(layer_2[859]), .out(far_3_3513_0[1]));
    assign layer_3[453] = far_3_3513_0[0] & far_3_3513_0[1]; 
    assign layer_3[454] = layer_2[277]; 
    assign layer_3[455] = ~layer_2[768]; 
    wire [1:0] far_3_3516_0;    relay_conn far_3_3516_0_a(.in(layer_2[702]), .out(far_3_3516_0[0]));    relay_conn far_3_3516_0_b(.in(layer_2[583]), .out(far_3_3516_0[1]));
    wire [1:0] far_3_3516_1;    relay_conn far_3_3516_1_a(.in(far_3_3516_0[0]), .out(far_3_3516_1[0]));    relay_conn far_3_3516_1_b(.in(far_3_3516_0[1]), .out(far_3_3516_1[1]));
    wire [1:0] far_3_3516_2;    relay_conn far_3_3516_2_a(.in(far_3_3516_1[0]), .out(far_3_3516_2[0]));    relay_conn far_3_3516_2_b(.in(far_3_3516_1[1]), .out(far_3_3516_2[1]));
    assign layer_3[456] = ~far_3_3516_2[1] | (far_3_3516_2[0] & far_3_3516_2[1]); 
    assign layer_3[457] = ~(layer_2[915] & layer_2[907]); 
    wire [1:0] far_3_3518_0;    relay_conn far_3_3518_0_a(.in(layer_2[845]), .out(far_3_3518_0[0]));    relay_conn far_3_3518_0_b(.in(layer_2[757]), .out(far_3_3518_0[1]));
    wire [1:0] far_3_3518_1;    relay_conn far_3_3518_1_a(.in(far_3_3518_0[0]), .out(far_3_3518_1[0]));    relay_conn far_3_3518_1_b(.in(far_3_3518_0[1]), .out(far_3_3518_1[1]));
    assign layer_3[458] = far_3_3518_1[0]; 
    wire [1:0] far_3_3519_0;    relay_conn far_3_3519_0_a(.in(layer_2[61]), .out(far_3_3519_0[0]));    relay_conn far_3_3519_0_b(.in(layer_2[138]), .out(far_3_3519_0[1]));
    wire [1:0] far_3_3519_1;    relay_conn far_3_3519_1_a(.in(far_3_3519_0[0]), .out(far_3_3519_1[0]));    relay_conn far_3_3519_1_b(.in(far_3_3519_0[1]), .out(far_3_3519_1[1]));
    assign layer_3[459] = far_3_3519_1[0] & far_3_3519_1[1]; 
    wire [1:0] far_3_3520_0;    relay_conn far_3_3520_0_a(.in(layer_2[818]), .out(far_3_3520_0[0]));    relay_conn far_3_3520_0_b(.in(layer_2[920]), .out(far_3_3520_0[1]));
    wire [1:0] far_3_3520_1;    relay_conn far_3_3520_1_a(.in(far_3_3520_0[0]), .out(far_3_3520_1[0]));    relay_conn far_3_3520_1_b(.in(far_3_3520_0[1]), .out(far_3_3520_1[1]));
    wire [1:0] far_3_3520_2;    relay_conn far_3_3520_2_a(.in(far_3_3520_1[0]), .out(far_3_3520_2[0]));    relay_conn far_3_3520_2_b(.in(far_3_3520_1[1]), .out(far_3_3520_2[1]));
    assign layer_3[460] = ~(far_3_3520_2[0] | far_3_3520_2[1]); 
    assign layer_3[461] = layer_2[390] & ~layer_2[370]; 
    assign layer_3[462] = layer_2[709]; 
    wire [1:0] far_3_3523_0;    relay_conn far_3_3523_0_a(.in(layer_2[250]), .out(far_3_3523_0[0]));    relay_conn far_3_3523_0_b(.in(layer_2[339]), .out(far_3_3523_0[1]));
    wire [1:0] far_3_3523_1;    relay_conn far_3_3523_1_a(.in(far_3_3523_0[0]), .out(far_3_3523_1[0]));    relay_conn far_3_3523_1_b(.in(far_3_3523_0[1]), .out(far_3_3523_1[1]));
    assign layer_3[463] = far_3_3523_1[1]; 
    wire [1:0] far_3_3524_0;    relay_conn far_3_3524_0_a(.in(layer_2[531]), .out(far_3_3524_0[0]));    relay_conn far_3_3524_0_b(.in(layer_2[641]), .out(far_3_3524_0[1]));
    wire [1:0] far_3_3524_1;    relay_conn far_3_3524_1_a(.in(far_3_3524_0[0]), .out(far_3_3524_1[0]));    relay_conn far_3_3524_1_b(.in(far_3_3524_0[1]), .out(far_3_3524_1[1]));
    wire [1:0] far_3_3524_2;    relay_conn far_3_3524_2_a(.in(far_3_3524_1[0]), .out(far_3_3524_2[0]));    relay_conn far_3_3524_2_b(.in(far_3_3524_1[1]), .out(far_3_3524_2[1]));
    assign layer_3[464] = ~far_3_3524_2[0] | (far_3_3524_2[0] & far_3_3524_2[1]); 
    wire [1:0] far_3_3525_0;    relay_conn far_3_3525_0_a(.in(layer_2[985]), .out(far_3_3525_0[0]));    relay_conn far_3_3525_0_b(.in(layer_2[926]), .out(far_3_3525_0[1]));
    assign layer_3[465] = ~far_3_3525_0[0] | (far_3_3525_0[0] & far_3_3525_0[1]); 
    wire [1:0] far_3_3526_0;    relay_conn far_3_3526_0_a(.in(layer_2[508]), .out(far_3_3526_0[0]));    relay_conn far_3_3526_0_b(.in(layer_2[421]), .out(far_3_3526_0[1]));
    wire [1:0] far_3_3526_1;    relay_conn far_3_3526_1_a(.in(far_3_3526_0[0]), .out(far_3_3526_1[0]));    relay_conn far_3_3526_1_b(.in(far_3_3526_0[1]), .out(far_3_3526_1[1]));
    assign layer_3[466] = far_3_3526_1[1] & ~far_3_3526_1[0]; 
    assign layer_3[467] = ~(layer_2[76] & layer_2[71]); 
    assign layer_3[468] = ~(layer_2[933] & layer_2[902]); 
    wire [1:0] far_3_3529_0;    relay_conn far_3_3529_0_a(.in(layer_2[1]), .out(far_3_3529_0[0]));    relay_conn far_3_3529_0_b(.in(layer_2[108]), .out(far_3_3529_0[1]));
    wire [1:0] far_3_3529_1;    relay_conn far_3_3529_1_a(.in(far_3_3529_0[0]), .out(far_3_3529_1[0]));    relay_conn far_3_3529_1_b(.in(far_3_3529_0[1]), .out(far_3_3529_1[1]));
    wire [1:0] far_3_3529_2;    relay_conn far_3_3529_2_a(.in(far_3_3529_1[0]), .out(far_3_3529_2[0]));    relay_conn far_3_3529_2_b(.in(far_3_3529_1[1]), .out(far_3_3529_2[1]));
    assign layer_3[469] = far_3_3529_2[1]; 
    wire [1:0] far_3_3530_0;    relay_conn far_3_3530_0_a(.in(layer_2[90]), .out(far_3_3530_0[0]));    relay_conn far_3_3530_0_b(.in(layer_2[18]), .out(far_3_3530_0[1]));
    wire [1:0] far_3_3530_1;    relay_conn far_3_3530_1_a(.in(far_3_3530_0[0]), .out(far_3_3530_1[0]));    relay_conn far_3_3530_1_b(.in(far_3_3530_0[1]), .out(far_3_3530_1[1]));
    assign layer_3[470] = ~far_3_3530_1[1] | (far_3_3530_1[0] & far_3_3530_1[1]); 
    wire [1:0] far_3_3531_0;    relay_conn far_3_3531_0_a(.in(layer_2[878]), .out(far_3_3531_0[0]));    relay_conn far_3_3531_0_b(.in(layer_2[920]), .out(far_3_3531_0[1]));
    assign layer_3[471] = ~(far_3_3531_0[0] & far_3_3531_0[1]); 
    assign layer_3[472] = layer_2[248] & ~layer_2[219]; 
    wire [1:0] far_3_3533_0;    relay_conn far_3_3533_0_a(.in(layer_2[670]), .out(far_3_3533_0[0]));    relay_conn far_3_3533_0_b(.in(layer_2[774]), .out(far_3_3533_0[1]));
    wire [1:0] far_3_3533_1;    relay_conn far_3_3533_1_a(.in(far_3_3533_0[0]), .out(far_3_3533_1[0]));    relay_conn far_3_3533_1_b(.in(far_3_3533_0[1]), .out(far_3_3533_1[1]));
    wire [1:0] far_3_3533_2;    relay_conn far_3_3533_2_a(.in(far_3_3533_1[0]), .out(far_3_3533_2[0]));    relay_conn far_3_3533_2_b(.in(far_3_3533_1[1]), .out(far_3_3533_2[1]));
    assign layer_3[473] = far_3_3533_2[0] ^ far_3_3533_2[1]; 
    assign layer_3[474] = ~layer_2[664] | (layer_2[673] & layer_2[664]); 
    wire [1:0] far_3_3535_0;    relay_conn far_3_3535_0_a(.in(layer_2[180]), .out(far_3_3535_0[0]));    relay_conn far_3_3535_0_b(.in(layer_2[287]), .out(far_3_3535_0[1]));
    wire [1:0] far_3_3535_1;    relay_conn far_3_3535_1_a(.in(far_3_3535_0[0]), .out(far_3_3535_1[0]));    relay_conn far_3_3535_1_b(.in(far_3_3535_0[1]), .out(far_3_3535_1[1]));
    wire [1:0] far_3_3535_2;    relay_conn far_3_3535_2_a(.in(far_3_3535_1[0]), .out(far_3_3535_2[0]));    relay_conn far_3_3535_2_b(.in(far_3_3535_1[1]), .out(far_3_3535_2[1]));
    assign layer_3[475] = far_3_3535_2[1]; 
    assign layer_3[476] = layer_2[208] & ~layer_2[221]; 
    assign layer_3[477] = ~layer_2[637]; 
    assign layer_3[478] = ~(layer_2[208] | layer_2[235]); 
    assign layer_3[479] = layer_2[824] ^ layer_2[794]; 
    assign layer_3[480] = layer_2[852] & ~layer_2[877]; 
    wire [1:0] far_3_3541_0;    relay_conn far_3_3541_0_a(.in(layer_2[1009]), .out(far_3_3541_0[0]));    relay_conn far_3_3541_0_b(.in(layer_2[934]), .out(far_3_3541_0[1]));
    wire [1:0] far_3_3541_1;    relay_conn far_3_3541_1_a(.in(far_3_3541_0[0]), .out(far_3_3541_1[0]));    relay_conn far_3_3541_1_b(.in(far_3_3541_0[1]), .out(far_3_3541_1[1]));
    assign layer_3[481] = far_3_3541_1[1] & ~far_3_3541_1[0]; 
    wire [1:0] far_3_3542_0;    relay_conn far_3_3542_0_a(.in(layer_2[859]), .out(far_3_3542_0[0]));    relay_conn far_3_3542_0_b(.in(layer_2[807]), .out(far_3_3542_0[1]));
    assign layer_3[482] = ~(far_3_3542_0[0] ^ far_3_3542_0[1]); 
    wire [1:0] far_3_3543_0;    relay_conn far_3_3543_0_a(.in(layer_2[813]), .out(far_3_3543_0[0]));    relay_conn far_3_3543_0_b(.in(layer_2[899]), .out(far_3_3543_0[1]));
    wire [1:0] far_3_3543_1;    relay_conn far_3_3543_1_a(.in(far_3_3543_0[0]), .out(far_3_3543_1[0]));    relay_conn far_3_3543_1_b(.in(far_3_3543_0[1]), .out(far_3_3543_1[1]));
    assign layer_3[483] = ~far_3_3543_1[0]; 
    assign layer_3[484] = layer_2[126] & ~layer_2[133]; 
    wire [1:0] far_3_3545_0;    relay_conn far_3_3545_0_a(.in(layer_2[50]), .out(far_3_3545_0[0]));    relay_conn far_3_3545_0_b(.in(layer_2[118]), .out(far_3_3545_0[1]));
    wire [1:0] far_3_3545_1;    relay_conn far_3_3545_1_a(.in(far_3_3545_0[0]), .out(far_3_3545_1[0]));    relay_conn far_3_3545_1_b(.in(far_3_3545_0[1]), .out(far_3_3545_1[1]));
    assign layer_3[485] = ~(far_3_3545_1[0] | far_3_3545_1[1]); 
    wire [1:0] far_3_3546_0;    relay_conn far_3_3546_0_a(.in(layer_2[741]), .out(far_3_3546_0[0]));    relay_conn far_3_3546_0_b(.in(layer_2[812]), .out(far_3_3546_0[1]));
    wire [1:0] far_3_3546_1;    relay_conn far_3_3546_1_a(.in(far_3_3546_0[0]), .out(far_3_3546_1[0]));    relay_conn far_3_3546_1_b(.in(far_3_3546_0[1]), .out(far_3_3546_1[1]));
    assign layer_3[486] = ~far_3_3546_1[1] | (far_3_3546_1[0] & far_3_3546_1[1]); 
    wire [1:0] far_3_3547_0;    relay_conn far_3_3547_0_a(.in(layer_2[347]), .out(far_3_3547_0[0]));    relay_conn far_3_3547_0_b(.in(layer_2[398]), .out(far_3_3547_0[1]));
    assign layer_3[487] = far_3_3547_0[0] ^ far_3_3547_0[1]; 
    assign layer_3[488] = layer_2[151] | layer_2[143]; 
    assign layer_3[489] = layer_2[50]; 
    wire [1:0] far_3_3550_0;    relay_conn far_3_3550_0_a(.in(layer_2[631]), .out(far_3_3550_0[0]));    relay_conn far_3_3550_0_b(.in(layer_2[741]), .out(far_3_3550_0[1]));
    wire [1:0] far_3_3550_1;    relay_conn far_3_3550_1_a(.in(far_3_3550_0[0]), .out(far_3_3550_1[0]));    relay_conn far_3_3550_1_b(.in(far_3_3550_0[1]), .out(far_3_3550_1[1]));
    wire [1:0] far_3_3550_2;    relay_conn far_3_3550_2_a(.in(far_3_3550_1[0]), .out(far_3_3550_2[0]));    relay_conn far_3_3550_2_b(.in(far_3_3550_1[1]), .out(far_3_3550_2[1]));
    assign layer_3[490] = far_3_3550_2[1]; 
    wire [1:0] far_3_3551_0;    relay_conn far_3_3551_0_a(.in(layer_2[371]), .out(far_3_3551_0[0]));    relay_conn far_3_3551_0_b(.in(layer_2[276]), .out(far_3_3551_0[1]));
    wire [1:0] far_3_3551_1;    relay_conn far_3_3551_1_a(.in(far_3_3551_0[0]), .out(far_3_3551_1[0]));    relay_conn far_3_3551_1_b(.in(far_3_3551_0[1]), .out(far_3_3551_1[1]));
    assign layer_3[491] = far_3_3551_1[0] & far_3_3551_1[1]; 
    wire [1:0] far_3_3552_0;    relay_conn far_3_3552_0_a(.in(layer_2[107]), .out(far_3_3552_0[0]));    relay_conn far_3_3552_0_b(.in(layer_2[178]), .out(far_3_3552_0[1]));
    wire [1:0] far_3_3552_1;    relay_conn far_3_3552_1_a(.in(far_3_3552_0[0]), .out(far_3_3552_1[0]));    relay_conn far_3_3552_1_b(.in(far_3_3552_0[1]), .out(far_3_3552_1[1]));
    assign layer_3[492] = far_3_3552_1[1] & ~far_3_3552_1[0]; 
    wire [1:0] far_3_3553_0;    relay_conn far_3_3553_0_a(.in(layer_2[623]), .out(far_3_3553_0[0]));    relay_conn far_3_3553_0_b(.in(layer_2[673]), .out(far_3_3553_0[1]));
    assign layer_3[493] = far_3_3553_0[0] ^ far_3_3553_0[1]; 
    assign layer_3[494] = layer_2[453] & ~layer_2[467]; 
    assign layer_3[495] = layer_2[205] & ~layer_2[235]; 
    wire [1:0] far_3_3556_0;    relay_conn far_3_3556_0_a(.in(layer_2[191]), .out(far_3_3556_0[0]));    relay_conn far_3_3556_0_b(.in(layer_2[304]), .out(far_3_3556_0[1]));
    wire [1:0] far_3_3556_1;    relay_conn far_3_3556_1_a(.in(far_3_3556_0[0]), .out(far_3_3556_1[0]));    relay_conn far_3_3556_1_b(.in(far_3_3556_0[1]), .out(far_3_3556_1[1]));
    wire [1:0] far_3_3556_2;    relay_conn far_3_3556_2_a(.in(far_3_3556_1[0]), .out(far_3_3556_2[0]));    relay_conn far_3_3556_2_b(.in(far_3_3556_1[1]), .out(far_3_3556_2[1]));
    assign layer_3[496] = far_3_3556_2[1] & ~far_3_3556_2[0]; 
    wire [1:0] far_3_3557_0;    relay_conn far_3_3557_0_a(.in(layer_2[663]), .out(far_3_3557_0[0]));    relay_conn far_3_3557_0_b(.in(layer_2[791]), .out(far_3_3557_0[1]));
    wire [1:0] far_3_3557_1;    relay_conn far_3_3557_1_a(.in(far_3_3557_0[0]), .out(far_3_3557_1[0]));    relay_conn far_3_3557_1_b(.in(far_3_3557_0[1]), .out(far_3_3557_1[1]));
    wire [1:0] far_3_3557_2;    relay_conn far_3_3557_2_a(.in(far_3_3557_1[0]), .out(far_3_3557_2[0]));    relay_conn far_3_3557_2_b(.in(far_3_3557_1[1]), .out(far_3_3557_2[1]));
    wire [1:0] far_3_3557_3;    relay_conn far_3_3557_3_a(.in(far_3_3557_2[0]), .out(far_3_3557_3[0]));    relay_conn far_3_3557_3_b(.in(far_3_3557_2[1]), .out(far_3_3557_3[1]));
    assign layer_3[497] = ~(far_3_3557_3[0] & far_3_3557_3[1]); 
    wire [1:0] far_3_3558_0;    relay_conn far_3_3558_0_a(.in(layer_2[463]), .out(far_3_3558_0[0]));    relay_conn far_3_3558_0_b(.in(layer_2[519]), .out(far_3_3558_0[1]));
    assign layer_3[498] = ~(far_3_3558_0[0] & far_3_3558_0[1]); 
    wire [1:0] far_3_3559_0;    relay_conn far_3_3559_0_a(.in(layer_2[627]), .out(far_3_3559_0[0]));    relay_conn far_3_3559_0_b(.in(layer_2[661]), .out(far_3_3559_0[1]));
    assign layer_3[499] = ~(far_3_3559_0[0] & far_3_3559_0[1]); 
    wire [1:0] far_3_3560_0;    relay_conn far_3_3560_0_a(.in(layer_2[1005]), .out(far_3_3560_0[0]));    relay_conn far_3_3560_0_b(.in(layer_2[916]), .out(far_3_3560_0[1]));
    wire [1:0] far_3_3560_1;    relay_conn far_3_3560_1_a(.in(far_3_3560_0[0]), .out(far_3_3560_1[0]));    relay_conn far_3_3560_1_b(.in(far_3_3560_0[1]), .out(far_3_3560_1[1]));
    assign layer_3[500] = ~far_3_3560_1[0] | (far_3_3560_1[0] & far_3_3560_1[1]); 
    wire [1:0] far_3_3561_0;    relay_conn far_3_3561_0_a(.in(layer_2[714]), .out(far_3_3561_0[0]));    relay_conn far_3_3561_0_b(.in(layer_2[777]), .out(far_3_3561_0[1]));
    assign layer_3[501] = ~(far_3_3561_0[0] & far_3_3561_0[1]); 
    assign layer_3[502] = ~(layer_2[654] | layer_2[626]); 
    wire [1:0] far_3_3563_0;    relay_conn far_3_3563_0_a(.in(layer_2[791]), .out(far_3_3563_0[0]));    relay_conn far_3_3563_0_b(.in(layer_2[891]), .out(far_3_3563_0[1]));
    wire [1:0] far_3_3563_1;    relay_conn far_3_3563_1_a(.in(far_3_3563_0[0]), .out(far_3_3563_1[0]));    relay_conn far_3_3563_1_b(.in(far_3_3563_0[1]), .out(far_3_3563_1[1]));
    wire [1:0] far_3_3563_2;    relay_conn far_3_3563_2_a(.in(far_3_3563_1[0]), .out(far_3_3563_2[0]));    relay_conn far_3_3563_2_b(.in(far_3_3563_1[1]), .out(far_3_3563_2[1]));
    assign layer_3[503] = far_3_3563_2[1] & ~far_3_3563_2[0]; 
    wire [1:0] far_3_3564_0;    relay_conn far_3_3564_0_a(.in(layer_2[423]), .out(far_3_3564_0[0]));    relay_conn far_3_3564_0_b(.in(layer_2[307]), .out(far_3_3564_0[1]));
    wire [1:0] far_3_3564_1;    relay_conn far_3_3564_1_a(.in(far_3_3564_0[0]), .out(far_3_3564_1[0]));    relay_conn far_3_3564_1_b(.in(far_3_3564_0[1]), .out(far_3_3564_1[1]));
    wire [1:0] far_3_3564_2;    relay_conn far_3_3564_2_a(.in(far_3_3564_1[0]), .out(far_3_3564_2[0]));    relay_conn far_3_3564_2_b(.in(far_3_3564_1[1]), .out(far_3_3564_2[1]));
    assign layer_3[504] = far_3_3564_2[0] & ~far_3_3564_2[1]; 
    wire [1:0] far_3_3565_0;    relay_conn far_3_3565_0_a(.in(layer_2[134]), .out(far_3_3565_0[0]));    relay_conn far_3_3565_0_b(.in(layer_2[52]), .out(far_3_3565_0[1]));
    wire [1:0] far_3_3565_1;    relay_conn far_3_3565_1_a(.in(far_3_3565_0[0]), .out(far_3_3565_1[0]));    relay_conn far_3_3565_1_b(.in(far_3_3565_0[1]), .out(far_3_3565_1[1]));
    assign layer_3[505] = ~(far_3_3565_1[0] & far_3_3565_1[1]); 
    wire [1:0] far_3_3566_0;    relay_conn far_3_3566_0_a(.in(layer_2[496]), .out(far_3_3566_0[0]));    relay_conn far_3_3566_0_b(.in(layer_2[433]), .out(far_3_3566_0[1]));
    assign layer_3[506] = ~(far_3_3566_0[0] | far_3_3566_0[1]); 
    assign layer_3[507] = layer_2[374] & layer_2[380]; 
    wire [1:0] far_3_3568_0;    relay_conn far_3_3568_0_a(.in(layer_2[670]), .out(far_3_3568_0[0]));    relay_conn far_3_3568_0_b(.in(layer_2[761]), .out(far_3_3568_0[1]));
    wire [1:0] far_3_3568_1;    relay_conn far_3_3568_1_a(.in(far_3_3568_0[0]), .out(far_3_3568_1[0]));    relay_conn far_3_3568_1_b(.in(far_3_3568_0[1]), .out(far_3_3568_1[1]));
    assign layer_3[508] = far_3_3568_1[1]; 
    wire [1:0] far_3_3569_0;    relay_conn far_3_3569_0_a(.in(layer_2[509]), .out(far_3_3569_0[0]));    relay_conn far_3_3569_0_b(.in(layer_2[434]), .out(far_3_3569_0[1]));
    wire [1:0] far_3_3569_1;    relay_conn far_3_3569_1_a(.in(far_3_3569_0[0]), .out(far_3_3569_1[0]));    relay_conn far_3_3569_1_b(.in(far_3_3569_0[1]), .out(far_3_3569_1[1]));
    assign layer_3[509] = far_3_3569_1[0] & ~far_3_3569_1[1]; 
    wire [1:0] far_3_3570_0;    relay_conn far_3_3570_0_a(.in(layer_2[75]), .out(far_3_3570_0[0]));    relay_conn far_3_3570_0_b(.in(layer_2[140]), .out(far_3_3570_0[1]));
    wire [1:0] far_3_3570_1;    relay_conn far_3_3570_1_a(.in(far_3_3570_0[0]), .out(far_3_3570_1[0]));    relay_conn far_3_3570_1_b(.in(far_3_3570_0[1]), .out(far_3_3570_1[1]));
    assign layer_3[510] = far_3_3570_1[0] ^ far_3_3570_1[1]; 
    wire [1:0] far_3_3571_0;    relay_conn far_3_3571_0_a(.in(layer_2[4]), .out(far_3_3571_0[0]));    relay_conn far_3_3571_0_b(.in(layer_2[54]), .out(far_3_3571_0[1]));
    assign layer_3[511] = far_3_3571_0[0] & far_3_3571_0[1]; 
    wire [1:0] far_3_3572_0;    relay_conn far_3_3572_0_a(.in(layer_2[126]), .out(far_3_3572_0[0]));    relay_conn far_3_3572_0_b(.in(layer_2[56]), .out(far_3_3572_0[1]));
    wire [1:0] far_3_3572_1;    relay_conn far_3_3572_1_a(.in(far_3_3572_0[0]), .out(far_3_3572_1[0]));    relay_conn far_3_3572_1_b(.in(far_3_3572_0[1]), .out(far_3_3572_1[1]));
    assign layer_3[512] = far_3_3572_1[1]; 
    wire [1:0] far_3_3573_0;    relay_conn far_3_3573_0_a(.in(layer_2[25]), .out(far_3_3573_0[0]));    relay_conn far_3_3573_0_b(.in(layer_2[120]), .out(far_3_3573_0[1]));
    wire [1:0] far_3_3573_1;    relay_conn far_3_3573_1_a(.in(far_3_3573_0[0]), .out(far_3_3573_1[0]));    relay_conn far_3_3573_1_b(.in(far_3_3573_0[1]), .out(far_3_3573_1[1]));
    assign layer_3[513] = far_3_3573_1[1]; 
    wire [1:0] far_3_3574_0;    relay_conn far_3_3574_0_a(.in(layer_2[133]), .out(far_3_3574_0[0]));    relay_conn far_3_3574_0_b(.in(layer_2[252]), .out(far_3_3574_0[1]));
    wire [1:0] far_3_3574_1;    relay_conn far_3_3574_1_a(.in(far_3_3574_0[0]), .out(far_3_3574_1[0]));    relay_conn far_3_3574_1_b(.in(far_3_3574_0[1]), .out(far_3_3574_1[1]));
    wire [1:0] far_3_3574_2;    relay_conn far_3_3574_2_a(.in(far_3_3574_1[0]), .out(far_3_3574_2[0]));    relay_conn far_3_3574_2_b(.in(far_3_3574_1[1]), .out(far_3_3574_2[1]));
    assign layer_3[514] = far_3_3574_2[0] & far_3_3574_2[1]; 
    assign layer_3[515] = layer_2[506] ^ layer_2[500]; 
    wire [1:0] far_3_3576_0;    relay_conn far_3_3576_0_a(.in(layer_2[915]), .out(far_3_3576_0[0]));    relay_conn far_3_3576_0_b(.in(layer_2[836]), .out(far_3_3576_0[1]));
    wire [1:0] far_3_3576_1;    relay_conn far_3_3576_1_a(.in(far_3_3576_0[0]), .out(far_3_3576_1[0]));    relay_conn far_3_3576_1_b(.in(far_3_3576_0[1]), .out(far_3_3576_1[1]));
    assign layer_3[516] = ~far_3_3576_1[0]; 
    assign layer_3[517] = ~layer_2[348]; 
    wire [1:0] far_3_3578_0;    relay_conn far_3_3578_0_a(.in(layer_2[1017]), .out(far_3_3578_0[0]));    relay_conn far_3_3578_0_b(.in(layer_2[903]), .out(far_3_3578_0[1]));
    wire [1:0] far_3_3578_1;    relay_conn far_3_3578_1_a(.in(far_3_3578_0[0]), .out(far_3_3578_1[0]));    relay_conn far_3_3578_1_b(.in(far_3_3578_0[1]), .out(far_3_3578_1[1]));
    wire [1:0] far_3_3578_2;    relay_conn far_3_3578_2_a(.in(far_3_3578_1[0]), .out(far_3_3578_2[0]));    relay_conn far_3_3578_2_b(.in(far_3_3578_1[1]), .out(far_3_3578_2[1]));
    assign layer_3[518] = far_3_3578_2[0]; 
    wire [1:0] far_3_3579_0;    relay_conn far_3_3579_0_a(.in(layer_2[550]), .out(far_3_3579_0[0]));    relay_conn far_3_3579_0_b(.in(layer_2[498]), .out(far_3_3579_0[1]));
    assign layer_3[519] = ~(far_3_3579_0[0] | far_3_3579_0[1]); 
    wire [1:0] far_3_3580_0;    relay_conn far_3_3580_0_a(.in(layer_2[335]), .out(far_3_3580_0[0]));    relay_conn far_3_3580_0_b(.in(layer_2[379]), .out(far_3_3580_0[1]));
    assign layer_3[520] = far_3_3580_0[0] & ~far_3_3580_0[1]; 
    assign layer_3[521] = ~(layer_2[995] & layer_2[1013]); 
    wire [1:0] far_3_3582_0;    relay_conn far_3_3582_0_a(.in(layer_2[225]), .out(far_3_3582_0[0]));    relay_conn far_3_3582_0_b(.in(layer_2[310]), .out(far_3_3582_0[1]));
    wire [1:0] far_3_3582_1;    relay_conn far_3_3582_1_a(.in(far_3_3582_0[0]), .out(far_3_3582_1[0]));    relay_conn far_3_3582_1_b(.in(far_3_3582_0[1]), .out(far_3_3582_1[1]));
    assign layer_3[522] = far_3_3582_1[0] & far_3_3582_1[1]; 
    wire [1:0] far_3_3583_0;    relay_conn far_3_3583_0_a(.in(layer_2[248]), .out(far_3_3583_0[0]));    relay_conn far_3_3583_0_b(.in(layer_2[298]), .out(far_3_3583_0[1]));
    assign layer_3[523] = ~(far_3_3583_0[0] & far_3_3583_0[1]); 
    assign layer_3[524] = ~layer_2[203] | (layer_2[203] & layer_2[205]); 
    assign layer_3[525] = ~layer_2[154] | (layer_2[163] & layer_2[154]); 
    wire [1:0] far_3_3586_0;    relay_conn far_3_3586_0_a(.in(layer_2[791]), .out(far_3_3586_0[0]));    relay_conn far_3_3586_0_b(.in(layer_2[916]), .out(far_3_3586_0[1]));
    wire [1:0] far_3_3586_1;    relay_conn far_3_3586_1_a(.in(far_3_3586_0[0]), .out(far_3_3586_1[0]));    relay_conn far_3_3586_1_b(.in(far_3_3586_0[1]), .out(far_3_3586_1[1]));
    wire [1:0] far_3_3586_2;    relay_conn far_3_3586_2_a(.in(far_3_3586_1[0]), .out(far_3_3586_2[0]));    relay_conn far_3_3586_2_b(.in(far_3_3586_1[1]), .out(far_3_3586_2[1]));
    assign layer_3[526] = ~far_3_3586_2[1] | (far_3_3586_2[0] & far_3_3586_2[1]); 
    wire [1:0] far_3_3587_0;    relay_conn far_3_3587_0_a(.in(layer_2[134]), .out(far_3_3587_0[0]));    relay_conn far_3_3587_0_b(.in(layer_2[192]), .out(far_3_3587_0[1]));
    assign layer_3[527] = ~far_3_3587_0[1] | (far_3_3587_0[0] & far_3_3587_0[1]); 
    wire [1:0] far_3_3588_0;    relay_conn far_3_3588_0_a(.in(layer_2[558]), .out(far_3_3588_0[0]));    relay_conn far_3_3588_0_b(.in(layer_2[667]), .out(far_3_3588_0[1]));
    wire [1:0] far_3_3588_1;    relay_conn far_3_3588_1_a(.in(far_3_3588_0[0]), .out(far_3_3588_1[0]));    relay_conn far_3_3588_1_b(.in(far_3_3588_0[1]), .out(far_3_3588_1[1]));
    wire [1:0] far_3_3588_2;    relay_conn far_3_3588_2_a(.in(far_3_3588_1[0]), .out(far_3_3588_2[0]));    relay_conn far_3_3588_2_b(.in(far_3_3588_1[1]), .out(far_3_3588_2[1]));
    assign layer_3[528] = ~(far_3_3588_2[0] ^ far_3_3588_2[1]); 
    wire [1:0] far_3_3589_0;    relay_conn far_3_3589_0_a(.in(layer_2[553]), .out(far_3_3589_0[0]));    relay_conn far_3_3589_0_b(.in(layer_2[610]), .out(far_3_3589_0[1]));
    assign layer_3[529] = ~(far_3_3589_0[0] | far_3_3589_0[1]); 
    assign layer_3[530] = ~(layer_2[292] | layer_2[265]); 
    assign layer_3[531] = ~(layer_2[200] | layer_2[177]); 
    wire [1:0] far_3_3592_0;    relay_conn far_3_3592_0_a(.in(layer_2[882]), .out(far_3_3592_0[0]));    relay_conn far_3_3592_0_b(.in(layer_2[840]), .out(far_3_3592_0[1]));
    assign layer_3[532] = far_3_3592_0[0] & ~far_3_3592_0[1]; 
    wire [1:0] far_3_3593_0;    relay_conn far_3_3593_0_a(.in(layer_2[345]), .out(far_3_3593_0[0]));    relay_conn far_3_3593_0_b(.in(layer_2[235]), .out(far_3_3593_0[1]));
    wire [1:0] far_3_3593_1;    relay_conn far_3_3593_1_a(.in(far_3_3593_0[0]), .out(far_3_3593_1[0]));    relay_conn far_3_3593_1_b(.in(far_3_3593_0[1]), .out(far_3_3593_1[1]));
    wire [1:0] far_3_3593_2;    relay_conn far_3_3593_2_a(.in(far_3_3593_1[0]), .out(far_3_3593_2[0]));    relay_conn far_3_3593_2_b(.in(far_3_3593_1[1]), .out(far_3_3593_2[1]));
    assign layer_3[533] = far_3_3593_2[0] ^ far_3_3593_2[1]; 
    wire [1:0] far_3_3594_0;    relay_conn far_3_3594_0_a(.in(layer_2[995]), .out(far_3_3594_0[0]));    relay_conn far_3_3594_0_b(.in(layer_2[880]), .out(far_3_3594_0[1]));
    wire [1:0] far_3_3594_1;    relay_conn far_3_3594_1_a(.in(far_3_3594_0[0]), .out(far_3_3594_1[0]));    relay_conn far_3_3594_1_b(.in(far_3_3594_0[1]), .out(far_3_3594_1[1]));
    wire [1:0] far_3_3594_2;    relay_conn far_3_3594_2_a(.in(far_3_3594_1[0]), .out(far_3_3594_2[0]));    relay_conn far_3_3594_2_b(.in(far_3_3594_1[1]), .out(far_3_3594_2[1]));
    assign layer_3[534] = ~far_3_3594_2[1] | (far_3_3594_2[0] & far_3_3594_2[1]); 
    wire [1:0] far_3_3595_0;    relay_conn far_3_3595_0_a(.in(layer_2[912]), .out(far_3_3595_0[0]));    relay_conn far_3_3595_0_b(.in(layer_2[785]), .out(far_3_3595_0[1]));
    wire [1:0] far_3_3595_1;    relay_conn far_3_3595_1_a(.in(far_3_3595_0[0]), .out(far_3_3595_1[0]));    relay_conn far_3_3595_1_b(.in(far_3_3595_0[1]), .out(far_3_3595_1[1]));
    wire [1:0] far_3_3595_2;    relay_conn far_3_3595_2_a(.in(far_3_3595_1[0]), .out(far_3_3595_2[0]));    relay_conn far_3_3595_2_b(.in(far_3_3595_1[1]), .out(far_3_3595_2[1]));
    assign layer_3[535] = far_3_3595_2[0] & ~far_3_3595_2[1]; 
    assign layer_3[536] = ~layer_2[920] | (layer_2[949] & layer_2[920]); 
    wire [1:0] far_3_3597_0;    relay_conn far_3_3597_0_a(.in(layer_2[971]), .out(far_3_3597_0[0]));    relay_conn far_3_3597_0_b(.in(layer_2[1016]), .out(far_3_3597_0[1]));
    assign layer_3[537] = far_3_3597_0[1] & ~far_3_3597_0[0]; 
    wire [1:0] far_3_3598_0;    relay_conn far_3_3598_0_a(.in(layer_2[986]), .out(far_3_3598_0[0]));    relay_conn far_3_3598_0_b(.in(layer_2[927]), .out(far_3_3598_0[1]));
    assign layer_3[538] = ~far_3_3598_0[0]; 
    wire [1:0] far_3_3599_0;    relay_conn far_3_3599_0_a(.in(layer_2[748]), .out(far_3_3599_0[0]));    relay_conn far_3_3599_0_b(.in(layer_2[703]), .out(far_3_3599_0[1]));
    assign layer_3[539] = far_3_3599_0[1]; 
    wire [1:0] far_3_3600_0;    relay_conn far_3_3600_0_a(.in(layer_2[1005]), .out(far_3_3600_0[0]));    relay_conn far_3_3600_0_b(.in(layer_2[884]), .out(far_3_3600_0[1]));
    wire [1:0] far_3_3600_1;    relay_conn far_3_3600_1_a(.in(far_3_3600_0[0]), .out(far_3_3600_1[0]));    relay_conn far_3_3600_1_b(.in(far_3_3600_0[1]), .out(far_3_3600_1[1]));
    wire [1:0] far_3_3600_2;    relay_conn far_3_3600_2_a(.in(far_3_3600_1[0]), .out(far_3_3600_2[0]));    relay_conn far_3_3600_2_b(.in(far_3_3600_1[1]), .out(far_3_3600_2[1]));
    assign layer_3[540] = far_3_3600_2[1]; 
    wire [1:0] far_3_3601_0;    relay_conn far_3_3601_0_a(.in(layer_2[949]), .out(far_3_3601_0[0]));    relay_conn far_3_3601_0_b(.in(layer_2[997]), .out(far_3_3601_0[1]));
    assign layer_3[541] = ~far_3_3601_0[0] | (far_3_3601_0[0] & far_3_3601_0[1]); 
    assign layer_3[542] = ~layer_2[64]; 
    wire [1:0] far_3_3603_0;    relay_conn far_3_3603_0_a(.in(layer_2[774]), .out(far_3_3603_0[0]));    relay_conn far_3_3603_0_b(.in(layer_2[680]), .out(far_3_3603_0[1]));
    wire [1:0] far_3_3603_1;    relay_conn far_3_3603_1_a(.in(far_3_3603_0[0]), .out(far_3_3603_1[0]));    relay_conn far_3_3603_1_b(.in(far_3_3603_0[1]), .out(far_3_3603_1[1]));
    assign layer_3[543] = ~far_3_3603_1[0]; 
    wire [1:0] far_3_3604_0;    relay_conn far_3_3604_0_a(.in(layer_2[912]), .out(far_3_3604_0[0]));    relay_conn far_3_3604_0_b(.in(layer_2[859]), .out(far_3_3604_0[1]));
    assign layer_3[544] = ~(far_3_3604_0[0] & far_3_3604_0[1]); 
    assign layer_3[545] = layer_2[735] | layer_2[749]; 
    wire [1:0] far_3_3606_0;    relay_conn far_3_3606_0_a(.in(layer_2[206]), .out(far_3_3606_0[0]));    relay_conn far_3_3606_0_b(.in(layer_2[309]), .out(far_3_3606_0[1]));
    wire [1:0] far_3_3606_1;    relay_conn far_3_3606_1_a(.in(far_3_3606_0[0]), .out(far_3_3606_1[0]));    relay_conn far_3_3606_1_b(.in(far_3_3606_0[1]), .out(far_3_3606_1[1]));
    wire [1:0] far_3_3606_2;    relay_conn far_3_3606_2_a(.in(far_3_3606_1[0]), .out(far_3_3606_2[0]));    relay_conn far_3_3606_2_b(.in(far_3_3606_1[1]), .out(far_3_3606_2[1]));
    assign layer_3[546] = ~far_3_3606_2[1] | (far_3_3606_2[0] & far_3_3606_2[1]); 
    wire [1:0] far_3_3607_0;    relay_conn far_3_3607_0_a(.in(layer_2[340]), .out(far_3_3607_0[0]));    relay_conn far_3_3607_0_b(.in(layer_2[444]), .out(far_3_3607_0[1]));
    wire [1:0] far_3_3607_1;    relay_conn far_3_3607_1_a(.in(far_3_3607_0[0]), .out(far_3_3607_1[0]));    relay_conn far_3_3607_1_b(.in(far_3_3607_0[1]), .out(far_3_3607_1[1]));
    wire [1:0] far_3_3607_2;    relay_conn far_3_3607_2_a(.in(far_3_3607_1[0]), .out(far_3_3607_2[0]));    relay_conn far_3_3607_2_b(.in(far_3_3607_1[1]), .out(far_3_3607_2[1]));
    assign layer_3[547] = far_3_3607_2[0] | far_3_3607_2[1]; 
    wire [1:0] far_3_3608_0;    relay_conn far_3_3608_0_a(.in(layer_2[126]), .out(far_3_3608_0[0]));    relay_conn far_3_3608_0_b(.in(layer_2[6]), .out(far_3_3608_0[1]));
    wire [1:0] far_3_3608_1;    relay_conn far_3_3608_1_a(.in(far_3_3608_0[0]), .out(far_3_3608_1[0]));    relay_conn far_3_3608_1_b(.in(far_3_3608_0[1]), .out(far_3_3608_1[1]));
    wire [1:0] far_3_3608_2;    relay_conn far_3_3608_2_a(.in(far_3_3608_1[0]), .out(far_3_3608_2[0]));    relay_conn far_3_3608_2_b(.in(far_3_3608_1[1]), .out(far_3_3608_2[1]));
    assign layer_3[548] = ~(far_3_3608_2[0] | far_3_3608_2[1]); 
    wire [1:0] far_3_3609_0;    relay_conn far_3_3609_0_a(.in(layer_2[644]), .out(far_3_3609_0[0]));    relay_conn far_3_3609_0_b(.in(layer_2[610]), .out(far_3_3609_0[1]));
    assign layer_3[549] = ~(far_3_3609_0[0] ^ far_3_3609_0[1]); 
    wire [1:0] far_3_3610_0;    relay_conn far_3_3610_0_a(.in(layer_2[1017]), .out(far_3_3610_0[0]));    relay_conn far_3_3610_0_b(.in(layer_2[910]), .out(far_3_3610_0[1]));
    wire [1:0] far_3_3610_1;    relay_conn far_3_3610_1_a(.in(far_3_3610_0[0]), .out(far_3_3610_1[0]));    relay_conn far_3_3610_1_b(.in(far_3_3610_0[1]), .out(far_3_3610_1[1]));
    wire [1:0] far_3_3610_2;    relay_conn far_3_3610_2_a(.in(far_3_3610_1[0]), .out(far_3_3610_2[0]));    relay_conn far_3_3610_2_b(.in(far_3_3610_1[1]), .out(far_3_3610_2[1]));
    assign layer_3[550] = ~(far_3_3610_2[0] | far_3_3610_2[1]); 
    wire [1:0] far_3_3611_0;    relay_conn far_3_3611_0_a(.in(layer_2[681]), .out(far_3_3611_0[0]));    relay_conn far_3_3611_0_b(.in(layer_2[553]), .out(far_3_3611_0[1]));
    wire [1:0] far_3_3611_1;    relay_conn far_3_3611_1_a(.in(far_3_3611_0[0]), .out(far_3_3611_1[0]));    relay_conn far_3_3611_1_b(.in(far_3_3611_0[1]), .out(far_3_3611_1[1]));
    wire [1:0] far_3_3611_2;    relay_conn far_3_3611_2_a(.in(far_3_3611_1[0]), .out(far_3_3611_2[0]));    relay_conn far_3_3611_2_b(.in(far_3_3611_1[1]), .out(far_3_3611_2[1]));
    wire [1:0] far_3_3611_3;    relay_conn far_3_3611_3_a(.in(far_3_3611_2[0]), .out(far_3_3611_3[0]));    relay_conn far_3_3611_3_b(.in(far_3_3611_2[1]), .out(far_3_3611_3[1]));
    assign layer_3[551] = ~(far_3_3611_3[0] ^ far_3_3611_3[1]); 
    wire [1:0] far_3_3612_0;    relay_conn far_3_3612_0_a(.in(layer_2[433]), .out(far_3_3612_0[0]));    relay_conn far_3_3612_0_b(.in(layer_2[307]), .out(far_3_3612_0[1]));
    wire [1:0] far_3_3612_1;    relay_conn far_3_3612_1_a(.in(far_3_3612_0[0]), .out(far_3_3612_1[0]));    relay_conn far_3_3612_1_b(.in(far_3_3612_0[1]), .out(far_3_3612_1[1]));
    wire [1:0] far_3_3612_2;    relay_conn far_3_3612_2_a(.in(far_3_3612_1[0]), .out(far_3_3612_2[0]));    relay_conn far_3_3612_2_b(.in(far_3_3612_1[1]), .out(far_3_3612_2[1]));
    assign layer_3[552] = far_3_3612_2[0] | far_3_3612_2[1]; 
    wire [1:0] far_3_3613_0;    relay_conn far_3_3613_0_a(.in(layer_2[781]), .out(far_3_3613_0[0]));    relay_conn far_3_3613_0_b(.in(layer_2[822]), .out(far_3_3613_0[1]));
    assign layer_3[553] = ~(far_3_3613_0[0] ^ far_3_3613_0[1]); 
    wire [1:0] far_3_3614_0;    relay_conn far_3_3614_0_a(.in(layer_2[29]), .out(far_3_3614_0[0]));    relay_conn far_3_3614_0_b(.in(layer_2[61]), .out(far_3_3614_0[1]));
    assign layer_3[554] = ~far_3_3614_0[1]; 
    assign layer_3[555] = layer_2[341]; 
    wire [1:0] far_3_3616_0;    relay_conn far_3_3616_0_a(.in(layer_2[396]), .out(far_3_3616_0[0]));    relay_conn far_3_3616_0_b(.in(layer_2[340]), .out(far_3_3616_0[1]));
    assign layer_3[556] = ~far_3_3616_0[1]; 
    wire [1:0] far_3_3617_0;    relay_conn far_3_3617_0_a(.in(layer_2[265]), .out(far_3_3617_0[0]));    relay_conn far_3_3617_0_b(.in(layer_2[194]), .out(far_3_3617_0[1]));
    wire [1:0] far_3_3617_1;    relay_conn far_3_3617_1_a(.in(far_3_3617_0[0]), .out(far_3_3617_1[0]));    relay_conn far_3_3617_1_b(.in(far_3_3617_0[1]), .out(far_3_3617_1[1]));
    assign layer_3[557] = ~far_3_3617_1[1]; 
    wire [1:0] far_3_3618_0;    relay_conn far_3_3618_0_a(.in(layer_2[222]), .out(far_3_3618_0[0]));    relay_conn far_3_3618_0_b(.in(layer_2[120]), .out(far_3_3618_0[1]));
    wire [1:0] far_3_3618_1;    relay_conn far_3_3618_1_a(.in(far_3_3618_0[0]), .out(far_3_3618_1[0]));    relay_conn far_3_3618_1_b(.in(far_3_3618_0[1]), .out(far_3_3618_1[1]));
    wire [1:0] far_3_3618_2;    relay_conn far_3_3618_2_a(.in(far_3_3618_1[0]), .out(far_3_3618_2[0]));    relay_conn far_3_3618_2_b(.in(far_3_3618_1[1]), .out(far_3_3618_2[1]));
    assign layer_3[558] = far_3_3618_2[0] & ~far_3_3618_2[1]; 
    assign layer_3[559] = ~layer_2[521] | (layer_2[543] & layer_2[521]); 
    assign layer_3[560] = layer_2[172] ^ layer_2[183]; 
    assign layer_3[561] = ~(layer_2[252] & layer_2[244]); 
    wire [1:0] far_3_3622_0;    relay_conn far_3_3622_0_a(.in(layer_2[324]), .out(far_3_3622_0[0]));    relay_conn far_3_3622_0_b(.in(layer_2[262]), .out(far_3_3622_0[1]));
    assign layer_3[562] = far_3_3622_0[0] & far_3_3622_0[1]; 
    wire [1:0] far_3_3623_0;    relay_conn far_3_3623_0_a(.in(layer_2[87]), .out(far_3_3623_0[0]));    relay_conn far_3_3623_0_b(.in(layer_2[190]), .out(far_3_3623_0[1]));
    wire [1:0] far_3_3623_1;    relay_conn far_3_3623_1_a(.in(far_3_3623_0[0]), .out(far_3_3623_1[0]));    relay_conn far_3_3623_1_b(.in(far_3_3623_0[1]), .out(far_3_3623_1[1]));
    wire [1:0] far_3_3623_2;    relay_conn far_3_3623_2_a(.in(far_3_3623_1[0]), .out(far_3_3623_2[0]));    relay_conn far_3_3623_2_b(.in(far_3_3623_1[1]), .out(far_3_3623_2[1]));
    assign layer_3[563] = ~far_3_3623_2[0] | (far_3_3623_2[0] & far_3_3623_2[1]); 
    assign layer_3[564] = layer_2[877] & ~layer_2[852]; 
    wire [1:0] far_3_3625_0;    relay_conn far_3_3625_0_a(.in(layer_2[129]), .out(far_3_3625_0[0]));    relay_conn far_3_3625_0_b(.in(layer_2[200]), .out(far_3_3625_0[1]));
    wire [1:0] far_3_3625_1;    relay_conn far_3_3625_1_a(.in(far_3_3625_0[0]), .out(far_3_3625_1[0]));    relay_conn far_3_3625_1_b(.in(far_3_3625_0[1]), .out(far_3_3625_1[1]));
    assign layer_3[565] = ~(far_3_3625_1[0] | far_3_3625_1[1]); 
    wire [1:0] far_3_3626_0;    relay_conn far_3_3626_0_a(.in(layer_2[132]), .out(far_3_3626_0[0]));    relay_conn far_3_3626_0_b(.in(layer_2[28]), .out(far_3_3626_0[1]));
    wire [1:0] far_3_3626_1;    relay_conn far_3_3626_1_a(.in(far_3_3626_0[0]), .out(far_3_3626_1[0]));    relay_conn far_3_3626_1_b(.in(far_3_3626_0[1]), .out(far_3_3626_1[1]));
    wire [1:0] far_3_3626_2;    relay_conn far_3_3626_2_a(.in(far_3_3626_1[0]), .out(far_3_3626_2[0]));    relay_conn far_3_3626_2_b(.in(far_3_3626_1[1]), .out(far_3_3626_2[1]));
    assign layer_3[566] = far_3_3626_2[0] & far_3_3626_2[1]; 
    wire [1:0] far_3_3627_0;    relay_conn far_3_3627_0_a(.in(layer_2[855]), .out(far_3_3627_0[0]));    relay_conn far_3_3627_0_b(.in(layer_2[748]), .out(far_3_3627_0[1]));
    wire [1:0] far_3_3627_1;    relay_conn far_3_3627_1_a(.in(far_3_3627_0[0]), .out(far_3_3627_1[0]));    relay_conn far_3_3627_1_b(.in(far_3_3627_0[1]), .out(far_3_3627_1[1]));
    wire [1:0] far_3_3627_2;    relay_conn far_3_3627_2_a(.in(far_3_3627_1[0]), .out(far_3_3627_2[0]));    relay_conn far_3_3627_2_b(.in(far_3_3627_1[1]), .out(far_3_3627_2[1]));
    assign layer_3[567] = ~(far_3_3627_2[0] & far_3_3627_2[1]); 
    wire [1:0] far_3_3628_0;    relay_conn far_3_3628_0_a(.in(layer_2[603]), .out(far_3_3628_0[0]));    relay_conn far_3_3628_0_b(.in(layer_2[509]), .out(far_3_3628_0[1]));
    wire [1:0] far_3_3628_1;    relay_conn far_3_3628_1_a(.in(far_3_3628_0[0]), .out(far_3_3628_1[0]));    relay_conn far_3_3628_1_b(.in(far_3_3628_0[1]), .out(far_3_3628_1[1]));
    assign layer_3[568] = ~(far_3_3628_1[0] & far_3_3628_1[1]); 
    wire [1:0] far_3_3629_0;    relay_conn far_3_3629_0_a(.in(layer_2[244]), .out(far_3_3629_0[0]));    relay_conn far_3_3629_0_b(.in(layer_2[185]), .out(far_3_3629_0[1]));
    assign layer_3[569] = ~far_3_3629_0[0]; 
    wire [1:0] far_3_3630_0;    relay_conn far_3_3630_0_a(.in(layer_2[730]), .out(far_3_3630_0[0]));    relay_conn far_3_3630_0_b(.in(layer_2[855]), .out(far_3_3630_0[1]));
    wire [1:0] far_3_3630_1;    relay_conn far_3_3630_1_a(.in(far_3_3630_0[0]), .out(far_3_3630_1[0]));    relay_conn far_3_3630_1_b(.in(far_3_3630_0[1]), .out(far_3_3630_1[1]));
    wire [1:0] far_3_3630_2;    relay_conn far_3_3630_2_a(.in(far_3_3630_1[0]), .out(far_3_3630_2[0]));    relay_conn far_3_3630_2_b(.in(far_3_3630_1[1]), .out(far_3_3630_2[1]));
    assign layer_3[570] = ~far_3_3630_2[1]; 
    wire [1:0] far_3_3631_0;    relay_conn far_3_3631_0_a(.in(layer_2[299]), .out(far_3_3631_0[0]));    relay_conn far_3_3631_0_b(.in(layer_2[379]), .out(far_3_3631_0[1]));
    wire [1:0] far_3_3631_1;    relay_conn far_3_3631_1_a(.in(far_3_3631_0[0]), .out(far_3_3631_1[0]));    relay_conn far_3_3631_1_b(.in(far_3_3631_0[1]), .out(far_3_3631_1[1]));
    assign layer_3[571] = far_3_3631_1[0] & ~far_3_3631_1[1]; 
    wire [1:0] far_3_3632_0;    relay_conn far_3_3632_0_a(.in(layer_2[465]), .out(far_3_3632_0[0]));    relay_conn far_3_3632_0_b(.in(layer_2[383]), .out(far_3_3632_0[1]));
    wire [1:0] far_3_3632_1;    relay_conn far_3_3632_1_a(.in(far_3_3632_0[0]), .out(far_3_3632_1[0]));    relay_conn far_3_3632_1_b(.in(far_3_3632_0[1]), .out(far_3_3632_1[1]));
    assign layer_3[572] = far_3_3632_1[1]; 
    assign layer_3[573] = ~layer_2[670] | (layer_2[670] & layer_2[681]); 
    wire [1:0] far_3_3634_0;    relay_conn far_3_3634_0_a(.in(layer_2[652]), .out(far_3_3634_0[0]));    relay_conn far_3_3634_0_b(.in(layer_2[576]), .out(far_3_3634_0[1]));
    wire [1:0] far_3_3634_1;    relay_conn far_3_3634_1_a(.in(far_3_3634_0[0]), .out(far_3_3634_1[0]));    relay_conn far_3_3634_1_b(.in(far_3_3634_0[1]), .out(far_3_3634_1[1]));
    assign layer_3[574] = far_3_3634_1[1]; 
    wire [1:0] far_3_3635_0;    relay_conn far_3_3635_0_a(.in(layer_2[185]), .out(far_3_3635_0[0]));    relay_conn far_3_3635_0_b(.in(layer_2[139]), .out(far_3_3635_0[1]));
    assign layer_3[575] = far_3_3635_0[0] & ~far_3_3635_0[1]; 
    wire [1:0] far_3_3636_0;    relay_conn far_3_3636_0_a(.in(layer_2[827]), .out(far_3_3636_0[0]));    relay_conn far_3_3636_0_b(.in(layer_2[726]), .out(far_3_3636_0[1]));
    wire [1:0] far_3_3636_1;    relay_conn far_3_3636_1_a(.in(far_3_3636_0[0]), .out(far_3_3636_1[0]));    relay_conn far_3_3636_1_b(.in(far_3_3636_0[1]), .out(far_3_3636_1[1]));
    wire [1:0] far_3_3636_2;    relay_conn far_3_3636_2_a(.in(far_3_3636_1[0]), .out(far_3_3636_2[0]));    relay_conn far_3_3636_2_b(.in(far_3_3636_1[1]), .out(far_3_3636_2[1]));
    assign layer_3[576] = far_3_3636_2[0] & ~far_3_3636_2[1]; 
    wire [1:0] far_3_3637_0;    relay_conn far_3_3637_0_a(.in(layer_2[771]), .out(far_3_3637_0[0]));    relay_conn far_3_3637_0_b(.in(layer_2[646]), .out(far_3_3637_0[1]));
    wire [1:0] far_3_3637_1;    relay_conn far_3_3637_1_a(.in(far_3_3637_0[0]), .out(far_3_3637_1[0]));    relay_conn far_3_3637_1_b(.in(far_3_3637_0[1]), .out(far_3_3637_1[1]));
    wire [1:0] far_3_3637_2;    relay_conn far_3_3637_2_a(.in(far_3_3637_1[0]), .out(far_3_3637_2[0]));    relay_conn far_3_3637_2_b(.in(far_3_3637_1[1]), .out(far_3_3637_2[1]));
    assign layer_3[577] = ~far_3_3637_2[1] | (far_3_3637_2[0] & far_3_3637_2[1]); 
    assign layer_3[578] = layer_2[830] | layer_2[836]; 
    wire [1:0] far_3_3639_0;    relay_conn far_3_3639_0_a(.in(layer_2[836]), .out(far_3_3639_0[0]));    relay_conn far_3_3639_0_b(.in(layer_2[899]), .out(far_3_3639_0[1]));
    assign layer_3[579] = ~far_3_3639_0[1] | (far_3_3639_0[0] & far_3_3639_0[1]); 
    assign layer_3[580] = ~layer_2[381]; 
    wire [1:0] far_3_3641_0;    relay_conn far_3_3641_0_a(.in(layer_2[517]), .out(far_3_3641_0[0]));    relay_conn far_3_3641_0_b(.in(layer_2[565]), .out(far_3_3641_0[1]));
    assign layer_3[581] = ~(far_3_3641_0[0] ^ far_3_3641_0[1]); 
    assign layer_3[582] = layer_2[807]; 
    wire [1:0] far_3_3643_0;    relay_conn far_3_3643_0_a(.in(layer_2[23]), .out(far_3_3643_0[0]));    relay_conn far_3_3643_0_b(.in(layer_2[138]), .out(far_3_3643_0[1]));
    wire [1:0] far_3_3643_1;    relay_conn far_3_3643_1_a(.in(far_3_3643_0[0]), .out(far_3_3643_1[0]));    relay_conn far_3_3643_1_b(.in(far_3_3643_0[1]), .out(far_3_3643_1[1]));
    wire [1:0] far_3_3643_2;    relay_conn far_3_3643_2_a(.in(far_3_3643_1[0]), .out(far_3_3643_2[0]));    relay_conn far_3_3643_2_b(.in(far_3_3643_1[1]), .out(far_3_3643_2[1]));
    assign layer_3[583] = ~(far_3_3643_2[0] & far_3_3643_2[1]); 
    wire [1:0] far_3_3644_0;    relay_conn far_3_3644_0_a(.in(layer_2[762]), .out(far_3_3644_0[0]));    relay_conn far_3_3644_0_b(.in(layer_2[709]), .out(far_3_3644_0[1]));
    assign layer_3[584] = far_3_3644_0[1]; 
    wire [1:0] far_3_3645_0;    relay_conn far_3_3645_0_a(.in(layer_2[209]), .out(far_3_3645_0[0]));    relay_conn far_3_3645_0_b(.in(layer_2[120]), .out(far_3_3645_0[1]));
    wire [1:0] far_3_3645_1;    relay_conn far_3_3645_1_a(.in(far_3_3645_0[0]), .out(far_3_3645_1[0]));    relay_conn far_3_3645_1_b(.in(far_3_3645_0[1]), .out(far_3_3645_1[1]));
    assign layer_3[585] = far_3_3645_1[1] & ~far_3_3645_1[0]; 
    wire [1:0] far_3_3646_0;    relay_conn far_3_3646_0_a(.in(layer_2[928]), .out(far_3_3646_0[0]));    relay_conn far_3_3646_0_b(.in(layer_2[835]), .out(far_3_3646_0[1]));
    wire [1:0] far_3_3646_1;    relay_conn far_3_3646_1_a(.in(far_3_3646_0[0]), .out(far_3_3646_1[0]));    relay_conn far_3_3646_1_b(.in(far_3_3646_0[1]), .out(far_3_3646_1[1]));
    assign layer_3[586] = ~far_3_3646_1[1]; 
    wire [1:0] far_3_3647_0;    relay_conn far_3_3647_0_a(.in(layer_2[969]), .out(far_3_3647_0[0]));    relay_conn far_3_3647_0_b(.in(layer_2[856]), .out(far_3_3647_0[1]));
    wire [1:0] far_3_3647_1;    relay_conn far_3_3647_1_a(.in(far_3_3647_0[0]), .out(far_3_3647_1[0]));    relay_conn far_3_3647_1_b(.in(far_3_3647_0[1]), .out(far_3_3647_1[1]));
    wire [1:0] far_3_3647_2;    relay_conn far_3_3647_2_a(.in(far_3_3647_1[0]), .out(far_3_3647_2[0]));    relay_conn far_3_3647_2_b(.in(far_3_3647_1[1]), .out(far_3_3647_2[1]));
    assign layer_3[587] = far_3_3647_2[0] & ~far_3_3647_2[1]; 
    wire [1:0] far_3_3648_0;    relay_conn far_3_3648_0_a(.in(layer_2[604]), .out(far_3_3648_0[0]));    relay_conn far_3_3648_0_b(.in(layer_2[714]), .out(far_3_3648_0[1]));
    wire [1:0] far_3_3648_1;    relay_conn far_3_3648_1_a(.in(far_3_3648_0[0]), .out(far_3_3648_1[0]));    relay_conn far_3_3648_1_b(.in(far_3_3648_0[1]), .out(far_3_3648_1[1]));
    wire [1:0] far_3_3648_2;    relay_conn far_3_3648_2_a(.in(far_3_3648_1[0]), .out(far_3_3648_2[0]));    relay_conn far_3_3648_2_b(.in(far_3_3648_1[1]), .out(far_3_3648_2[1]));
    assign layer_3[588] = ~far_3_3648_2[1] | (far_3_3648_2[0] & far_3_3648_2[1]); 
    wire [1:0] far_3_3649_0;    relay_conn far_3_3649_0_a(.in(layer_2[460]), .out(far_3_3649_0[0]));    relay_conn far_3_3649_0_b(.in(layer_2[509]), .out(far_3_3649_0[1]));
    assign layer_3[589] = far_3_3649_0[0] & far_3_3649_0[1]; 
    assign layer_3[590] = ~layer_2[738] | (layer_2[758] & layer_2[738]); 
    wire [1:0] far_3_3651_0;    relay_conn far_3_3651_0_a(.in(layer_2[950]), .out(far_3_3651_0[0]));    relay_conn far_3_3651_0_b(.in(layer_2[880]), .out(far_3_3651_0[1]));
    wire [1:0] far_3_3651_1;    relay_conn far_3_3651_1_a(.in(far_3_3651_0[0]), .out(far_3_3651_1[0]));    relay_conn far_3_3651_1_b(.in(far_3_3651_0[1]), .out(far_3_3651_1[1]));
    assign layer_3[591] = ~far_3_3651_1[0] | (far_3_3651_1[0] & far_3_3651_1[1]); 
    wire [1:0] far_3_3652_0;    relay_conn far_3_3652_0_a(.in(layer_2[685]), .out(far_3_3652_0[0]));    relay_conn far_3_3652_0_b(.in(layer_2[560]), .out(far_3_3652_0[1]));
    wire [1:0] far_3_3652_1;    relay_conn far_3_3652_1_a(.in(far_3_3652_0[0]), .out(far_3_3652_1[0]));    relay_conn far_3_3652_1_b(.in(far_3_3652_0[1]), .out(far_3_3652_1[1]));
    wire [1:0] far_3_3652_2;    relay_conn far_3_3652_2_a(.in(far_3_3652_1[0]), .out(far_3_3652_2[0]));    relay_conn far_3_3652_2_b(.in(far_3_3652_1[1]), .out(far_3_3652_2[1]));
    assign layer_3[592] = ~(far_3_3652_2[0] | far_3_3652_2[1]); 
    wire [1:0] far_3_3653_0;    relay_conn far_3_3653_0_a(.in(layer_2[452]), .out(far_3_3653_0[0]));    relay_conn far_3_3653_0_b(.in(layer_2[336]), .out(far_3_3653_0[1]));
    wire [1:0] far_3_3653_1;    relay_conn far_3_3653_1_a(.in(far_3_3653_0[0]), .out(far_3_3653_1[0]));    relay_conn far_3_3653_1_b(.in(far_3_3653_0[1]), .out(far_3_3653_1[1]));
    wire [1:0] far_3_3653_2;    relay_conn far_3_3653_2_a(.in(far_3_3653_1[0]), .out(far_3_3653_2[0]));    relay_conn far_3_3653_2_b(.in(far_3_3653_1[1]), .out(far_3_3653_2[1]));
    assign layer_3[593] = far_3_3653_2[0] | far_3_3653_2[1]; 
    assign layer_3[594] = layer_2[958] & ~layer_2[927]; 
    wire [1:0] far_3_3655_0;    relay_conn far_3_3655_0_a(.in(layer_2[830]), .out(far_3_3655_0[0]));    relay_conn far_3_3655_0_b(.in(layer_2[748]), .out(far_3_3655_0[1]));
    wire [1:0] far_3_3655_1;    relay_conn far_3_3655_1_a(.in(far_3_3655_0[0]), .out(far_3_3655_1[0]));    relay_conn far_3_3655_1_b(.in(far_3_3655_0[1]), .out(far_3_3655_1[1]));
    assign layer_3[595] = far_3_3655_1[0] & far_3_3655_1[1]; 
    wire [1:0] far_3_3656_0;    relay_conn far_3_3656_0_a(.in(layer_2[79]), .out(far_3_3656_0[0]));    relay_conn far_3_3656_0_b(.in(layer_2[151]), .out(far_3_3656_0[1]));
    wire [1:0] far_3_3656_1;    relay_conn far_3_3656_1_a(.in(far_3_3656_0[0]), .out(far_3_3656_1[0]));    relay_conn far_3_3656_1_b(.in(far_3_3656_0[1]), .out(far_3_3656_1[1]));
    assign layer_3[596] = far_3_3656_1[0] | far_3_3656_1[1]; 
    wire [1:0] far_3_3657_0;    relay_conn far_3_3657_0_a(.in(layer_2[379]), .out(far_3_3657_0[0]));    relay_conn far_3_3657_0_b(.in(layer_2[253]), .out(far_3_3657_0[1]));
    wire [1:0] far_3_3657_1;    relay_conn far_3_3657_1_a(.in(far_3_3657_0[0]), .out(far_3_3657_1[0]));    relay_conn far_3_3657_1_b(.in(far_3_3657_0[1]), .out(far_3_3657_1[1]));
    wire [1:0] far_3_3657_2;    relay_conn far_3_3657_2_a(.in(far_3_3657_1[0]), .out(far_3_3657_2[0]));    relay_conn far_3_3657_2_b(.in(far_3_3657_1[1]), .out(far_3_3657_2[1]));
    assign layer_3[597] = ~(far_3_3657_2[0] ^ far_3_3657_2[1]); 
    wire [1:0] far_3_3658_0;    relay_conn far_3_3658_0_a(.in(layer_2[892]), .out(far_3_3658_0[0]));    relay_conn far_3_3658_0_b(.in(layer_2[830]), .out(far_3_3658_0[1]));
    assign layer_3[598] = far_3_3658_0[0] & far_3_3658_0[1]; 
    wire [1:0] far_3_3659_0;    relay_conn far_3_3659_0_a(.in(layer_2[102]), .out(far_3_3659_0[0]));    relay_conn far_3_3659_0_b(.in(layer_2[43]), .out(far_3_3659_0[1]));
    assign layer_3[599] = far_3_3659_0[0] & ~far_3_3659_0[1]; 
    wire [1:0] far_3_3660_0;    relay_conn far_3_3660_0_a(.in(layer_2[757]), .out(far_3_3660_0[0]));    relay_conn far_3_3660_0_b(.in(layer_2[866]), .out(far_3_3660_0[1]));
    wire [1:0] far_3_3660_1;    relay_conn far_3_3660_1_a(.in(far_3_3660_0[0]), .out(far_3_3660_1[0]));    relay_conn far_3_3660_1_b(.in(far_3_3660_0[1]), .out(far_3_3660_1[1]));
    wire [1:0] far_3_3660_2;    relay_conn far_3_3660_2_a(.in(far_3_3660_1[0]), .out(far_3_3660_2[0]));    relay_conn far_3_3660_2_b(.in(far_3_3660_1[1]), .out(far_3_3660_2[1]));
    assign layer_3[600] = far_3_3660_2[0] | far_3_3660_2[1]; 
    assign layer_3[601] = ~layer_2[245] | (layer_2[245] & layer_2[260]); 
    wire [1:0] far_3_3662_0;    relay_conn far_3_3662_0_a(.in(layer_2[525]), .out(far_3_3662_0[0]));    relay_conn far_3_3662_0_b(.in(layer_2[411]), .out(far_3_3662_0[1]));
    wire [1:0] far_3_3662_1;    relay_conn far_3_3662_1_a(.in(far_3_3662_0[0]), .out(far_3_3662_1[0]));    relay_conn far_3_3662_1_b(.in(far_3_3662_0[1]), .out(far_3_3662_1[1]));
    wire [1:0] far_3_3662_2;    relay_conn far_3_3662_2_a(.in(far_3_3662_1[0]), .out(far_3_3662_2[0]));    relay_conn far_3_3662_2_b(.in(far_3_3662_1[1]), .out(far_3_3662_2[1]));
    assign layer_3[602] = ~(far_3_3662_2[0] & far_3_3662_2[1]); 
    assign layer_3[603] = layer_2[556] | layer_2[565]; 
    wire [1:0] far_3_3664_0;    relay_conn far_3_3664_0_a(.in(layer_2[803]), .out(far_3_3664_0[0]));    relay_conn far_3_3664_0_b(.in(layer_2[915]), .out(far_3_3664_0[1]));
    wire [1:0] far_3_3664_1;    relay_conn far_3_3664_1_a(.in(far_3_3664_0[0]), .out(far_3_3664_1[0]));    relay_conn far_3_3664_1_b(.in(far_3_3664_0[1]), .out(far_3_3664_1[1]));
    wire [1:0] far_3_3664_2;    relay_conn far_3_3664_2_a(.in(far_3_3664_1[0]), .out(far_3_3664_2[0]));    relay_conn far_3_3664_2_b(.in(far_3_3664_1[1]), .out(far_3_3664_2[1]));
    assign layer_3[604] = ~far_3_3664_2[1]; 
    wire [1:0] far_3_3665_0;    relay_conn far_3_3665_0_a(.in(layer_2[998]), .out(far_3_3665_0[0]));    relay_conn far_3_3665_0_b(.in(layer_2[915]), .out(far_3_3665_0[1]));
    wire [1:0] far_3_3665_1;    relay_conn far_3_3665_1_a(.in(far_3_3665_0[0]), .out(far_3_3665_1[0]));    relay_conn far_3_3665_1_b(.in(far_3_3665_0[1]), .out(far_3_3665_1[1]));
    assign layer_3[605] = far_3_3665_1[1]; 
    assign layer_3[606] = layer_2[233]; 
    wire [1:0] far_3_3667_0;    relay_conn far_3_3667_0_a(.in(layer_2[379]), .out(far_3_3667_0[0]));    relay_conn far_3_3667_0_b(.in(layer_2[313]), .out(far_3_3667_0[1]));
    wire [1:0] far_3_3667_1;    relay_conn far_3_3667_1_a(.in(far_3_3667_0[0]), .out(far_3_3667_1[0]));    relay_conn far_3_3667_1_b(.in(far_3_3667_0[1]), .out(far_3_3667_1[1]));
    assign layer_3[607] = far_3_3667_1[1] & ~far_3_3667_1[0]; 
    wire [1:0] far_3_3668_0;    relay_conn far_3_3668_0_a(.in(layer_2[620]), .out(far_3_3668_0[0]));    relay_conn far_3_3668_0_b(.in(layer_2[688]), .out(far_3_3668_0[1]));
    wire [1:0] far_3_3668_1;    relay_conn far_3_3668_1_a(.in(far_3_3668_0[0]), .out(far_3_3668_1[0]));    relay_conn far_3_3668_1_b(.in(far_3_3668_0[1]), .out(far_3_3668_1[1]));
    assign layer_3[608] = far_3_3668_1[0] ^ far_3_3668_1[1]; 
    assign layer_3[609] = ~layer_2[803]; 
    wire [1:0] far_3_3670_0;    relay_conn far_3_3670_0_a(.in(layer_2[129]), .out(far_3_3670_0[0]));    relay_conn far_3_3670_0_b(.in(layer_2[85]), .out(far_3_3670_0[1]));
    assign layer_3[610] = far_3_3670_0[1]; 
    assign layer_3[611] = ~layer_2[415] | (layer_2[400] & layer_2[415]); 
    wire [1:0] far_3_3672_0;    relay_conn far_3_3672_0_a(.in(layer_2[835]), .out(far_3_3672_0[0]));    relay_conn far_3_3672_0_b(.in(layer_2[715]), .out(far_3_3672_0[1]));
    wire [1:0] far_3_3672_1;    relay_conn far_3_3672_1_a(.in(far_3_3672_0[0]), .out(far_3_3672_1[0]));    relay_conn far_3_3672_1_b(.in(far_3_3672_0[1]), .out(far_3_3672_1[1]));
    wire [1:0] far_3_3672_2;    relay_conn far_3_3672_2_a(.in(far_3_3672_1[0]), .out(far_3_3672_2[0]));    relay_conn far_3_3672_2_b(.in(far_3_3672_1[1]), .out(far_3_3672_2[1]));
    assign layer_3[612] = ~(far_3_3672_2[0] & far_3_3672_2[1]); 
    wire [1:0] far_3_3673_0;    relay_conn far_3_3673_0_a(.in(layer_2[956]), .out(far_3_3673_0[0]));    relay_conn far_3_3673_0_b(.in(layer_2[910]), .out(far_3_3673_0[1]));
    assign layer_3[613] = far_3_3673_0[1] & ~far_3_3673_0[0]; 
    assign layer_3[614] = ~(layer_2[881] & layer_2[912]); 
    wire [1:0] far_3_3675_0;    relay_conn far_3_3675_0_a(.in(layer_2[603]), .out(far_3_3675_0[0]));    relay_conn far_3_3675_0_b(.in(layer_2[524]), .out(far_3_3675_0[1]));
    wire [1:0] far_3_3675_1;    relay_conn far_3_3675_1_a(.in(far_3_3675_0[0]), .out(far_3_3675_1[0]));    relay_conn far_3_3675_1_b(.in(far_3_3675_0[1]), .out(far_3_3675_1[1]));
    assign layer_3[615] = ~(far_3_3675_1[0] & far_3_3675_1[1]); 
    assign layer_3[616] = ~(layer_2[737] | layer_2[716]); 
    wire [1:0] far_3_3677_0;    relay_conn far_3_3677_0_a(.in(layer_2[195]), .out(far_3_3677_0[0]));    relay_conn far_3_3677_0_b(.in(layer_2[309]), .out(far_3_3677_0[1]));
    wire [1:0] far_3_3677_1;    relay_conn far_3_3677_1_a(.in(far_3_3677_0[0]), .out(far_3_3677_1[0]));    relay_conn far_3_3677_1_b(.in(far_3_3677_0[1]), .out(far_3_3677_1[1]));
    wire [1:0] far_3_3677_2;    relay_conn far_3_3677_2_a(.in(far_3_3677_1[0]), .out(far_3_3677_2[0]));    relay_conn far_3_3677_2_b(.in(far_3_3677_1[1]), .out(far_3_3677_2[1]));
    assign layer_3[617] = ~far_3_3677_2[1]; 
    wire [1:0] far_3_3678_0;    relay_conn far_3_3678_0_a(.in(layer_2[757]), .out(far_3_3678_0[0]));    relay_conn far_3_3678_0_b(.in(layer_2[845]), .out(far_3_3678_0[1]));
    wire [1:0] far_3_3678_1;    relay_conn far_3_3678_1_a(.in(far_3_3678_0[0]), .out(far_3_3678_1[0]));    relay_conn far_3_3678_1_b(.in(far_3_3678_0[1]), .out(far_3_3678_1[1]));
    assign layer_3[618] = ~far_3_3678_1[1] | (far_3_3678_1[0] & far_3_3678_1[1]); 
    wire [1:0] far_3_3679_0;    relay_conn far_3_3679_0_a(.in(layer_2[726]), .out(far_3_3679_0[0]));    relay_conn far_3_3679_0_b(.in(layer_2[836]), .out(far_3_3679_0[1]));
    wire [1:0] far_3_3679_1;    relay_conn far_3_3679_1_a(.in(far_3_3679_0[0]), .out(far_3_3679_1[0]));    relay_conn far_3_3679_1_b(.in(far_3_3679_0[1]), .out(far_3_3679_1[1]));
    wire [1:0] far_3_3679_2;    relay_conn far_3_3679_2_a(.in(far_3_3679_1[0]), .out(far_3_3679_2[0]));    relay_conn far_3_3679_2_b(.in(far_3_3679_1[1]), .out(far_3_3679_2[1]));
    assign layer_3[619] = far_3_3679_2[0] | far_3_3679_2[1]; 
    wire [1:0] far_3_3680_0;    relay_conn far_3_3680_0_a(.in(layer_2[341]), .out(far_3_3680_0[0]));    relay_conn far_3_3680_0_b(.in(layer_2[248]), .out(far_3_3680_0[1]));
    wire [1:0] far_3_3680_1;    relay_conn far_3_3680_1_a(.in(far_3_3680_0[0]), .out(far_3_3680_1[0]));    relay_conn far_3_3680_1_b(.in(far_3_3680_0[1]), .out(far_3_3680_1[1]));
    assign layer_3[620] = ~far_3_3680_1[1]; 
    wire [1:0] far_3_3681_0;    relay_conn far_3_3681_0_a(.in(layer_2[75]), .out(far_3_3681_0[0]));    relay_conn far_3_3681_0_b(.in(layer_2[2]), .out(far_3_3681_0[1]));
    wire [1:0] far_3_3681_1;    relay_conn far_3_3681_1_a(.in(far_3_3681_0[0]), .out(far_3_3681_1[0]));    relay_conn far_3_3681_1_b(.in(far_3_3681_0[1]), .out(far_3_3681_1[1]));
    assign layer_3[621] = ~(far_3_3681_1[0] ^ far_3_3681_1[1]); 
    wire [1:0] far_3_3682_0;    relay_conn far_3_3682_0_a(.in(layer_2[910]), .out(far_3_3682_0[0]));    relay_conn far_3_3682_0_b(.in(layer_2[977]), .out(far_3_3682_0[1]));
    wire [1:0] far_3_3682_1;    relay_conn far_3_3682_1_a(.in(far_3_3682_0[0]), .out(far_3_3682_1[0]));    relay_conn far_3_3682_1_b(.in(far_3_3682_0[1]), .out(far_3_3682_1[1]));
    assign layer_3[622] = far_3_3682_1[0] & ~far_3_3682_1[1]; 
    wire [1:0] far_3_3683_0;    relay_conn far_3_3683_0_a(.in(layer_2[41]), .out(far_3_3683_0[0]));    relay_conn far_3_3683_0_b(.in(layer_2[85]), .out(far_3_3683_0[1]));
    assign layer_3[623] = far_3_3683_0[0] & far_3_3683_0[1]; 
    assign layer_3[624] = layer_2[707]; 
    wire [1:0] far_3_3685_0;    relay_conn far_3_3685_0_a(.in(layer_2[341]), .out(far_3_3685_0[0]));    relay_conn far_3_3685_0_b(.in(layer_2[428]), .out(far_3_3685_0[1]));
    wire [1:0] far_3_3685_1;    relay_conn far_3_3685_1_a(.in(far_3_3685_0[0]), .out(far_3_3685_1[0]));    relay_conn far_3_3685_1_b(.in(far_3_3685_0[1]), .out(far_3_3685_1[1]));
    assign layer_3[625] = far_3_3685_1[0] & ~far_3_3685_1[1]; 
    wire [1:0] far_3_3686_0;    relay_conn far_3_3686_0_a(.in(layer_2[330]), .out(far_3_3686_0[0]));    relay_conn far_3_3686_0_b(.in(layer_2[376]), .out(far_3_3686_0[1]));
    assign layer_3[626] = far_3_3686_0[0] | far_3_3686_0[1]; 
    assign layer_3[627] = ~layer_2[348] | (layer_2[336] & layer_2[348]); 
    wire [1:0] far_3_3688_0;    relay_conn far_3_3688_0_a(.in(layer_2[38]), .out(far_3_3688_0[0]));    relay_conn far_3_3688_0_b(.in(layer_2[3]), .out(far_3_3688_0[1]));
    assign layer_3[628] = ~far_3_3688_0[0] | (far_3_3688_0[0] & far_3_3688_0[1]); 
    assign layer_3[629] = ~layer_2[532]; 
    wire [1:0] far_3_3690_0;    relay_conn far_3_3690_0_a(.in(layer_2[245]), .out(far_3_3690_0[0]));    relay_conn far_3_3690_0_b(.in(layer_2[143]), .out(far_3_3690_0[1]));
    wire [1:0] far_3_3690_1;    relay_conn far_3_3690_1_a(.in(far_3_3690_0[0]), .out(far_3_3690_1[0]));    relay_conn far_3_3690_1_b(.in(far_3_3690_0[1]), .out(far_3_3690_1[1]));
    wire [1:0] far_3_3690_2;    relay_conn far_3_3690_2_a(.in(far_3_3690_1[0]), .out(far_3_3690_2[0]));    relay_conn far_3_3690_2_b(.in(far_3_3690_1[1]), .out(far_3_3690_2[1]));
    assign layer_3[630] = ~far_3_3690_2[0]; 
    assign layer_3[631] = ~(layer_2[43] | layer_2[56]); 
    wire [1:0] far_3_3692_0;    relay_conn far_3_3692_0_a(.in(layer_2[827]), .out(far_3_3692_0[0]));    relay_conn far_3_3692_0_b(.in(layer_2[784]), .out(far_3_3692_0[1]));
    assign layer_3[632] = ~far_3_3692_0[0]; 
    wire [1:0] far_3_3693_0;    relay_conn far_3_3693_0_a(.in(layer_2[716]), .out(far_3_3693_0[0]));    relay_conn far_3_3693_0_b(.in(layer_2[749]), .out(far_3_3693_0[1]));
    assign layer_3[633] = far_3_3693_0[1] & ~far_3_3693_0[0]; 
    wire [1:0] far_3_3694_0;    relay_conn far_3_3694_0_a(.in(layer_2[83]), .out(far_3_3694_0[0]));    relay_conn far_3_3694_0_b(.in(layer_2[35]), .out(far_3_3694_0[1]));
    assign layer_3[634] = ~far_3_3694_0[1]; 
    wire [1:0] far_3_3695_0;    relay_conn far_3_3695_0_a(.in(layer_2[281]), .out(far_3_3695_0[0]));    relay_conn far_3_3695_0_b(.in(layer_2[188]), .out(far_3_3695_0[1]));
    wire [1:0] far_3_3695_1;    relay_conn far_3_3695_1_a(.in(far_3_3695_0[0]), .out(far_3_3695_1[0]));    relay_conn far_3_3695_1_b(.in(far_3_3695_0[1]), .out(far_3_3695_1[1]));
    assign layer_3[635] = ~(far_3_3695_1[0] ^ far_3_3695_1[1]); 
    wire [1:0] far_3_3696_0;    relay_conn far_3_3696_0_a(.in(layer_2[709]), .out(far_3_3696_0[0]));    relay_conn far_3_3696_0_b(.in(layer_2[643]), .out(far_3_3696_0[1]));
    wire [1:0] far_3_3696_1;    relay_conn far_3_3696_1_a(.in(far_3_3696_0[0]), .out(far_3_3696_1[0]));    relay_conn far_3_3696_1_b(.in(far_3_3696_0[1]), .out(far_3_3696_1[1]));
    assign layer_3[636] = far_3_3696_1[0] & ~far_3_3696_1[1]; 
    wire [1:0] far_3_3697_0;    relay_conn far_3_3697_0_a(.in(layer_2[708]), .out(far_3_3697_0[0]));    relay_conn far_3_3697_0_b(.in(layer_2[580]), .out(far_3_3697_0[1]));
    wire [1:0] far_3_3697_1;    relay_conn far_3_3697_1_a(.in(far_3_3697_0[0]), .out(far_3_3697_1[0]));    relay_conn far_3_3697_1_b(.in(far_3_3697_0[1]), .out(far_3_3697_1[1]));
    wire [1:0] far_3_3697_2;    relay_conn far_3_3697_2_a(.in(far_3_3697_1[0]), .out(far_3_3697_2[0]));    relay_conn far_3_3697_2_b(.in(far_3_3697_1[1]), .out(far_3_3697_2[1]));
    wire [1:0] far_3_3697_3;    relay_conn far_3_3697_3_a(.in(far_3_3697_2[0]), .out(far_3_3697_3[0]));    relay_conn far_3_3697_3_b(.in(far_3_3697_2[1]), .out(far_3_3697_3[1]));
    assign layer_3[637] = far_3_3697_3[0] | far_3_3697_3[1]; 
    wire [1:0] far_3_3698_0;    relay_conn far_3_3698_0_a(.in(layer_2[433]), .out(far_3_3698_0[0]));    relay_conn far_3_3698_0_b(.in(layer_2[330]), .out(far_3_3698_0[1]));
    wire [1:0] far_3_3698_1;    relay_conn far_3_3698_1_a(.in(far_3_3698_0[0]), .out(far_3_3698_1[0]));    relay_conn far_3_3698_1_b(.in(far_3_3698_0[1]), .out(far_3_3698_1[1]));
    wire [1:0] far_3_3698_2;    relay_conn far_3_3698_2_a(.in(far_3_3698_1[0]), .out(far_3_3698_2[0]));    relay_conn far_3_3698_2_b(.in(far_3_3698_1[1]), .out(far_3_3698_2[1]));
    assign layer_3[638] = ~(far_3_3698_2[0] ^ far_3_3698_2[1]); 
    wire [1:0] far_3_3699_0;    relay_conn far_3_3699_0_a(.in(layer_2[915]), .out(far_3_3699_0[0]));    relay_conn far_3_3699_0_b(.in(layer_2[955]), .out(far_3_3699_0[1]));
    assign layer_3[639] = ~far_3_3699_0[1]; 
    wire [1:0] far_3_3700_0;    relay_conn far_3_3700_0_a(.in(layer_2[949]), .out(far_3_3700_0[0]));    relay_conn far_3_3700_0_b(.in(layer_2[987]), .out(far_3_3700_0[1]));
    assign layer_3[640] = far_3_3700_0[1]; 
    wire [1:0] far_3_3701_0;    relay_conn far_3_3701_0_a(.in(layer_2[257]), .out(far_3_3701_0[0]));    relay_conn far_3_3701_0_b(.in(layer_2[306]), .out(far_3_3701_0[1]));
    assign layer_3[641] = ~far_3_3701_0[1]; 
    wire [1:0] far_3_3702_0;    relay_conn far_3_3702_0_a(.in(layer_2[855]), .out(far_3_3702_0[0]));    relay_conn far_3_3702_0_b(.in(layer_2[949]), .out(far_3_3702_0[1]));
    wire [1:0] far_3_3702_1;    relay_conn far_3_3702_1_a(.in(far_3_3702_0[0]), .out(far_3_3702_1[0]));    relay_conn far_3_3702_1_b(.in(far_3_3702_0[1]), .out(far_3_3702_1[1]));
    assign layer_3[642] = ~far_3_3702_1[1] | (far_3_3702_1[0] & far_3_3702_1[1]); 
    wire [1:0] far_3_3703_0;    relay_conn far_3_3703_0_a(.in(layer_2[191]), .out(far_3_3703_0[0]));    relay_conn far_3_3703_0_b(.in(layer_2[118]), .out(far_3_3703_0[1]));
    wire [1:0] far_3_3703_1;    relay_conn far_3_3703_1_a(.in(far_3_3703_0[0]), .out(far_3_3703_1[0]));    relay_conn far_3_3703_1_b(.in(far_3_3703_0[1]), .out(far_3_3703_1[1]));
    assign layer_3[643] = ~far_3_3703_1[0] | (far_3_3703_1[0] & far_3_3703_1[1]); 
    wire [1:0] far_3_3704_0;    relay_conn far_3_3704_0_a(.in(layer_2[548]), .out(far_3_3704_0[0]));    relay_conn far_3_3704_0_b(.in(layer_2[673]), .out(far_3_3704_0[1]));
    wire [1:0] far_3_3704_1;    relay_conn far_3_3704_1_a(.in(far_3_3704_0[0]), .out(far_3_3704_1[0]));    relay_conn far_3_3704_1_b(.in(far_3_3704_0[1]), .out(far_3_3704_1[1]));
    wire [1:0] far_3_3704_2;    relay_conn far_3_3704_2_a(.in(far_3_3704_1[0]), .out(far_3_3704_2[0]));    relay_conn far_3_3704_2_b(.in(far_3_3704_1[1]), .out(far_3_3704_2[1]));
    assign layer_3[644] = ~far_3_3704_2[0] | (far_3_3704_2[0] & far_3_3704_2[1]); 
    assign layer_3[645] = layer_2[513] & layer_2[539]; 
    wire [1:0] far_3_3706_0;    relay_conn far_3_3706_0_a(.in(layer_2[507]), .out(far_3_3706_0[0]));    relay_conn far_3_3706_0_b(.in(layer_2[610]), .out(far_3_3706_0[1]));
    wire [1:0] far_3_3706_1;    relay_conn far_3_3706_1_a(.in(far_3_3706_0[0]), .out(far_3_3706_1[0]));    relay_conn far_3_3706_1_b(.in(far_3_3706_0[1]), .out(far_3_3706_1[1]));
    wire [1:0] far_3_3706_2;    relay_conn far_3_3706_2_a(.in(far_3_3706_1[0]), .out(far_3_3706_2[0]));    relay_conn far_3_3706_2_b(.in(far_3_3706_1[1]), .out(far_3_3706_2[1]));
    assign layer_3[646] = far_3_3706_2[0]; 
    wire [1:0] far_3_3707_0;    relay_conn far_3_3707_0_a(.in(layer_2[239]), .out(far_3_3707_0[0]));    relay_conn far_3_3707_0_b(.in(layer_2[129]), .out(far_3_3707_0[1]));
    wire [1:0] far_3_3707_1;    relay_conn far_3_3707_1_a(.in(far_3_3707_0[0]), .out(far_3_3707_1[0]));    relay_conn far_3_3707_1_b(.in(far_3_3707_0[1]), .out(far_3_3707_1[1]));
    wire [1:0] far_3_3707_2;    relay_conn far_3_3707_2_a(.in(far_3_3707_1[0]), .out(far_3_3707_2[0]));    relay_conn far_3_3707_2_b(.in(far_3_3707_1[1]), .out(far_3_3707_2[1]));
    assign layer_3[647] = far_3_3707_2[0] & ~far_3_3707_2[1]; 
    wire [1:0] far_3_3708_0;    relay_conn far_3_3708_0_a(.in(layer_2[839]), .out(far_3_3708_0[0]));    relay_conn far_3_3708_0_b(.in(layer_2[910]), .out(far_3_3708_0[1]));
    wire [1:0] far_3_3708_1;    relay_conn far_3_3708_1_a(.in(far_3_3708_0[0]), .out(far_3_3708_1[0]));    relay_conn far_3_3708_1_b(.in(far_3_3708_0[1]), .out(far_3_3708_1[1]));
    assign layer_3[648] = far_3_3708_1[0] & far_3_3708_1[1]; 
    wire [1:0] far_3_3709_0;    relay_conn far_3_3709_0_a(.in(layer_2[300]), .out(far_3_3709_0[0]));    relay_conn far_3_3709_0_b(.in(layer_2[205]), .out(far_3_3709_0[1]));
    wire [1:0] far_3_3709_1;    relay_conn far_3_3709_1_a(.in(far_3_3709_0[0]), .out(far_3_3709_1[0]));    relay_conn far_3_3709_1_b(.in(far_3_3709_0[1]), .out(far_3_3709_1[1]));
    assign layer_3[649] = far_3_3709_1[0] & far_3_3709_1[1]; 
    wire [1:0] far_3_3710_0;    relay_conn far_3_3710_0_a(.in(layer_2[906]), .out(far_3_3710_0[0]));    relay_conn far_3_3710_0_b(.in(layer_2[1015]), .out(far_3_3710_0[1]));
    wire [1:0] far_3_3710_1;    relay_conn far_3_3710_1_a(.in(far_3_3710_0[0]), .out(far_3_3710_1[0]));    relay_conn far_3_3710_1_b(.in(far_3_3710_0[1]), .out(far_3_3710_1[1]));
    wire [1:0] far_3_3710_2;    relay_conn far_3_3710_2_a(.in(far_3_3710_1[0]), .out(far_3_3710_2[0]));    relay_conn far_3_3710_2_b(.in(far_3_3710_1[1]), .out(far_3_3710_2[1]));
    assign layer_3[650] = far_3_3710_2[0] & far_3_3710_2[1]; 
    assign layer_3[651] = layer_2[907] | layer_2[891]; 
    assign layer_3[652] = ~layer_2[281]; 
    assign layer_3[653] = ~layer_2[738] | (layer_2[757] & layer_2[738]); 
    wire [1:0] far_3_3714_0;    relay_conn far_3_3714_0_a(.in(layer_2[143]), .out(far_3_3714_0[0]));    relay_conn far_3_3714_0_b(.in(layer_2[215]), .out(far_3_3714_0[1]));
    wire [1:0] far_3_3714_1;    relay_conn far_3_3714_1_a(.in(far_3_3714_0[0]), .out(far_3_3714_1[0]));    relay_conn far_3_3714_1_b(.in(far_3_3714_0[1]), .out(far_3_3714_1[1]));
    assign layer_3[654] = far_3_3714_1[0] & ~far_3_3714_1[1]; 
    wire [1:0] far_3_3715_0;    relay_conn far_3_3715_0_a(.in(layer_2[129]), .out(far_3_3715_0[0]));    relay_conn far_3_3715_0_b(.in(layer_2[208]), .out(far_3_3715_0[1]));
    wire [1:0] far_3_3715_1;    relay_conn far_3_3715_1_a(.in(far_3_3715_0[0]), .out(far_3_3715_1[0]));    relay_conn far_3_3715_1_b(.in(far_3_3715_0[1]), .out(far_3_3715_1[1]));
    assign layer_3[655] = ~(far_3_3715_1[0] & far_3_3715_1[1]); 
    wire [1:0] far_3_3716_0;    relay_conn far_3_3716_0_a(.in(layer_2[912]), .out(far_3_3716_0[0]));    relay_conn far_3_3716_0_b(.in(layer_2[859]), .out(far_3_3716_0[1]));
    assign layer_3[656] = ~far_3_3716_0[0] | (far_3_3716_0[0] & far_3_3716_0[1]); 
    assign layer_3[657] = layer_2[958] & ~layer_2[927]; 
    wire [1:0] far_3_3718_0;    relay_conn far_3_3718_0_a(.in(layer_2[854]), .out(far_3_3718_0[0]));    relay_conn far_3_3718_0_b(.in(layer_2[970]), .out(far_3_3718_0[1]));
    wire [1:0] far_3_3718_1;    relay_conn far_3_3718_1_a(.in(far_3_3718_0[0]), .out(far_3_3718_1[0]));    relay_conn far_3_3718_1_b(.in(far_3_3718_0[1]), .out(far_3_3718_1[1]));
    wire [1:0] far_3_3718_2;    relay_conn far_3_3718_2_a(.in(far_3_3718_1[0]), .out(far_3_3718_2[0]));    relay_conn far_3_3718_2_b(.in(far_3_3718_1[1]), .out(far_3_3718_2[1]));
    assign layer_3[658] = far_3_3718_2[0] & ~far_3_3718_2[1]; 
    wire [1:0] far_3_3719_0;    relay_conn far_3_3719_0_a(.in(layer_2[777]), .out(far_3_3719_0[0]));    relay_conn far_3_3719_0_b(.in(layer_2[845]), .out(far_3_3719_0[1]));
    wire [1:0] far_3_3719_1;    relay_conn far_3_3719_1_a(.in(far_3_3719_0[0]), .out(far_3_3719_1[0]));    relay_conn far_3_3719_1_b(.in(far_3_3719_0[1]), .out(far_3_3719_1[1]));
    assign layer_3[659] = far_3_3719_1[0]; 
    wire [1:0] far_3_3720_0;    relay_conn far_3_3720_0_a(.in(layer_2[120]), .out(far_3_3720_0[0]));    relay_conn far_3_3720_0_b(.in(layer_2[239]), .out(far_3_3720_0[1]));
    wire [1:0] far_3_3720_1;    relay_conn far_3_3720_1_a(.in(far_3_3720_0[0]), .out(far_3_3720_1[0]));    relay_conn far_3_3720_1_b(.in(far_3_3720_0[1]), .out(far_3_3720_1[1]));
    wire [1:0] far_3_3720_2;    relay_conn far_3_3720_2_a(.in(far_3_3720_1[0]), .out(far_3_3720_2[0]));    relay_conn far_3_3720_2_b(.in(far_3_3720_1[1]), .out(far_3_3720_2[1]));
    assign layer_3[660] = far_3_3720_2[0] & ~far_3_3720_2[1]; 
    assign layer_3[661] = ~(layer_2[779] & layer_2[785]); 
    assign layer_3[662] = ~(layer_2[234] ^ layer_2[238]); 
    assign layer_3[663] = ~(layer_2[144] & layer_2[137]); 
    assign layer_3[664] = layer_2[341] | layer_2[320]; 
    wire [1:0] far_3_3725_0;    relay_conn far_3_3725_0_a(.in(layer_2[332]), .out(far_3_3725_0[0]));    relay_conn far_3_3725_0_b(.in(layer_2[378]), .out(far_3_3725_0[1]));
    assign layer_3[665] = far_3_3725_0[0]; 
    wire [1:0] far_3_3726_0;    relay_conn far_3_3726_0_a(.in(layer_2[241]), .out(far_3_3726_0[0]));    relay_conn far_3_3726_0_b(.in(layer_2[289]), .out(far_3_3726_0[1]));
    assign layer_3[666] = ~far_3_3726_0[0] | (far_3_3726_0[0] & far_3_3726_0[1]); 
    wire [1:0] far_3_3727_0;    relay_conn far_3_3727_0_a(.in(layer_2[233]), .out(far_3_3727_0[0]));    relay_conn far_3_3727_0_b(.in(layer_2[167]), .out(far_3_3727_0[1]));
    wire [1:0] far_3_3727_1;    relay_conn far_3_3727_1_a(.in(far_3_3727_0[0]), .out(far_3_3727_1[0]));    relay_conn far_3_3727_1_b(.in(far_3_3727_0[1]), .out(far_3_3727_1[1]));
    assign layer_3[667] = ~(far_3_3727_1[0] & far_3_3727_1[1]); 
    wire [1:0] far_3_3728_0;    relay_conn far_3_3728_0_a(.in(layer_2[646]), .out(far_3_3728_0[0]));    relay_conn far_3_3728_0_b(.in(layer_2[769]), .out(far_3_3728_0[1]));
    wire [1:0] far_3_3728_1;    relay_conn far_3_3728_1_a(.in(far_3_3728_0[0]), .out(far_3_3728_1[0]));    relay_conn far_3_3728_1_b(.in(far_3_3728_0[1]), .out(far_3_3728_1[1]));
    wire [1:0] far_3_3728_2;    relay_conn far_3_3728_2_a(.in(far_3_3728_1[0]), .out(far_3_3728_2[0]));    relay_conn far_3_3728_2_b(.in(far_3_3728_1[1]), .out(far_3_3728_2[1]));
    assign layer_3[668] = ~far_3_3728_2[0]; 
    assign layer_3[669] = layer_2[136] | layer_2[126]; 
    wire [1:0] far_3_3730_0;    relay_conn far_3_3730_0_a(.in(layer_2[1002]), .out(far_3_3730_0[0]));    relay_conn far_3_3730_0_b(.in(layer_2[970]), .out(far_3_3730_0[1]));
    assign layer_3[670] = far_3_3730_0[0] & far_3_3730_0[1]; 
    wire [1:0] far_3_3731_0;    relay_conn far_3_3731_0_a(.in(layer_2[920]), .out(far_3_3731_0[0]));    relay_conn far_3_3731_0_b(.in(layer_2[839]), .out(far_3_3731_0[1]));
    wire [1:0] far_3_3731_1;    relay_conn far_3_3731_1_a(.in(far_3_3731_0[0]), .out(far_3_3731_1[0]));    relay_conn far_3_3731_1_b(.in(far_3_3731_0[1]), .out(far_3_3731_1[1]));
    assign layer_3[671] = far_3_3731_1[1]; 
    wire [1:0] far_3_3732_0;    relay_conn far_3_3732_0_a(.in(layer_2[748]), .out(far_3_3732_0[0]));    relay_conn far_3_3732_0_b(.in(layer_2[844]), .out(far_3_3732_0[1]));
    wire [1:0] far_3_3732_1;    relay_conn far_3_3732_1_a(.in(far_3_3732_0[0]), .out(far_3_3732_1[0]));    relay_conn far_3_3732_1_b(.in(far_3_3732_0[1]), .out(far_3_3732_1[1]));
    wire [1:0] far_3_3732_2;    relay_conn far_3_3732_2_a(.in(far_3_3732_1[0]), .out(far_3_3732_2[0]));    relay_conn far_3_3732_2_b(.in(far_3_3732_1[1]), .out(far_3_3732_2[1]));
    assign layer_3[672] = ~far_3_3732_2[0] | (far_3_3732_2[0] & far_3_3732_2[1]); 
    wire [1:0] far_3_3733_0;    relay_conn far_3_3733_0_a(.in(layer_2[245]), .out(far_3_3733_0[0]));    relay_conn far_3_3733_0_b(.in(layer_2[303]), .out(far_3_3733_0[1]));
    assign layer_3[673] = ~far_3_3733_0[0]; 
    wire [1:0] far_3_3734_0;    relay_conn far_3_3734_0_a(.in(layer_2[766]), .out(far_3_3734_0[0]));    relay_conn far_3_3734_0_b(.in(layer_2[888]), .out(far_3_3734_0[1]));
    wire [1:0] far_3_3734_1;    relay_conn far_3_3734_1_a(.in(far_3_3734_0[0]), .out(far_3_3734_1[0]));    relay_conn far_3_3734_1_b(.in(far_3_3734_0[1]), .out(far_3_3734_1[1]));
    wire [1:0] far_3_3734_2;    relay_conn far_3_3734_2_a(.in(far_3_3734_1[0]), .out(far_3_3734_2[0]));    relay_conn far_3_3734_2_b(.in(far_3_3734_1[1]), .out(far_3_3734_2[1]));
    assign layer_3[674] = far_3_3734_2[0] | far_3_3734_2[1]; 
    assign layer_3[675] = layer_2[775] & layer_2[802]; 
    wire [1:0] far_3_3736_0;    relay_conn far_3_3736_0_a(.in(layer_2[1001]), .out(far_3_3736_0[0]));    relay_conn far_3_3736_0_b(.in(layer_2[960]), .out(far_3_3736_0[1]));
    assign layer_3[676] = far_3_3736_0[0] | far_3_3736_0[1]; 
    assign layer_3[677] = ~(layer_2[27] | layer_2[23]); 
    wire [1:0] far_3_3738_0;    relay_conn far_3_3738_0_a(.in(layer_2[693]), .out(far_3_3738_0[0]));    relay_conn far_3_3738_0_b(.in(layer_2[752]), .out(far_3_3738_0[1]));
    assign layer_3[678] = far_3_3738_0[1] & ~far_3_3738_0[0]; 
    wire [1:0] far_3_3739_0;    relay_conn far_3_3739_0_a(.in(layer_2[252]), .out(far_3_3739_0[0]));    relay_conn far_3_3739_0_b(.in(layer_2[354]), .out(far_3_3739_0[1]));
    wire [1:0] far_3_3739_1;    relay_conn far_3_3739_1_a(.in(far_3_3739_0[0]), .out(far_3_3739_1[0]));    relay_conn far_3_3739_1_b(.in(far_3_3739_0[1]), .out(far_3_3739_1[1]));
    wire [1:0] far_3_3739_2;    relay_conn far_3_3739_2_a(.in(far_3_3739_1[0]), .out(far_3_3739_2[0]));    relay_conn far_3_3739_2_b(.in(far_3_3739_1[1]), .out(far_3_3739_2[1]));
    assign layer_3[679] = ~far_3_3739_2[1]; 
    wire [1:0] far_3_3740_0;    relay_conn far_3_3740_0_a(.in(layer_2[108]), .out(far_3_3740_0[0]));    relay_conn far_3_3740_0_b(.in(layer_2[56]), .out(far_3_3740_0[1]));
    assign layer_3[680] = far_3_3740_0[0] & far_3_3740_0[1]; 
    assign layer_3[681] = ~(layer_2[927] | layer_2[949]); 
    wire [1:0] far_3_3742_0;    relay_conn far_3_3742_0_a(.in(layer_2[1004]), .out(far_3_3742_0[0]));    relay_conn far_3_3742_0_b(.in(layer_2[927]), .out(far_3_3742_0[1]));
    wire [1:0] far_3_3742_1;    relay_conn far_3_3742_1_a(.in(far_3_3742_0[0]), .out(far_3_3742_1[0]));    relay_conn far_3_3742_1_b(.in(far_3_3742_0[1]), .out(far_3_3742_1[1]));
    assign layer_3[682] = ~(far_3_3742_1[0] | far_3_3742_1[1]); 
    wire [1:0] far_3_3743_0;    relay_conn far_3_3743_0_a(.in(layer_2[514]), .out(far_3_3743_0[0]));    relay_conn far_3_3743_0_b(.in(layer_2[389]), .out(far_3_3743_0[1]));
    wire [1:0] far_3_3743_1;    relay_conn far_3_3743_1_a(.in(far_3_3743_0[0]), .out(far_3_3743_1[0]));    relay_conn far_3_3743_1_b(.in(far_3_3743_0[1]), .out(far_3_3743_1[1]));
    wire [1:0] far_3_3743_2;    relay_conn far_3_3743_2_a(.in(far_3_3743_1[0]), .out(far_3_3743_2[0]));    relay_conn far_3_3743_2_b(.in(far_3_3743_1[1]), .out(far_3_3743_2[1]));
    assign layer_3[683] = ~(far_3_3743_2[0] ^ far_3_3743_2[1]); 
    wire [1:0] far_3_3744_0;    relay_conn far_3_3744_0_a(.in(layer_2[997]), .out(far_3_3744_0[0]));    relay_conn far_3_3744_0_b(.in(layer_2[913]), .out(far_3_3744_0[1]));
    wire [1:0] far_3_3744_1;    relay_conn far_3_3744_1_a(.in(far_3_3744_0[0]), .out(far_3_3744_1[0]));    relay_conn far_3_3744_1_b(.in(far_3_3744_0[1]), .out(far_3_3744_1[1]));
    assign layer_3[684] = far_3_3744_1[0] ^ far_3_3744_1[1]; 
    wire [1:0] far_3_3745_0;    relay_conn far_3_3745_0_a(.in(layer_2[191]), .out(far_3_3745_0[0]));    relay_conn far_3_3745_0_b(.in(layer_2[93]), .out(far_3_3745_0[1]));
    wire [1:0] far_3_3745_1;    relay_conn far_3_3745_1_a(.in(far_3_3745_0[0]), .out(far_3_3745_1[0]));    relay_conn far_3_3745_1_b(.in(far_3_3745_0[1]), .out(far_3_3745_1[1]));
    wire [1:0] far_3_3745_2;    relay_conn far_3_3745_2_a(.in(far_3_3745_1[0]), .out(far_3_3745_2[0]));    relay_conn far_3_3745_2_b(.in(far_3_3745_1[1]), .out(far_3_3745_2[1]));
    assign layer_3[685] = far_3_3745_2[1]; 
    wire [1:0] far_3_3746_0;    relay_conn far_3_3746_0_a(.in(layer_2[463]), .out(far_3_3746_0[0]));    relay_conn far_3_3746_0_b(.in(layer_2[379]), .out(far_3_3746_0[1]));
    wire [1:0] far_3_3746_1;    relay_conn far_3_3746_1_a(.in(far_3_3746_0[0]), .out(far_3_3746_1[0]));    relay_conn far_3_3746_1_b(.in(far_3_3746_0[1]), .out(far_3_3746_1[1]));
    assign layer_3[686] = ~(far_3_3746_1[0] & far_3_3746_1[1]); 
    wire [1:0] far_3_3747_0;    relay_conn far_3_3747_0_a(.in(layer_2[345]), .out(far_3_3747_0[0]));    relay_conn far_3_3747_0_b(.in(layer_2[412]), .out(far_3_3747_0[1]));
    wire [1:0] far_3_3747_1;    relay_conn far_3_3747_1_a(.in(far_3_3747_0[0]), .out(far_3_3747_1[0]));    relay_conn far_3_3747_1_b(.in(far_3_3747_0[1]), .out(far_3_3747_1[1]));
    assign layer_3[687] = ~(far_3_3747_1[0] ^ far_3_3747_1[1]); 
    wire [1:0] far_3_3748_0;    relay_conn far_3_3748_0_a(.in(layer_2[683]), .out(far_3_3748_0[0]));    relay_conn far_3_3748_0_b(.in(layer_2[801]), .out(far_3_3748_0[1]));
    wire [1:0] far_3_3748_1;    relay_conn far_3_3748_1_a(.in(far_3_3748_0[0]), .out(far_3_3748_1[0]));    relay_conn far_3_3748_1_b(.in(far_3_3748_0[1]), .out(far_3_3748_1[1]));
    wire [1:0] far_3_3748_2;    relay_conn far_3_3748_2_a(.in(far_3_3748_1[0]), .out(far_3_3748_2[0]));    relay_conn far_3_3748_2_b(.in(far_3_3748_1[1]), .out(far_3_3748_2[1]));
    assign layer_3[688] = ~(far_3_3748_2[0] | far_3_3748_2[1]); 
    assign layer_3[689] = ~layer_2[58] | (layer_2[58] & layer_2[75]); 
    wire [1:0] far_3_3750_0;    relay_conn far_3_3750_0_a(.in(layer_2[463]), .out(far_3_3750_0[0]));    relay_conn far_3_3750_0_b(.in(layer_2[508]), .out(far_3_3750_0[1]));
    assign layer_3[690] = ~far_3_3750_0[0]; 
    wire [1:0] far_3_3751_0;    relay_conn far_3_3751_0_a(.in(layer_2[716]), .out(far_3_3751_0[0]));    relay_conn far_3_3751_0_b(.in(layer_2[597]), .out(far_3_3751_0[1]));
    wire [1:0] far_3_3751_1;    relay_conn far_3_3751_1_a(.in(far_3_3751_0[0]), .out(far_3_3751_1[0]));    relay_conn far_3_3751_1_b(.in(far_3_3751_0[1]), .out(far_3_3751_1[1]));
    wire [1:0] far_3_3751_2;    relay_conn far_3_3751_2_a(.in(far_3_3751_1[0]), .out(far_3_3751_2[0]));    relay_conn far_3_3751_2_b(.in(far_3_3751_1[1]), .out(far_3_3751_2[1]));
    assign layer_3[691] = far_3_3751_2[1] & ~far_3_3751_2[0]; 
    assign layer_3[692] = layer_2[865] & ~layer_2[866]; 
    wire [1:0] far_3_3753_0;    relay_conn far_3_3753_0_a(.in(layer_2[462]), .out(far_3_3753_0[0]));    relay_conn far_3_3753_0_b(.in(layer_2[543]), .out(far_3_3753_0[1]));
    wire [1:0] far_3_3753_1;    relay_conn far_3_3753_1_a(.in(far_3_3753_0[0]), .out(far_3_3753_1[0]));    relay_conn far_3_3753_1_b(.in(far_3_3753_0[1]), .out(far_3_3753_1[1]));
    assign layer_3[693] = ~far_3_3753_1[0]; 
    wire [1:0] far_3_3754_0;    relay_conn far_3_3754_0_a(.in(layer_2[768]), .out(far_3_3754_0[0]));    relay_conn far_3_3754_0_b(.in(layer_2[709]), .out(far_3_3754_0[1]));
    assign layer_3[694] = ~far_3_3754_0[0] | (far_3_3754_0[0] & far_3_3754_0[1]); 
    wire [1:0] far_3_3755_0;    relay_conn far_3_3755_0_a(.in(layer_2[341]), .out(far_3_3755_0[0]));    relay_conn far_3_3755_0_b(.in(layer_2[434]), .out(far_3_3755_0[1]));
    wire [1:0] far_3_3755_1;    relay_conn far_3_3755_1_a(.in(far_3_3755_0[0]), .out(far_3_3755_1[0]));    relay_conn far_3_3755_1_b(.in(far_3_3755_0[1]), .out(far_3_3755_1[1]));
    assign layer_3[695] = ~far_3_3755_1[0] | (far_3_3755_1[0] & far_3_3755_1[1]); 
    wire [1:0] far_3_3756_0;    relay_conn far_3_3756_0_a(.in(layer_2[742]), .out(far_3_3756_0[0]));    relay_conn far_3_3756_0_b(.in(layer_2[687]), .out(far_3_3756_0[1]));
    assign layer_3[696] = far_3_3756_0[0] & ~far_3_3756_0[1]; 
    wire [1:0] far_3_3757_0;    relay_conn far_3_3757_0_a(.in(layer_2[227]), .out(far_3_3757_0[0]));    relay_conn far_3_3757_0_b(.in(layer_2[132]), .out(far_3_3757_0[1]));
    wire [1:0] far_3_3757_1;    relay_conn far_3_3757_1_a(.in(far_3_3757_0[0]), .out(far_3_3757_1[0]));    relay_conn far_3_3757_1_b(.in(far_3_3757_0[1]), .out(far_3_3757_1[1]));
    assign layer_3[697] = ~far_3_3757_1[0]; 
    wire [1:0] far_3_3758_0;    relay_conn far_3_3758_0_a(.in(layer_2[785]), .out(far_3_3758_0[0]));    relay_conn far_3_3758_0_b(.in(layer_2[910]), .out(far_3_3758_0[1]));
    wire [1:0] far_3_3758_1;    relay_conn far_3_3758_1_a(.in(far_3_3758_0[0]), .out(far_3_3758_1[0]));    relay_conn far_3_3758_1_b(.in(far_3_3758_0[1]), .out(far_3_3758_1[1]));
    wire [1:0] far_3_3758_2;    relay_conn far_3_3758_2_a(.in(far_3_3758_1[0]), .out(far_3_3758_2[0]));    relay_conn far_3_3758_2_b(.in(far_3_3758_1[1]), .out(far_3_3758_2[1]));
    assign layer_3[698] = far_3_3758_2[0] | far_3_3758_2[1]; 
    wire [1:0] far_3_3759_0;    relay_conn far_3_3759_0_a(.in(layer_2[500]), .out(far_3_3759_0[0]));    relay_conn far_3_3759_0_b(.in(layer_2[440]), .out(far_3_3759_0[1]));
    assign layer_3[699] = ~(far_3_3759_0[0] | far_3_3759_0[1]); 
    assign layer_3[700] = layer_2[774] & ~layer_2[794]; 
    assign layer_3[701] = ~layer_2[892] | (layer_2[892] & layer_2[877]); 
    wire [1:0] far_3_3762_0;    relay_conn far_3_3762_0_a(.in(layer_2[539]), .out(far_3_3762_0[0]));    relay_conn far_3_3762_0_b(.in(layer_2[492]), .out(far_3_3762_0[1]));
    assign layer_3[702] = ~(far_3_3762_0[0] & far_3_3762_0[1]); 
    assign layer_3[703] = ~layer_2[844] | (layer_2[844] & layer_2[819]); 
    wire [1:0] far_3_3764_0;    relay_conn far_3_3764_0_a(.in(layer_2[256]), .out(far_3_3764_0[0]));    relay_conn far_3_3764_0_b(.in(layer_2[325]), .out(far_3_3764_0[1]));
    wire [1:0] far_3_3764_1;    relay_conn far_3_3764_1_a(.in(far_3_3764_0[0]), .out(far_3_3764_1[0]));    relay_conn far_3_3764_1_b(.in(far_3_3764_0[1]), .out(far_3_3764_1[1]));
    assign layer_3[704] = far_3_3764_1[0] | far_3_3764_1[1]; 
    wire [1:0] far_3_3765_0;    relay_conn far_3_3765_0_a(.in(layer_2[200]), .out(far_3_3765_0[0]));    relay_conn far_3_3765_0_b(.in(layer_2[284]), .out(far_3_3765_0[1]));
    wire [1:0] far_3_3765_1;    relay_conn far_3_3765_1_a(.in(far_3_3765_0[0]), .out(far_3_3765_1[0]));    relay_conn far_3_3765_1_b(.in(far_3_3765_0[1]), .out(far_3_3765_1[1]));
    assign layer_3[705] = far_3_3765_1[1]; 
    wire [1:0] far_3_3766_0;    relay_conn far_3_3766_0_a(.in(layer_2[1011]), .out(far_3_3766_0[0]));    relay_conn far_3_3766_0_b(.in(layer_2[891]), .out(far_3_3766_0[1]));
    wire [1:0] far_3_3766_1;    relay_conn far_3_3766_1_a(.in(far_3_3766_0[0]), .out(far_3_3766_1[0]));    relay_conn far_3_3766_1_b(.in(far_3_3766_0[1]), .out(far_3_3766_1[1]));
    wire [1:0] far_3_3766_2;    relay_conn far_3_3766_2_a(.in(far_3_3766_1[0]), .out(far_3_3766_2[0]));    relay_conn far_3_3766_2_b(.in(far_3_3766_1[1]), .out(far_3_3766_2[1]));
    assign layer_3[706] = ~far_3_3766_2[0] | (far_3_3766_2[0] & far_3_3766_2[1]); 
    wire [1:0] far_3_3767_0;    relay_conn far_3_3767_0_a(.in(layer_2[198]), .out(far_3_3767_0[0]));    relay_conn far_3_3767_0_b(.in(layer_2[232]), .out(far_3_3767_0[1]));
    assign layer_3[707] = ~(far_3_3767_0[0] | far_3_3767_0[1]); 
    wire [1:0] far_3_3768_0;    relay_conn far_3_3768_0_a(.in(layer_2[836]), .out(far_3_3768_0[0]));    relay_conn far_3_3768_0_b(.in(layer_2[791]), .out(far_3_3768_0[1]));
    assign layer_3[708] = ~far_3_3768_0[1]; 
    assign layer_3[709] = layer_2[6]; 
    wire [1:0] far_3_3770_0;    relay_conn far_3_3770_0_a(.in(layer_2[685]), .out(far_3_3770_0[0]));    relay_conn far_3_3770_0_b(.in(layer_2[774]), .out(far_3_3770_0[1]));
    wire [1:0] far_3_3770_1;    relay_conn far_3_3770_1_a(.in(far_3_3770_0[0]), .out(far_3_3770_1[0]));    relay_conn far_3_3770_1_b(.in(far_3_3770_0[1]), .out(far_3_3770_1[1]));
    assign layer_3[710] = far_3_3770_1[0] | far_3_3770_1[1]; 
    wire [1:0] far_3_3771_0;    relay_conn far_3_3771_0_a(.in(layer_2[850]), .out(far_3_3771_0[0]));    relay_conn far_3_3771_0_b(.in(layer_2[927]), .out(far_3_3771_0[1]));
    wire [1:0] far_3_3771_1;    relay_conn far_3_3771_1_a(.in(far_3_3771_0[0]), .out(far_3_3771_1[0]));    relay_conn far_3_3771_1_b(.in(far_3_3771_0[1]), .out(far_3_3771_1[1]));
    assign layer_3[711] = ~far_3_3771_1[1]; 
    assign layer_3[712] = layer_2[960] | layer_2[988]; 
    wire [1:0] far_3_3773_0;    relay_conn far_3_3773_0_a(.in(layer_2[1014]), .out(far_3_3773_0[0]));    relay_conn far_3_3773_0_b(.in(layer_2[978]), .out(far_3_3773_0[1]));
    assign layer_3[713] = ~far_3_3773_0[1] | (far_3_3773_0[0] & far_3_3773_0[1]); 
    wire [1:0] far_3_3774_0;    relay_conn far_3_3774_0_a(.in(layer_2[212]), .out(far_3_3774_0[0]));    relay_conn far_3_3774_0_b(.in(layer_2[284]), .out(far_3_3774_0[1]));
    wire [1:0] far_3_3774_1;    relay_conn far_3_3774_1_a(.in(far_3_3774_0[0]), .out(far_3_3774_1[0]));    relay_conn far_3_3774_1_b(.in(far_3_3774_0[1]), .out(far_3_3774_1[1]));
    assign layer_3[714] = far_3_3774_1[1] & ~far_3_3774_1[0]; 
    assign layer_3[715] = layer_2[498]; 
    assign layer_3[716] = ~(layer_2[211] & layer_2[205]); 
    wire [1:0] far_3_3777_0;    relay_conn far_3_3777_0_a(.in(layer_2[742]), .out(far_3_3777_0[0]));    relay_conn far_3_3777_0_b(.in(layer_2[824]), .out(far_3_3777_0[1]));
    wire [1:0] far_3_3777_1;    relay_conn far_3_3777_1_a(.in(far_3_3777_0[0]), .out(far_3_3777_1[0]));    relay_conn far_3_3777_1_b(.in(far_3_3777_0[1]), .out(far_3_3777_1[1]));
    assign layer_3[717] = far_3_3777_1[1]; 
    wire [1:0] far_3_3778_0;    relay_conn far_3_3778_0_a(.in(layer_2[246]), .out(far_3_3778_0[0]));    relay_conn far_3_3778_0_b(.in(layer_2[357]), .out(far_3_3778_0[1]));
    wire [1:0] far_3_3778_1;    relay_conn far_3_3778_1_a(.in(far_3_3778_0[0]), .out(far_3_3778_1[0]));    relay_conn far_3_3778_1_b(.in(far_3_3778_0[1]), .out(far_3_3778_1[1]));
    wire [1:0] far_3_3778_2;    relay_conn far_3_3778_2_a(.in(far_3_3778_1[0]), .out(far_3_3778_2[0]));    relay_conn far_3_3778_2_b(.in(far_3_3778_1[1]), .out(far_3_3778_2[1]));
    assign layer_3[718] = far_3_3778_2[0]; 
    assign layer_3[719] = layer_2[440]; 
    wire [1:0] far_3_3780_0;    relay_conn far_3_3780_0_a(.in(layer_2[328]), .out(far_3_3780_0[0]));    relay_conn far_3_3780_0_b(.in(layer_2[381]), .out(far_3_3780_0[1]));
    assign layer_3[720] = ~(far_3_3780_0[0] ^ far_3_3780_0[1]); 
    wire [1:0] far_3_3781_0;    relay_conn far_3_3781_0_a(.in(layer_2[872]), .out(far_3_3781_0[0]));    relay_conn far_3_3781_0_b(.in(layer_2[952]), .out(far_3_3781_0[1]));
    wire [1:0] far_3_3781_1;    relay_conn far_3_3781_1_a(.in(far_3_3781_0[0]), .out(far_3_3781_1[0]));    relay_conn far_3_3781_1_b(.in(far_3_3781_0[1]), .out(far_3_3781_1[1]));
    assign layer_3[721] = ~far_3_3781_1[1]; 
    wire [1:0] far_3_3782_0;    relay_conn far_3_3782_0_a(.in(layer_2[485]), .out(far_3_3782_0[0]));    relay_conn far_3_3782_0_b(.in(layer_2[357]), .out(far_3_3782_0[1]));
    wire [1:0] far_3_3782_1;    relay_conn far_3_3782_1_a(.in(far_3_3782_0[0]), .out(far_3_3782_1[0]));    relay_conn far_3_3782_1_b(.in(far_3_3782_0[1]), .out(far_3_3782_1[1]));
    wire [1:0] far_3_3782_2;    relay_conn far_3_3782_2_a(.in(far_3_3782_1[0]), .out(far_3_3782_2[0]));    relay_conn far_3_3782_2_b(.in(far_3_3782_1[1]), .out(far_3_3782_2[1]));
    wire [1:0] far_3_3782_3;    relay_conn far_3_3782_3_a(.in(far_3_3782_2[0]), .out(far_3_3782_3[0]));    relay_conn far_3_3782_3_b(.in(far_3_3782_2[1]), .out(far_3_3782_3[1]));
    assign layer_3[722] = ~far_3_3782_3[1] | (far_3_3782_3[0] & far_3_3782_3[1]); 
    wire [1:0] far_3_3783_0;    relay_conn far_3_3783_0_a(.in(layer_2[283]), .out(far_3_3783_0[0]));    relay_conn far_3_3783_0_b(.in(layer_2[361]), .out(far_3_3783_0[1]));
    wire [1:0] far_3_3783_1;    relay_conn far_3_3783_1_a(.in(far_3_3783_0[0]), .out(far_3_3783_1[0]));    relay_conn far_3_3783_1_b(.in(far_3_3783_0[1]), .out(far_3_3783_1[1]));
    assign layer_3[723] = ~(far_3_3783_1[0] ^ far_3_3783_1[1]); 
    wire [1:0] far_3_3784_0;    relay_conn far_3_3784_0_a(.in(layer_2[35]), .out(far_3_3784_0[0]));    relay_conn far_3_3784_0_b(.in(layer_2[126]), .out(far_3_3784_0[1]));
    wire [1:0] far_3_3784_1;    relay_conn far_3_3784_1_a(.in(far_3_3784_0[0]), .out(far_3_3784_1[0]));    relay_conn far_3_3784_1_b(.in(far_3_3784_0[1]), .out(far_3_3784_1[1]));
    assign layer_3[724] = far_3_3784_1[0] ^ far_3_3784_1[1]; 
    wire [1:0] far_3_3785_0;    relay_conn far_3_3785_0_a(.in(layer_2[341]), .out(far_3_3785_0[0]));    relay_conn far_3_3785_0_b(.in(layer_2[309]), .out(far_3_3785_0[1]));
    assign layer_3[725] = ~(far_3_3785_0[0] & far_3_3785_0[1]); 
    wire [1:0] far_3_3786_0;    relay_conn far_3_3786_0_a(.in(layer_2[921]), .out(far_3_3786_0[0]));    relay_conn far_3_3786_0_b(.in(layer_2[835]), .out(far_3_3786_0[1]));
    wire [1:0] far_3_3786_1;    relay_conn far_3_3786_1_a(.in(far_3_3786_0[0]), .out(far_3_3786_1[0]));    relay_conn far_3_3786_1_b(.in(far_3_3786_0[1]), .out(far_3_3786_1[1]));
    assign layer_3[726] = ~far_3_3786_1[0]; 
    assign layer_3[727] = layer_2[729] | layer_2[749]; 
    wire [1:0] far_3_3788_0;    relay_conn far_3_3788_0_a(.in(layer_2[267]), .out(far_3_3788_0[0]));    relay_conn far_3_3788_0_b(.in(layer_2[154]), .out(far_3_3788_0[1]));
    wire [1:0] far_3_3788_1;    relay_conn far_3_3788_1_a(.in(far_3_3788_0[0]), .out(far_3_3788_1[0]));    relay_conn far_3_3788_1_b(.in(far_3_3788_0[1]), .out(far_3_3788_1[1]));
    wire [1:0] far_3_3788_2;    relay_conn far_3_3788_2_a(.in(far_3_3788_1[0]), .out(far_3_3788_2[0]));    relay_conn far_3_3788_2_b(.in(far_3_3788_1[1]), .out(far_3_3788_2[1]));
    assign layer_3[728] = far_3_3788_2[1] & ~far_3_3788_2[0]; 
    assign layer_3[729] = layer_2[207]; 
    wire [1:0] far_3_3790_0;    relay_conn far_3_3790_0_a(.in(layer_2[299]), .out(far_3_3790_0[0]));    relay_conn far_3_3790_0_b(.in(layer_2[398]), .out(far_3_3790_0[1]));
    wire [1:0] far_3_3790_1;    relay_conn far_3_3790_1_a(.in(far_3_3790_0[0]), .out(far_3_3790_1[0]));    relay_conn far_3_3790_1_b(.in(far_3_3790_0[1]), .out(far_3_3790_1[1]));
    wire [1:0] far_3_3790_2;    relay_conn far_3_3790_2_a(.in(far_3_3790_1[0]), .out(far_3_3790_2[0]));    relay_conn far_3_3790_2_b(.in(far_3_3790_1[1]), .out(far_3_3790_2[1]));
    assign layer_3[730] = ~(far_3_3790_2[0] | far_3_3790_2[1]); 
    assign layer_3[731] = ~layer_2[649]; 
    wire [1:0] far_3_3792_0;    relay_conn far_3_3792_0_a(.in(layer_2[660]), .out(far_3_3792_0[0]));    relay_conn far_3_3792_0_b(.in(layer_2[573]), .out(far_3_3792_0[1]));
    wire [1:0] far_3_3792_1;    relay_conn far_3_3792_1_a(.in(far_3_3792_0[0]), .out(far_3_3792_1[0]));    relay_conn far_3_3792_1_b(.in(far_3_3792_0[1]), .out(far_3_3792_1[1]));
    assign layer_3[732] = ~(far_3_3792_1[0] & far_3_3792_1[1]); 
    wire [1:0] far_3_3793_0;    relay_conn far_3_3793_0_a(.in(layer_2[774]), .out(far_3_3793_0[0]));    relay_conn far_3_3793_0_b(.in(layer_2[651]), .out(far_3_3793_0[1]));
    wire [1:0] far_3_3793_1;    relay_conn far_3_3793_1_a(.in(far_3_3793_0[0]), .out(far_3_3793_1[0]));    relay_conn far_3_3793_1_b(.in(far_3_3793_0[1]), .out(far_3_3793_1[1]));
    wire [1:0] far_3_3793_2;    relay_conn far_3_3793_2_a(.in(far_3_3793_1[0]), .out(far_3_3793_2[0]));    relay_conn far_3_3793_2_b(.in(far_3_3793_1[1]), .out(far_3_3793_2[1]));
    assign layer_3[733] = ~(far_3_3793_2[0] & far_3_3793_2[1]); 
    wire [1:0] far_3_3794_0;    relay_conn far_3_3794_0_a(.in(layer_2[25]), .out(far_3_3794_0[0]));    relay_conn far_3_3794_0_b(.in(layer_2[126]), .out(far_3_3794_0[1]));
    wire [1:0] far_3_3794_1;    relay_conn far_3_3794_1_a(.in(far_3_3794_0[0]), .out(far_3_3794_1[0]));    relay_conn far_3_3794_1_b(.in(far_3_3794_0[1]), .out(far_3_3794_1[1]));
    wire [1:0] far_3_3794_2;    relay_conn far_3_3794_2_a(.in(far_3_3794_1[0]), .out(far_3_3794_2[0]));    relay_conn far_3_3794_2_b(.in(far_3_3794_1[1]), .out(far_3_3794_2[1]));
    assign layer_3[734] = far_3_3794_2[0] | far_3_3794_2[1]; 
    wire [1:0] far_3_3795_0;    relay_conn far_3_3795_0_a(.in(layer_2[813]), .out(far_3_3795_0[0]));    relay_conn far_3_3795_0_b(.in(layer_2[770]), .out(far_3_3795_0[1]));
    assign layer_3[735] = far_3_3795_0[0] ^ far_3_3795_0[1]; 
    wire [1:0] far_3_3796_0;    relay_conn far_3_3796_0_a(.in(layer_2[813]), .out(far_3_3796_0[0]));    relay_conn far_3_3796_0_b(.in(layer_2[845]), .out(far_3_3796_0[1]));
    assign layer_3[736] = far_3_3796_0[1]; 
    wire [1:0] far_3_3797_0;    relay_conn far_3_3797_0_a(.in(layer_2[623]), .out(far_3_3797_0[0]));    relay_conn far_3_3797_0_b(.in(layer_2[722]), .out(far_3_3797_0[1]));
    wire [1:0] far_3_3797_1;    relay_conn far_3_3797_1_a(.in(far_3_3797_0[0]), .out(far_3_3797_1[0]));    relay_conn far_3_3797_1_b(.in(far_3_3797_0[1]), .out(far_3_3797_1[1]));
    wire [1:0] far_3_3797_2;    relay_conn far_3_3797_2_a(.in(far_3_3797_1[0]), .out(far_3_3797_2[0]));    relay_conn far_3_3797_2_b(.in(far_3_3797_1[1]), .out(far_3_3797_2[1]));
    assign layer_3[737] = ~far_3_3797_2[1]; 
    wire [1:0] far_3_3798_0;    relay_conn far_3_3798_0_a(.in(layer_2[429]), .out(far_3_3798_0[0]));    relay_conn far_3_3798_0_b(.in(layer_2[350]), .out(far_3_3798_0[1]));
    wire [1:0] far_3_3798_1;    relay_conn far_3_3798_1_a(.in(far_3_3798_0[0]), .out(far_3_3798_1[0]));    relay_conn far_3_3798_1_b(.in(far_3_3798_0[1]), .out(far_3_3798_1[1]));
    assign layer_3[738] = far_3_3798_1[0]; 
    wire [1:0] far_3_3799_0;    relay_conn far_3_3799_0_a(.in(layer_2[434]), .out(far_3_3799_0[0]));    relay_conn far_3_3799_0_b(.in(layer_2[519]), .out(far_3_3799_0[1]));
    wire [1:0] far_3_3799_1;    relay_conn far_3_3799_1_a(.in(far_3_3799_0[0]), .out(far_3_3799_1[0]));    relay_conn far_3_3799_1_b(.in(far_3_3799_0[1]), .out(far_3_3799_1[1]));
    assign layer_3[739] = far_3_3799_1[0] ^ far_3_3799_1[1]; 
    assign layer_3[740] = layer_2[1012] ^ layer_2[1010]; 
    wire [1:0] far_3_3801_0;    relay_conn far_3_3801_0_a(.in(layer_2[246]), .out(far_3_3801_0[0]));    relay_conn far_3_3801_0_b(.in(layer_2[320]), .out(far_3_3801_0[1]));
    wire [1:0] far_3_3801_1;    relay_conn far_3_3801_1_a(.in(far_3_3801_0[0]), .out(far_3_3801_1[0]));    relay_conn far_3_3801_1_b(.in(far_3_3801_0[1]), .out(far_3_3801_1[1]));
    assign layer_3[741] = far_3_3801_1[0] & far_3_3801_1[1]; 
    wire [1:0] far_3_3802_0;    relay_conn far_3_3802_0_a(.in(layer_2[494]), .out(far_3_3802_0[0]));    relay_conn far_3_3802_0_b(.in(layer_2[433]), .out(far_3_3802_0[1]));
    assign layer_3[742] = ~far_3_3802_0[0] | (far_3_3802_0[0] & far_3_3802_0[1]); 
    wire [1:0] far_3_3803_0;    relay_conn far_3_3803_0_a(.in(layer_2[143]), .out(far_3_3803_0[0]));    relay_conn far_3_3803_0_b(.in(layer_2[32]), .out(far_3_3803_0[1]));
    wire [1:0] far_3_3803_1;    relay_conn far_3_3803_1_a(.in(far_3_3803_0[0]), .out(far_3_3803_1[0]));    relay_conn far_3_3803_1_b(.in(far_3_3803_0[1]), .out(far_3_3803_1[1]));
    wire [1:0] far_3_3803_2;    relay_conn far_3_3803_2_a(.in(far_3_3803_1[0]), .out(far_3_3803_2[0]));    relay_conn far_3_3803_2_b(.in(far_3_3803_1[1]), .out(far_3_3803_2[1]));
    assign layer_3[743] = ~(far_3_3803_2[0] ^ far_3_3803_2[1]); 
    assign layer_3[744] = layer_2[29] & ~layer_2[26]; 
    wire [1:0] far_3_3805_0;    relay_conn far_3_3805_0_a(.in(layer_2[159]), .out(far_3_3805_0[0]));    relay_conn far_3_3805_0_b(.in(layer_2[78]), .out(far_3_3805_0[1]));
    wire [1:0] far_3_3805_1;    relay_conn far_3_3805_1_a(.in(far_3_3805_0[0]), .out(far_3_3805_1[0]));    relay_conn far_3_3805_1_b(.in(far_3_3805_0[1]), .out(far_3_3805_1[1]));
    assign layer_3[745] = far_3_3805_1[0]; 
    assign layer_3[746] = layer_2[920] | layer_2[916]; 
    wire [1:0] far_3_3807_0;    relay_conn far_3_3807_0_a(.in(layer_2[368]), .out(far_3_3807_0[0]));    relay_conn far_3_3807_0_b(.in(layer_2[247]), .out(far_3_3807_0[1]));
    wire [1:0] far_3_3807_1;    relay_conn far_3_3807_1_a(.in(far_3_3807_0[0]), .out(far_3_3807_1[0]));    relay_conn far_3_3807_1_b(.in(far_3_3807_0[1]), .out(far_3_3807_1[1]));
    wire [1:0] far_3_3807_2;    relay_conn far_3_3807_2_a(.in(far_3_3807_1[0]), .out(far_3_3807_2[0]));    relay_conn far_3_3807_2_b(.in(far_3_3807_1[1]), .out(far_3_3807_2[1]));
    assign layer_3[747] = far_3_3807_2[1] & ~far_3_3807_2[0]; 
    wire [1:0] far_3_3808_0;    relay_conn far_3_3808_0_a(.in(layer_2[303]), .out(far_3_3808_0[0]));    relay_conn far_3_3808_0_b(.in(layer_2[205]), .out(far_3_3808_0[1]));
    wire [1:0] far_3_3808_1;    relay_conn far_3_3808_1_a(.in(far_3_3808_0[0]), .out(far_3_3808_1[0]));    relay_conn far_3_3808_1_b(.in(far_3_3808_0[1]), .out(far_3_3808_1[1]));
    wire [1:0] far_3_3808_2;    relay_conn far_3_3808_2_a(.in(far_3_3808_1[0]), .out(far_3_3808_2[0]));    relay_conn far_3_3808_2_b(.in(far_3_3808_1[1]), .out(far_3_3808_2[1]));
    assign layer_3[748] = far_3_3808_2[0] & far_3_3808_2[1]; 
    wire [1:0] far_3_3809_0;    relay_conn far_3_3809_0_a(.in(layer_2[113]), .out(far_3_3809_0[0]));    relay_conn far_3_3809_0_b(.in(layer_2[38]), .out(far_3_3809_0[1]));
    wire [1:0] far_3_3809_1;    relay_conn far_3_3809_1_a(.in(far_3_3809_0[0]), .out(far_3_3809_1[0]));    relay_conn far_3_3809_1_b(.in(far_3_3809_0[1]), .out(far_3_3809_1[1]));
    assign layer_3[749] = far_3_3809_1[0] & far_3_3809_1[1]; 
    wire [1:0] far_3_3810_0;    relay_conn far_3_3810_0_a(.in(layer_2[71]), .out(far_3_3810_0[0]));    relay_conn far_3_3810_0_b(.in(layer_2[185]), .out(far_3_3810_0[1]));
    wire [1:0] far_3_3810_1;    relay_conn far_3_3810_1_a(.in(far_3_3810_0[0]), .out(far_3_3810_1[0]));    relay_conn far_3_3810_1_b(.in(far_3_3810_0[1]), .out(far_3_3810_1[1]));
    wire [1:0] far_3_3810_2;    relay_conn far_3_3810_2_a(.in(far_3_3810_1[0]), .out(far_3_3810_2[0]));    relay_conn far_3_3810_2_b(.in(far_3_3810_1[1]), .out(far_3_3810_2[1]));
    assign layer_3[750] = far_3_3810_2[0] | far_3_3810_2[1]; 
    wire [1:0] far_3_3811_0;    relay_conn far_3_3811_0_a(.in(layer_2[264]), .out(far_3_3811_0[0]));    relay_conn far_3_3811_0_b(.in(layer_2[390]), .out(far_3_3811_0[1]));
    wire [1:0] far_3_3811_1;    relay_conn far_3_3811_1_a(.in(far_3_3811_0[0]), .out(far_3_3811_1[0]));    relay_conn far_3_3811_1_b(.in(far_3_3811_0[1]), .out(far_3_3811_1[1]));
    wire [1:0] far_3_3811_2;    relay_conn far_3_3811_2_a(.in(far_3_3811_1[0]), .out(far_3_3811_2[0]));    relay_conn far_3_3811_2_b(.in(far_3_3811_1[1]), .out(far_3_3811_2[1]));
    assign layer_3[751] = far_3_3811_2[1] & ~far_3_3811_2[0]; 
    wire [1:0] far_3_3812_0;    relay_conn far_3_3812_0_a(.in(layer_2[748]), .out(far_3_3812_0[0]));    relay_conn far_3_3812_0_b(.in(layer_2[806]), .out(far_3_3812_0[1]));
    assign layer_3[752] = ~far_3_3812_0[1] | (far_3_3812_0[0] & far_3_3812_0[1]); 
    assign layer_3[753] = ~layer_2[292]; 
    wire [1:0] far_3_3814_0;    relay_conn far_3_3814_0_a(.in(layer_2[916]), .out(far_3_3814_0[0]));    relay_conn far_3_3814_0_b(.in(layer_2[1019]), .out(far_3_3814_0[1]));
    wire [1:0] far_3_3814_1;    relay_conn far_3_3814_1_a(.in(far_3_3814_0[0]), .out(far_3_3814_1[0]));    relay_conn far_3_3814_1_b(.in(far_3_3814_0[1]), .out(far_3_3814_1[1]));
    wire [1:0] far_3_3814_2;    relay_conn far_3_3814_2_a(.in(far_3_3814_1[0]), .out(far_3_3814_2[0]));    relay_conn far_3_3814_2_b(.in(far_3_3814_1[1]), .out(far_3_3814_2[1]));
    assign layer_3[754] = ~(far_3_3814_2[0] | far_3_3814_2[1]); 
    assign layer_3[755] = layer_2[27] & ~layer_2[28]; 
    wire [1:0] far_3_3816_0;    relay_conn far_3_3816_0_a(.in(layer_2[589]), .out(far_3_3816_0[0]));    relay_conn far_3_3816_0_b(.in(layer_2[531]), .out(far_3_3816_0[1]));
    assign layer_3[756] = far_3_3816_0[0] & far_3_3816_0[1]; 
    wire [1:0] far_3_3817_0;    relay_conn far_3_3817_0_a(.in(layer_2[949]), .out(far_3_3817_0[0]));    relay_conn far_3_3817_0_b(.in(layer_2[1005]), .out(far_3_3817_0[1]));
    assign layer_3[757] = far_3_3817_0[0] & far_3_3817_0[1]; 
    wire [1:0] far_3_3818_0;    relay_conn far_3_3818_0_a(.in(layer_2[248]), .out(far_3_3818_0[0]));    relay_conn far_3_3818_0_b(.in(layer_2[283]), .out(far_3_3818_0[1]));
    assign layer_3[758] = far_3_3818_0[1]; 
    assign layer_3[759] = ~(layer_2[899] ^ layer_2[897]); 
    wire [1:0] far_3_3820_0;    relay_conn far_3_3820_0_a(.in(layer_2[276]), .out(far_3_3820_0[0]));    relay_conn far_3_3820_0_b(.in(layer_2[379]), .out(far_3_3820_0[1]));
    wire [1:0] far_3_3820_1;    relay_conn far_3_3820_1_a(.in(far_3_3820_0[0]), .out(far_3_3820_1[0]));    relay_conn far_3_3820_1_b(.in(far_3_3820_0[1]), .out(far_3_3820_1[1]));
    wire [1:0] far_3_3820_2;    relay_conn far_3_3820_2_a(.in(far_3_3820_1[0]), .out(far_3_3820_2[0]));    relay_conn far_3_3820_2_b(.in(far_3_3820_1[1]), .out(far_3_3820_2[1]));
    assign layer_3[760] = far_3_3820_2[1] & ~far_3_3820_2[0]; 
    assign layer_3[761] = layer_2[327] | layer_2[339]; 
    wire [1:0] far_3_3822_0;    relay_conn far_3_3822_0_a(.in(layer_2[57]), .out(far_3_3822_0[0]));    relay_conn far_3_3822_0_b(.in(layer_2[127]), .out(far_3_3822_0[1]));
    wire [1:0] far_3_3822_1;    relay_conn far_3_3822_1_a(.in(far_3_3822_0[0]), .out(far_3_3822_1[0]));    relay_conn far_3_3822_1_b(.in(far_3_3822_0[1]), .out(far_3_3822_1[1]));
    assign layer_3[762] = ~far_3_3822_1[0] | (far_3_3822_1[0] & far_3_3822_1[1]); 
    assign layer_3[763] = ~layer_2[90]; 
    wire [1:0] far_3_3824_0;    relay_conn far_3_3824_0_a(.in(layer_2[141]), .out(far_3_3824_0[0]));    relay_conn far_3_3824_0_b(.in(layer_2[215]), .out(far_3_3824_0[1]));
    wire [1:0] far_3_3824_1;    relay_conn far_3_3824_1_a(.in(far_3_3824_0[0]), .out(far_3_3824_1[0]));    relay_conn far_3_3824_1_b(.in(far_3_3824_0[1]), .out(far_3_3824_1[1]));
    assign layer_3[764] = ~far_3_3824_1[0] | (far_3_3824_1[0] & far_3_3824_1[1]); 
    assign layer_3[765] = ~(layer_2[232] ^ layer_2[219]); 
    wire [1:0] far_3_3826_0;    relay_conn far_3_3826_0_a(.in(layer_2[107]), .out(far_3_3826_0[0]));    relay_conn far_3_3826_0_b(.in(layer_2[196]), .out(far_3_3826_0[1]));
    wire [1:0] far_3_3826_1;    relay_conn far_3_3826_1_a(.in(far_3_3826_0[0]), .out(far_3_3826_1[0]));    relay_conn far_3_3826_1_b(.in(far_3_3826_0[1]), .out(far_3_3826_1[1]));
    assign layer_3[766] = ~far_3_3826_1[0]; 
    assign layer_3[767] = layer_2[499]; 
    assign layer_3[768] = layer_2[426] & ~layer_2[449]; 
    wire [1:0] far_3_3829_0;    relay_conn far_3_3829_0_a(.in(layer_2[418]), .out(far_3_3829_0[0]));    relay_conn far_3_3829_0_b(.in(layer_2[335]), .out(far_3_3829_0[1]));
    wire [1:0] far_3_3829_1;    relay_conn far_3_3829_1_a(.in(far_3_3829_0[0]), .out(far_3_3829_1[0]));    relay_conn far_3_3829_1_b(.in(far_3_3829_0[1]), .out(far_3_3829_1[1]));
    assign layer_3[769] = far_3_3829_1[1] & ~far_3_3829_1[0]; 
    wire [1:0] far_3_3830_0;    relay_conn far_3_3830_0_a(.in(layer_2[450]), .out(far_3_3830_0[0]));    relay_conn far_3_3830_0_b(.in(layer_2[539]), .out(far_3_3830_0[1]));
    wire [1:0] far_3_3830_1;    relay_conn far_3_3830_1_a(.in(far_3_3830_0[0]), .out(far_3_3830_1[0]));    relay_conn far_3_3830_1_b(.in(far_3_3830_0[1]), .out(far_3_3830_1[1]));
    assign layer_3[770] = ~far_3_3830_1[1] | (far_3_3830_1[0] & far_3_3830_1[1]); 
    assign layer_3[771] = ~layer_2[32] | (layer_2[32] & layer_2[57]); 
    wire [1:0] far_3_3832_0;    relay_conn far_3_3832_0_a(.in(layer_2[191]), .out(far_3_3832_0[0]));    relay_conn far_3_3832_0_b(.in(layer_2[79]), .out(far_3_3832_0[1]));
    wire [1:0] far_3_3832_1;    relay_conn far_3_3832_1_a(.in(far_3_3832_0[0]), .out(far_3_3832_1[0]));    relay_conn far_3_3832_1_b(.in(far_3_3832_0[1]), .out(far_3_3832_1[1]));
    wire [1:0] far_3_3832_2;    relay_conn far_3_3832_2_a(.in(far_3_3832_1[0]), .out(far_3_3832_2[0]));    relay_conn far_3_3832_2_b(.in(far_3_3832_1[1]), .out(far_3_3832_2[1]));
    assign layer_3[772] = ~far_3_3832_2[0] | (far_3_3832_2[0] & far_3_3832_2[1]); 
    assign layer_3[773] = ~layer_2[837]; 
    wire [1:0] far_3_3834_0;    relay_conn far_3_3834_0_a(.in(layer_2[542]), .out(far_3_3834_0[0]));    relay_conn far_3_3834_0_b(.in(layer_2[477]), .out(far_3_3834_0[1]));
    wire [1:0] far_3_3834_1;    relay_conn far_3_3834_1_a(.in(far_3_3834_0[0]), .out(far_3_3834_1[0]));    relay_conn far_3_3834_1_b(.in(far_3_3834_0[1]), .out(far_3_3834_1[1]));
    assign layer_3[774] = far_3_3834_1[1]; 
    wire [1:0] far_3_3835_0;    relay_conn far_3_3835_0_a(.in(layer_2[826]), .out(far_3_3835_0[0]));    relay_conn far_3_3835_0_b(.in(layer_2[902]), .out(far_3_3835_0[1]));
    wire [1:0] far_3_3835_1;    relay_conn far_3_3835_1_a(.in(far_3_3835_0[0]), .out(far_3_3835_1[0]));    relay_conn far_3_3835_1_b(.in(far_3_3835_0[1]), .out(far_3_3835_1[1]));
    assign layer_3[775] = far_3_3835_1[0] ^ far_3_3835_1[1]; 
    assign layer_3[776] = ~(layer_2[840] ^ layer_2[824]); 
    wire [1:0] far_3_3837_0;    relay_conn far_3_3837_0_a(.in(layer_2[350]), .out(far_3_3837_0[0]));    relay_conn far_3_3837_0_b(.in(layer_2[388]), .out(far_3_3837_0[1]));
    assign layer_3[777] = far_3_3837_0[0] & far_3_3837_0[1]; 
    wire [1:0] far_3_3838_0;    relay_conn far_3_3838_0_a(.in(layer_2[341]), .out(far_3_3838_0[0]));    relay_conn far_3_3838_0_b(.in(layer_2[460]), .out(far_3_3838_0[1]));
    wire [1:0] far_3_3838_1;    relay_conn far_3_3838_1_a(.in(far_3_3838_0[0]), .out(far_3_3838_1[0]));    relay_conn far_3_3838_1_b(.in(far_3_3838_0[1]), .out(far_3_3838_1[1]));
    wire [1:0] far_3_3838_2;    relay_conn far_3_3838_2_a(.in(far_3_3838_1[0]), .out(far_3_3838_2[0]));    relay_conn far_3_3838_2_b(.in(far_3_3838_1[1]), .out(far_3_3838_2[1]));
    assign layer_3[778] = far_3_3838_2[0] & far_3_3838_2[1]; 
    assign layer_3[779] = ~(layer_2[550] | layer_2[578]); 
    assign layer_3[780] = ~layer_2[126] | (layer_2[126] & layer_2[148]); 
    wire [1:0] far_3_3841_0;    relay_conn far_3_3841_0_a(.in(layer_2[246]), .out(far_3_3841_0[0]));    relay_conn far_3_3841_0_b(.in(layer_2[130]), .out(far_3_3841_0[1]));
    wire [1:0] far_3_3841_1;    relay_conn far_3_3841_1_a(.in(far_3_3841_0[0]), .out(far_3_3841_1[0]));    relay_conn far_3_3841_1_b(.in(far_3_3841_0[1]), .out(far_3_3841_1[1]));
    wire [1:0] far_3_3841_2;    relay_conn far_3_3841_2_a(.in(far_3_3841_1[0]), .out(far_3_3841_2[0]));    relay_conn far_3_3841_2_b(.in(far_3_3841_1[1]), .out(far_3_3841_2[1]));
    assign layer_3[781] = ~far_3_3841_2[0] | (far_3_3841_2[0] & far_3_3841_2[1]); 
    wire [1:0] far_3_3842_0;    relay_conn far_3_3842_0_a(.in(layer_2[265]), .out(far_3_3842_0[0]));    relay_conn far_3_3842_0_b(.in(layer_2[345]), .out(far_3_3842_0[1]));
    wire [1:0] far_3_3842_1;    relay_conn far_3_3842_1_a(.in(far_3_3842_0[0]), .out(far_3_3842_1[0]));    relay_conn far_3_3842_1_b(.in(far_3_3842_0[1]), .out(far_3_3842_1[1]));
    assign layer_3[782] = far_3_3842_1[1]; 
    assign layer_3[783] = ~(layer_2[100] & layer_2[107]); 
    assign layer_3[784] = layer_2[1005]; 
    wire [1:0] far_3_3845_0;    relay_conn far_3_3845_0_a(.in(layer_2[24]), .out(far_3_3845_0[0]));    relay_conn far_3_3845_0_b(.in(layer_2[141]), .out(far_3_3845_0[1]));
    wire [1:0] far_3_3845_1;    relay_conn far_3_3845_1_a(.in(far_3_3845_0[0]), .out(far_3_3845_1[0]));    relay_conn far_3_3845_1_b(.in(far_3_3845_0[1]), .out(far_3_3845_1[1]));
    wire [1:0] far_3_3845_2;    relay_conn far_3_3845_2_a(.in(far_3_3845_1[0]), .out(far_3_3845_2[0]));    relay_conn far_3_3845_2_b(.in(far_3_3845_1[1]), .out(far_3_3845_2[1]));
    assign layer_3[785] = far_3_3845_2[1] & ~far_3_3845_2[0]; 
    wire [1:0] far_3_3846_0;    relay_conn far_3_3846_0_a(.in(layer_2[542]), .out(far_3_3846_0[0]));    relay_conn far_3_3846_0_b(.in(layer_2[421]), .out(far_3_3846_0[1]));
    wire [1:0] far_3_3846_1;    relay_conn far_3_3846_1_a(.in(far_3_3846_0[0]), .out(far_3_3846_1[0]));    relay_conn far_3_3846_1_b(.in(far_3_3846_0[1]), .out(far_3_3846_1[1]));
    wire [1:0] far_3_3846_2;    relay_conn far_3_3846_2_a(.in(far_3_3846_1[0]), .out(far_3_3846_2[0]));    relay_conn far_3_3846_2_b(.in(far_3_3846_1[1]), .out(far_3_3846_2[1]));
    assign layer_3[786] = ~(far_3_3846_2[0] | far_3_3846_2[1]); 
    wire [1:0] far_3_3847_0;    relay_conn far_3_3847_0_a(.in(layer_2[155]), .out(far_3_3847_0[0]));    relay_conn far_3_3847_0_b(.in(layer_2[94]), .out(far_3_3847_0[1]));
    assign layer_3[787] = ~far_3_3847_0[1] | (far_3_3847_0[0] & far_3_3847_0[1]); 
    wire [1:0] far_3_3848_0;    relay_conn far_3_3848_0_a(.in(layer_2[323]), .out(far_3_3848_0[0]));    relay_conn far_3_3848_0_b(.in(layer_2[442]), .out(far_3_3848_0[1]));
    wire [1:0] far_3_3848_1;    relay_conn far_3_3848_1_a(.in(far_3_3848_0[0]), .out(far_3_3848_1[0]));    relay_conn far_3_3848_1_b(.in(far_3_3848_0[1]), .out(far_3_3848_1[1]));
    wire [1:0] far_3_3848_2;    relay_conn far_3_3848_2_a(.in(far_3_3848_1[0]), .out(far_3_3848_2[0]));    relay_conn far_3_3848_2_b(.in(far_3_3848_1[1]), .out(far_3_3848_2[1]));
    assign layer_3[788] = ~far_3_3848_2[1] | (far_3_3848_2[0] & far_3_3848_2[1]); 
    assign layer_3[789] = ~(layer_2[626] ^ layer_2[640]); 
    wire [1:0] far_3_3850_0;    relay_conn far_3_3850_0_a(.in(layer_2[526]), .out(far_3_3850_0[0]));    relay_conn far_3_3850_0_b(.in(layer_2[644]), .out(far_3_3850_0[1]));
    wire [1:0] far_3_3850_1;    relay_conn far_3_3850_1_a(.in(far_3_3850_0[0]), .out(far_3_3850_1[0]));    relay_conn far_3_3850_1_b(.in(far_3_3850_0[1]), .out(far_3_3850_1[1]));
    wire [1:0] far_3_3850_2;    relay_conn far_3_3850_2_a(.in(far_3_3850_1[0]), .out(far_3_3850_2[0]));    relay_conn far_3_3850_2_b(.in(far_3_3850_1[1]), .out(far_3_3850_2[1]));
    assign layer_3[790] = ~far_3_3850_2[0] | (far_3_3850_2[0] & far_3_3850_2[1]); 
    assign layer_3[791] = ~layer_2[180] | (layer_2[208] & layer_2[180]); 
    assign layer_3[792] = layer_2[892] & ~layer_2[891]; 
    wire [1:0] far_3_3853_0;    relay_conn far_3_3853_0_a(.in(layer_2[925]), .out(far_3_3853_0[0]));    relay_conn far_3_3853_0_b(.in(layer_2[970]), .out(far_3_3853_0[1]));
    assign layer_3[793] = far_3_3853_0[0] & ~far_3_3853_0[1]; 
    wire [1:0] far_3_3854_0;    relay_conn far_3_3854_0_a(.in(layer_2[663]), .out(far_3_3854_0[0]));    relay_conn far_3_3854_0_b(.in(layer_2[775]), .out(far_3_3854_0[1]));
    wire [1:0] far_3_3854_1;    relay_conn far_3_3854_1_a(.in(far_3_3854_0[0]), .out(far_3_3854_1[0]));    relay_conn far_3_3854_1_b(.in(far_3_3854_0[1]), .out(far_3_3854_1[1]));
    wire [1:0] far_3_3854_2;    relay_conn far_3_3854_2_a(.in(far_3_3854_1[0]), .out(far_3_3854_2[0]));    relay_conn far_3_3854_2_b(.in(far_3_3854_1[1]), .out(far_3_3854_2[1]));
    assign layer_3[794] = ~far_3_3854_2[1] | (far_3_3854_2[0] & far_3_3854_2[1]); 
    wire [1:0] far_3_3855_0;    relay_conn far_3_3855_0_a(.in(layer_2[798]), .out(far_3_3855_0[0]));    relay_conn far_3_3855_0_b(.in(layer_2[726]), .out(far_3_3855_0[1]));
    wire [1:0] far_3_3855_1;    relay_conn far_3_3855_1_a(.in(far_3_3855_0[0]), .out(far_3_3855_1[0]));    relay_conn far_3_3855_1_b(.in(far_3_3855_0[1]), .out(far_3_3855_1[1]));
    assign layer_3[795] = ~far_3_3855_1[0]; 
    wire [1:0] far_3_3856_0;    relay_conn far_3_3856_0_a(.in(layer_2[255]), .out(far_3_3856_0[0]));    relay_conn far_3_3856_0_b(.in(layer_2[383]), .out(far_3_3856_0[1]));
    wire [1:0] far_3_3856_1;    relay_conn far_3_3856_1_a(.in(far_3_3856_0[0]), .out(far_3_3856_1[0]));    relay_conn far_3_3856_1_b(.in(far_3_3856_0[1]), .out(far_3_3856_1[1]));
    wire [1:0] far_3_3856_2;    relay_conn far_3_3856_2_a(.in(far_3_3856_1[0]), .out(far_3_3856_2[0]));    relay_conn far_3_3856_2_b(.in(far_3_3856_1[1]), .out(far_3_3856_2[1]));
    wire [1:0] far_3_3856_3;    relay_conn far_3_3856_3_a(.in(far_3_3856_2[0]), .out(far_3_3856_3[0]));    relay_conn far_3_3856_3_b(.in(far_3_3856_2[1]), .out(far_3_3856_3[1]));
    assign layer_3[796] = far_3_3856_3[0] & far_3_3856_3[1]; 
    wire [1:0] far_3_3857_0;    relay_conn far_3_3857_0_a(.in(layer_2[721]), .out(far_3_3857_0[0]));    relay_conn far_3_3857_0_b(.in(layer_2[823]), .out(far_3_3857_0[1]));
    wire [1:0] far_3_3857_1;    relay_conn far_3_3857_1_a(.in(far_3_3857_0[0]), .out(far_3_3857_1[0]));    relay_conn far_3_3857_1_b(.in(far_3_3857_0[1]), .out(far_3_3857_1[1]));
    wire [1:0] far_3_3857_2;    relay_conn far_3_3857_2_a(.in(far_3_3857_1[0]), .out(far_3_3857_2[0]));    relay_conn far_3_3857_2_b(.in(far_3_3857_1[1]), .out(far_3_3857_2[1]));
    assign layer_3[797] = far_3_3857_2[0] & far_3_3857_2[1]; 
    wire [1:0] far_3_3858_0;    relay_conn far_3_3858_0_a(.in(layer_2[766]), .out(far_3_3858_0[0]));    relay_conn far_3_3858_0_b(.in(layer_2[663]), .out(far_3_3858_0[1]));
    wire [1:0] far_3_3858_1;    relay_conn far_3_3858_1_a(.in(far_3_3858_0[0]), .out(far_3_3858_1[0]));    relay_conn far_3_3858_1_b(.in(far_3_3858_0[1]), .out(far_3_3858_1[1]));
    wire [1:0] far_3_3858_2;    relay_conn far_3_3858_2_a(.in(far_3_3858_1[0]), .out(far_3_3858_2[0]));    relay_conn far_3_3858_2_b(.in(far_3_3858_1[1]), .out(far_3_3858_2[1]));
    assign layer_3[798] = far_3_3858_2[1]; 
    wire [1:0] far_3_3859_0;    relay_conn far_3_3859_0_a(.in(layer_2[559]), .out(far_3_3859_0[0]));    relay_conn far_3_3859_0_b(.in(layer_2[480]), .out(far_3_3859_0[1]));
    wire [1:0] far_3_3859_1;    relay_conn far_3_3859_1_a(.in(far_3_3859_0[0]), .out(far_3_3859_1[0]));    relay_conn far_3_3859_1_b(.in(far_3_3859_0[1]), .out(far_3_3859_1[1]));
    assign layer_3[799] = far_3_3859_1[0] & far_3_3859_1[1]; 
    wire [1:0] far_3_3860_0;    relay_conn far_3_3860_0_a(.in(layer_2[852]), .out(far_3_3860_0[0]));    relay_conn far_3_3860_0_b(.in(layer_2[763]), .out(far_3_3860_0[1]));
    wire [1:0] far_3_3860_1;    relay_conn far_3_3860_1_a(.in(far_3_3860_0[0]), .out(far_3_3860_1[0]));    relay_conn far_3_3860_1_b(.in(far_3_3860_0[1]), .out(far_3_3860_1[1]));
    assign layer_3[800] = ~far_3_3860_1[0] | (far_3_3860_1[0] & far_3_3860_1[1]); 
    wire [1:0] far_3_3861_0;    relay_conn far_3_3861_0_a(.in(layer_2[64]), .out(far_3_3861_0[0]));    relay_conn far_3_3861_0_b(.in(layer_2[188]), .out(far_3_3861_0[1]));
    wire [1:0] far_3_3861_1;    relay_conn far_3_3861_1_a(.in(far_3_3861_0[0]), .out(far_3_3861_1[0]));    relay_conn far_3_3861_1_b(.in(far_3_3861_0[1]), .out(far_3_3861_1[1]));
    wire [1:0] far_3_3861_2;    relay_conn far_3_3861_2_a(.in(far_3_3861_1[0]), .out(far_3_3861_2[0]));    relay_conn far_3_3861_2_b(.in(far_3_3861_1[1]), .out(far_3_3861_2[1]));
    assign layer_3[801] = far_3_3861_2[1] & ~far_3_3861_2[0]; 
    assign layer_3[802] = layer_2[1016] & layer_2[986]; 
    wire [1:0] far_3_3863_0;    relay_conn far_3_3863_0_a(.in(layer_2[141]), .out(far_3_3863_0[0]));    relay_conn far_3_3863_0_b(.in(layer_2[266]), .out(far_3_3863_0[1]));
    wire [1:0] far_3_3863_1;    relay_conn far_3_3863_1_a(.in(far_3_3863_0[0]), .out(far_3_3863_1[0]));    relay_conn far_3_3863_1_b(.in(far_3_3863_0[1]), .out(far_3_3863_1[1]));
    wire [1:0] far_3_3863_2;    relay_conn far_3_3863_2_a(.in(far_3_3863_1[0]), .out(far_3_3863_2[0]));    relay_conn far_3_3863_2_b(.in(far_3_3863_1[1]), .out(far_3_3863_2[1]));
    assign layer_3[803] = far_3_3863_2[0]; 
    wire [1:0] far_3_3864_0;    relay_conn far_3_3864_0_a(.in(layer_2[333]), .out(far_3_3864_0[0]));    relay_conn far_3_3864_0_b(.in(layer_2[208]), .out(far_3_3864_0[1]));
    wire [1:0] far_3_3864_1;    relay_conn far_3_3864_1_a(.in(far_3_3864_0[0]), .out(far_3_3864_1[0]));    relay_conn far_3_3864_1_b(.in(far_3_3864_0[1]), .out(far_3_3864_1[1]));
    wire [1:0] far_3_3864_2;    relay_conn far_3_3864_2_a(.in(far_3_3864_1[0]), .out(far_3_3864_2[0]));    relay_conn far_3_3864_2_b(.in(far_3_3864_1[1]), .out(far_3_3864_2[1]));
    assign layer_3[804] = far_3_3864_2[0]; 
    assign layer_3[805] = ~layer_2[218] | (layer_2[241] & layer_2[218]); 
    wire [1:0] far_3_3866_0;    relay_conn far_3_3866_0_a(.in(layer_2[946]), .out(far_3_3866_0[0]));    relay_conn far_3_3866_0_b(.in(layer_2[899]), .out(far_3_3866_0[1]));
    assign layer_3[806] = ~far_3_3866_0[1]; 
    wire [1:0] far_3_3867_0;    relay_conn far_3_3867_0_a(.in(layer_2[993]), .out(far_3_3867_0[0]));    relay_conn far_3_3867_0_b(.in(layer_2[915]), .out(far_3_3867_0[1]));
    wire [1:0] far_3_3867_1;    relay_conn far_3_3867_1_a(.in(far_3_3867_0[0]), .out(far_3_3867_1[0]));    relay_conn far_3_3867_1_b(.in(far_3_3867_0[1]), .out(far_3_3867_1[1]));
    assign layer_3[807] = far_3_3867_1[0]; 
    wire [1:0] far_3_3868_0;    relay_conn far_3_3868_0_a(.in(layer_2[859]), .out(far_3_3868_0[0]));    relay_conn far_3_3868_0_b(.in(layer_2[952]), .out(far_3_3868_0[1]));
    wire [1:0] far_3_3868_1;    relay_conn far_3_3868_1_a(.in(far_3_3868_0[0]), .out(far_3_3868_1[0]));    relay_conn far_3_3868_1_b(.in(far_3_3868_0[1]), .out(far_3_3868_1[1]));
    assign layer_3[808] = ~far_3_3868_1[1] | (far_3_3868_1[0] & far_3_3868_1[1]); 
    wire [1:0] far_3_3869_0;    relay_conn far_3_3869_0_a(.in(layer_2[340]), .out(far_3_3869_0[0]));    relay_conn far_3_3869_0_b(.in(layer_2[301]), .out(far_3_3869_0[1]));
    assign layer_3[809] = far_3_3869_0[1] & ~far_3_3869_0[0]; 
    assign layer_3[810] = layer_2[558]; 
    wire [1:0] far_3_3871_0;    relay_conn far_3_3871_0_a(.in(layer_2[960]), .out(far_3_3871_0[0]));    relay_conn far_3_3871_0_b(.in(layer_2[872]), .out(far_3_3871_0[1]));
    wire [1:0] far_3_3871_1;    relay_conn far_3_3871_1_a(.in(far_3_3871_0[0]), .out(far_3_3871_1[0]));    relay_conn far_3_3871_1_b(.in(far_3_3871_0[1]), .out(far_3_3871_1[1]));
    assign layer_3[811] = far_3_3871_1[0] ^ far_3_3871_1[1]; 
    wire [1:0] far_3_3872_0;    relay_conn far_3_3872_0_a(.in(layer_2[363]), .out(far_3_3872_0[0]));    relay_conn far_3_3872_0_b(.in(layer_2[245]), .out(far_3_3872_0[1]));
    wire [1:0] far_3_3872_1;    relay_conn far_3_3872_1_a(.in(far_3_3872_0[0]), .out(far_3_3872_1[0]));    relay_conn far_3_3872_1_b(.in(far_3_3872_0[1]), .out(far_3_3872_1[1]));
    wire [1:0] far_3_3872_2;    relay_conn far_3_3872_2_a(.in(far_3_3872_1[0]), .out(far_3_3872_2[0]));    relay_conn far_3_3872_2_b(.in(far_3_3872_1[1]), .out(far_3_3872_2[1]));
    assign layer_3[812] = far_3_3872_2[1] & ~far_3_3872_2[0]; 
    assign layer_3[813] = layer_2[262]; 
    wire [1:0] far_3_3874_0;    relay_conn far_3_3874_0_a(.in(layer_2[424]), .out(far_3_3874_0[0]));    relay_conn far_3_3874_0_b(.in(layer_2[516]), .out(far_3_3874_0[1]));
    wire [1:0] far_3_3874_1;    relay_conn far_3_3874_1_a(.in(far_3_3874_0[0]), .out(far_3_3874_1[0]));    relay_conn far_3_3874_1_b(.in(far_3_3874_0[1]), .out(far_3_3874_1[1]));
    assign layer_3[814] = ~(far_3_3874_1[0] | far_3_3874_1[1]); 
    assign layer_3[815] = ~layer_2[120] | (layer_2[120] & layer_2[151]); 
    wire [1:0] far_3_3876_0;    relay_conn far_3_3876_0_a(.in(layer_2[87]), .out(far_3_3876_0[0]));    relay_conn far_3_3876_0_b(.in(layer_2[191]), .out(far_3_3876_0[1]));
    wire [1:0] far_3_3876_1;    relay_conn far_3_3876_1_a(.in(far_3_3876_0[0]), .out(far_3_3876_1[0]));    relay_conn far_3_3876_1_b(.in(far_3_3876_0[1]), .out(far_3_3876_1[1]));
    wire [1:0] far_3_3876_2;    relay_conn far_3_3876_2_a(.in(far_3_3876_1[0]), .out(far_3_3876_2[0]));    relay_conn far_3_3876_2_b(.in(far_3_3876_1[1]), .out(far_3_3876_2[1]));
    assign layer_3[816] = ~(far_3_3876_2[0] ^ far_3_3876_2[1]); 
    wire [1:0] far_3_3877_0;    relay_conn far_3_3877_0_a(.in(layer_2[671]), .out(far_3_3877_0[0]));    relay_conn far_3_3877_0_b(.in(layer_2[785]), .out(far_3_3877_0[1]));
    wire [1:0] far_3_3877_1;    relay_conn far_3_3877_1_a(.in(far_3_3877_0[0]), .out(far_3_3877_1[0]));    relay_conn far_3_3877_1_b(.in(far_3_3877_0[1]), .out(far_3_3877_1[1]));
    wire [1:0] far_3_3877_2;    relay_conn far_3_3877_2_a(.in(far_3_3877_1[0]), .out(far_3_3877_2[0]));    relay_conn far_3_3877_2_b(.in(far_3_3877_1[1]), .out(far_3_3877_2[1]));
    assign layer_3[817] = far_3_3877_2[0] & ~far_3_3877_2[1]; 
    wire [1:0] far_3_3878_0;    relay_conn far_3_3878_0_a(.in(layer_2[164]), .out(far_3_3878_0[0]));    relay_conn far_3_3878_0_b(.in(layer_2[235]), .out(far_3_3878_0[1]));
    wire [1:0] far_3_3878_1;    relay_conn far_3_3878_1_a(.in(far_3_3878_0[0]), .out(far_3_3878_1[0]));    relay_conn far_3_3878_1_b(.in(far_3_3878_0[1]), .out(far_3_3878_1[1]));
    assign layer_3[818] = ~(far_3_3878_1[0] | far_3_3878_1[1]); 
    assign layer_3[819] = layer_2[926]; 
    wire [1:0] far_3_3880_0;    relay_conn far_3_3880_0_a(.in(layer_2[205]), .out(far_3_3880_0[0]));    relay_conn far_3_3880_0_b(.in(layer_2[327]), .out(far_3_3880_0[1]));
    wire [1:0] far_3_3880_1;    relay_conn far_3_3880_1_a(.in(far_3_3880_0[0]), .out(far_3_3880_1[0]));    relay_conn far_3_3880_1_b(.in(far_3_3880_0[1]), .out(far_3_3880_1[1]));
    wire [1:0] far_3_3880_2;    relay_conn far_3_3880_2_a(.in(far_3_3880_1[0]), .out(far_3_3880_2[0]));    relay_conn far_3_3880_2_b(.in(far_3_3880_1[1]), .out(far_3_3880_2[1]));
    assign layer_3[820] = ~far_3_3880_2[1]; 
    wire [1:0] far_3_3881_0;    relay_conn far_3_3881_0_a(.in(layer_2[796]), .out(far_3_3881_0[0]));    relay_conn far_3_3881_0_b(.in(layer_2[842]), .out(far_3_3881_0[1]));
    assign layer_3[821] = ~far_3_3881_0[1] | (far_3_3881_0[0] & far_3_3881_0[1]); 
    wire [1:0] far_3_3882_0;    relay_conn far_3_3882_0_a(.in(layer_2[429]), .out(far_3_3882_0[0]));    relay_conn far_3_3882_0_b(.in(layer_2[548]), .out(far_3_3882_0[1]));
    wire [1:0] far_3_3882_1;    relay_conn far_3_3882_1_a(.in(far_3_3882_0[0]), .out(far_3_3882_1[0]));    relay_conn far_3_3882_1_b(.in(far_3_3882_0[1]), .out(far_3_3882_1[1]));
    wire [1:0] far_3_3882_2;    relay_conn far_3_3882_2_a(.in(far_3_3882_1[0]), .out(far_3_3882_2[0]));    relay_conn far_3_3882_2_b(.in(far_3_3882_1[1]), .out(far_3_3882_2[1]));
    assign layer_3[822] = ~far_3_3882_2[0] | (far_3_3882_2[0] & far_3_3882_2[1]); 
    wire [1:0] far_3_3883_0;    relay_conn far_3_3883_0_a(.in(layer_2[302]), .out(far_3_3883_0[0]));    relay_conn far_3_3883_0_b(.in(layer_2[252]), .out(far_3_3883_0[1]));
    assign layer_3[823] = ~(far_3_3883_0[0] & far_3_3883_0[1]); 
    wire [1:0] far_3_3884_0;    relay_conn far_3_3884_0_a(.in(layer_2[621]), .out(far_3_3884_0[0]));    relay_conn far_3_3884_0_b(.in(layer_2[585]), .out(far_3_3884_0[1]));
    assign layer_3[824] = far_3_3884_0[1]; 
    wire [1:0] far_3_3885_0;    relay_conn far_3_3885_0_a(.in(layer_2[208]), .out(far_3_3885_0[0]));    relay_conn far_3_3885_0_b(.in(layer_2[277]), .out(far_3_3885_0[1]));
    wire [1:0] far_3_3885_1;    relay_conn far_3_3885_1_a(.in(far_3_3885_0[0]), .out(far_3_3885_1[0]));    relay_conn far_3_3885_1_b(.in(far_3_3885_0[1]), .out(far_3_3885_1[1]));
    assign layer_3[825] = ~far_3_3885_1[1]; 
    wire [1:0] far_3_3886_0;    relay_conn far_3_3886_0_a(.in(layer_2[543]), .out(far_3_3886_0[0]));    relay_conn far_3_3886_0_b(.in(layer_2[612]), .out(far_3_3886_0[1]));
    wire [1:0] far_3_3886_1;    relay_conn far_3_3886_1_a(.in(far_3_3886_0[0]), .out(far_3_3886_1[0]));    relay_conn far_3_3886_1_b(.in(far_3_3886_0[1]), .out(far_3_3886_1[1]));
    assign layer_3[826] = far_3_3886_1[0] & ~far_3_3886_1[1]; 
    assign layer_3[827] = ~layer_2[913] | (layer_2[913] & layer_2[927]); 
    wire [1:0] far_3_3888_0;    relay_conn far_3_3888_0_a(.in(layer_2[674]), .out(far_3_3888_0[0]));    relay_conn far_3_3888_0_b(.in(layer_2[762]), .out(far_3_3888_0[1]));
    wire [1:0] far_3_3888_1;    relay_conn far_3_3888_1_a(.in(far_3_3888_0[0]), .out(far_3_3888_1[0]));    relay_conn far_3_3888_1_b(.in(far_3_3888_0[1]), .out(far_3_3888_1[1]));
    assign layer_3[828] = far_3_3888_1[0] & far_3_3888_1[1]; 
    wire [1:0] far_3_3889_0;    relay_conn far_3_3889_0_a(.in(layer_2[200]), .out(far_3_3889_0[0]));    relay_conn far_3_3889_0_b(.in(layer_2[112]), .out(far_3_3889_0[1]));
    wire [1:0] far_3_3889_1;    relay_conn far_3_3889_1_a(.in(far_3_3889_0[0]), .out(far_3_3889_1[0]));    relay_conn far_3_3889_1_b(.in(far_3_3889_0[1]), .out(far_3_3889_1[1]));
    assign layer_3[829] = far_3_3889_1[0] | far_3_3889_1[1]; 
    wire [1:0] far_3_3890_0;    relay_conn far_3_3890_0_a(.in(layer_2[106]), .out(far_3_3890_0[0]));    relay_conn far_3_3890_0_b(.in(layer_2[1]), .out(far_3_3890_0[1]));
    wire [1:0] far_3_3890_1;    relay_conn far_3_3890_1_a(.in(far_3_3890_0[0]), .out(far_3_3890_1[0]));    relay_conn far_3_3890_1_b(.in(far_3_3890_0[1]), .out(far_3_3890_1[1]));
    wire [1:0] far_3_3890_2;    relay_conn far_3_3890_2_a(.in(far_3_3890_1[0]), .out(far_3_3890_2[0]));    relay_conn far_3_3890_2_b(.in(far_3_3890_1[1]), .out(far_3_3890_2[1]));
    assign layer_3[830] = far_3_3890_2[0] & ~far_3_3890_2[1]; 
    wire [1:0] far_3_3891_0;    relay_conn far_3_3891_0_a(.in(layer_2[3]), .out(far_3_3891_0[0]));    relay_conn far_3_3891_0_b(.in(layer_2[100]), .out(far_3_3891_0[1]));
    wire [1:0] far_3_3891_1;    relay_conn far_3_3891_1_a(.in(far_3_3891_0[0]), .out(far_3_3891_1[0]));    relay_conn far_3_3891_1_b(.in(far_3_3891_0[1]), .out(far_3_3891_1[1]));
    wire [1:0] far_3_3891_2;    relay_conn far_3_3891_2_a(.in(far_3_3891_1[0]), .out(far_3_3891_2[0]));    relay_conn far_3_3891_2_b(.in(far_3_3891_1[1]), .out(far_3_3891_2[1]));
    assign layer_3[831] = ~(far_3_3891_2[0] & far_3_3891_2[1]); 
    assign layer_3[832] = ~layer_2[244]; 
    wire [1:0] far_3_3893_0;    relay_conn far_3_3893_0_a(.in(layer_2[483]), .out(far_3_3893_0[0]));    relay_conn far_3_3893_0_b(.in(layer_2[577]), .out(far_3_3893_0[1]));
    wire [1:0] far_3_3893_1;    relay_conn far_3_3893_1_a(.in(far_3_3893_0[0]), .out(far_3_3893_1[0]));    relay_conn far_3_3893_1_b(.in(far_3_3893_0[1]), .out(far_3_3893_1[1]));
    assign layer_3[833] = far_3_3893_1[0] & ~far_3_3893_1[1]; 
    assign layer_3[834] = layer_2[151]; 
    wire [1:0] far_3_3895_0;    relay_conn far_3_3895_0_a(.in(layer_2[79]), .out(far_3_3895_0[0]));    relay_conn far_3_3895_0_b(.in(layer_2[140]), .out(far_3_3895_0[1]));
    assign layer_3[835] = far_3_3895_0[1] & ~far_3_3895_0[0]; 
    assign layer_3[836] = ~layer_2[307] | (layer_2[310] & layer_2[307]); 
    wire [1:0] far_3_3897_0;    relay_conn far_3_3897_0_a(.in(layer_2[725]), .out(far_3_3897_0[0]));    relay_conn far_3_3897_0_b(.in(layer_2[645]), .out(far_3_3897_0[1]));
    wire [1:0] far_3_3897_1;    relay_conn far_3_3897_1_a(.in(far_3_3897_0[0]), .out(far_3_3897_1[0]));    relay_conn far_3_3897_1_b(.in(far_3_3897_0[1]), .out(far_3_3897_1[1]));
    assign layer_3[837] = far_3_3897_1[1] & ~far_3_3897_1[0]; 
    wire [1:0] far_3_3898_0;    relay_conn far_3_3898_0_a(.in(layer_2[208]), .out(far_3_3898_0[0]));    relay_conn far_3_3898_0_b(.in(layer_2[306]), .out(far_3_3898_0[1]));
    wire [1:0] far_3_3898_1;    relay_conn far_3_3898_1_a(.in(far_3_3898_0[0]), .out(far_3_3898_1[0]));    relay_conn far_3_3898_1_b(.in(far_3_3898_0[1]), .out(far_3_3898_1[1]));
    wire [1:0] far_3_3898_2;    relay_conn far_3_3898_2_a(.in(far_3_3898_1[0]), .out(far_3_3898_2[0]));    relay_conn far_3_3898_2_b(.in(far_3_3898_1[1]), .out(far_3_3898_2[1]));
    assign layer_3[838] = far_3_3898_2[1] & ~far_3_3898_2[0]; 
    assign layer_3[839] = layer_2[798] & ~layer_2[780]; 
    wire [1:0] far_3_3900_0;    relay_conn far_3_3900_0_a(.in(layer_2[79]), .out(far_3_3900_0[0]));    relay_conn far_3_3900_0_b(.in(layer_2[198]), .out(far_3_3900_0[1]));
    wire [1:0] far_3_3900_1;    relay_conn far_3_3900_1_a(.in(far_3_3900_0[0]), .out(far_3_3900_1[0]));    relay_conn far_3_3900_1_b(.in(far_3_3900_0[1]), .out(far_3_3900_1[1]));
    wire [1:0] far_3_3900_2;    relay_conn far_3_3900_2_a(.in(far_3_3900_1[0]), .out(far_3_3900_2[0]));    relay_conn far_3_3900_2_b(.in(far_3_3900_1[1]), .out(far_3_3900_2[1]));
    assign layer_3[840] = ~far_3_3900_2[1] | (far_3_3900_2[0] & far_3_3900_2[1]); 
    wire [1:0] far_3_3901_0;    relay_conn far_3_3901_0_a(.in(layer_2[265]), .out(far_3_3901_0[0]));    relay_conn far_3_3901_0_b(.in(layer_2[345]), .out(far_3_3901_0[1]));
    wire [1:0] far_3_3901_1;    relay_conn far_3_3901_1_a(.in(far_3_3901_0[0]), .out(far_3_3901_1[0]));    relay_conn far_3_3901_1_b(.in(far_3_3901_0[1]), .out(far_3_3901_1[1]));
    assign layer_3[841] = far_3_3901_1[1] & ~far_3_3901_1[0]; 
    wire [1:0] far_3_3902_0;    relay_conn far_3_3902_0_a(.in(layer_2[178]), .out(far_3_3902_0[0]));    relay_conn far_3_3902_0_b(.in(layer_2[284]), .out(far_3_3902_0[1]));
    wire [1:0] far_3_3902_1;    relay_conn far_3_3902_1_a(.in(far_3_3902_0[0]), .out(far_3_3902_1[0]));    relay_conn far_3_3902_1_b(.in(far_3_3902_0[1]), .out(far_3_3902_1[1]));
    wire [1:0] far_3_3902_2;    relay_conn far_3_3902_2_a(.in(far_3_3902_1[0]), .out(far_3_3902_2[0]));    relay_conn far_3_3902_2_b(.in(far_3_3902_1[1]), .out(far_3_3902_2[1]));
    assign layer_3[842] = far_3_3902_2[1]; 
    assign layer_3[843] = ~layer_2[41]; 
    wire [1:0] far_3_3904_0;    relay_conn far_3_3904_0_a(.in(layer_2[777]), .out(far_3_3904_0[0]));    relay_conn far_3_3904_0_b(.in(layer_2[689]), .out(far_3_3904_0[1]));
    wire [1:0] far_3_3904_1;    relay_conn far_3_3904_1_a(.in(far_3_3904_0[0]), .out(far_3_3904_1[0]));    relay_conn far_3_3904_1_b(.in(far_3_3904_0[1]), .out(far_3_3904_1[1]));
    assign layer_3[844] = ~far_3_3904_1[0]; 
    wire [1:0] far_3_3905_0;    relay_conn far_3_3905_0_a(.in(layer_2[262]), .out(far_3_3905_0[0]));    relay_conn far_3_3905_0_b(.in(layer_2[137]), .out(far_3_3905_0[1]));
    wire [1:0] far_3_3905_1;    relay_conn far_3_3905_1_a(.in(far_3_3905_0[0]), .out(far_3_3905_1[0]));    relay_conn far_3_3905_1_b(.in(far_3_3905_0[1]), .out(far_3_3905_1[1]));
    wire [1:0] far_3_3905_2;    relay_conn far_3_3905_2_a(.in(far_3_3905_1[0]), .out(far_3_3905_2[0]));    relay_conn far_3_3905_2_b(.in(far_3_3905_1[1]), .out(far_3_3905_2[1]));
    assign layer_3[845] = ~(far_3_3905_2[0] & far_3_3905_2[1]); 
    assign layer_3[846] = ~layer_2[286] | (layer_2[286] & layer_2[287]); 
    assign layer_3[847] = layer_2[416] | layer_2[405]; 
    assign layer_3[848] = ~layer_2[703] | (layer_2[678] & layer_2[703]); 
    wire [1:0] far_3_3909_0;    relay_conn far_3_3909_0_a(.in(layer_2[298]), .out(far_3_3909_0[0]));    relay_conn far_3_3909_0_b(.in(layer_2[195]), .out(far_3_3909_0[1]));
    wire [1:0] far_3_3909_1;    relay_conn far_3_3909_1_a(.in(far_3_3909_0[0]), .out(far_3_3909_1[0]));    relay_conn far_3_3909_1_b(.in(far_3_3909_0[1]), .out(far_3_3909_1[1]));
    wire [1:0] far_3_3909_2;    relay_conn far_3_3909_2_a(.in(far_3_3909_1[0]), .out(far_3_3909_2[0]));    relay_conn far_3_3909_2_b(.in(far_3_3909_1[1]), .out(far_3_3909_2[1]));
    assign layer_3[849] = ~far_3_3909_2[0]; 
    assign layer_3[850] = ~(layer_2[1005] & layer_2[997]); 
    wire [1:0] far_3_3911_0;    relay_conn far_3_3911_0_a(.in(layer_2[206]), .out(far_3_3911_0[0]));    relay_conn far_3_3911_0_b(.in(layer_2[127]), .out(far_3_3911_0[1]));
    wire [1:0] far_3_3911_1;    relay_conn far_3_3911_1_a(.in(far_3_3911_0[0]), .out(far_3_3911_1[0]));    relay_conn far_3_3911_1_b(.in(far_3_3911_0[1]), .out(far_3_3911_1[1]));
    assign layer_3[851] = far_3_3911_1[1] & ~far_3_3911_1[0]; 
    wire [1:0] far_3_3912_0;    relay_conn far_3_3912_0_a(.in(layer_2[924]), .out(far_3_3912_0[0]));    relay_conn far_3_3912_0_b(.in(layer_2[975]), .out(far_3_3912_0[1]));
    assign layer_3[852] = far_3_3912_0[0] | far_3_3912_0[1]; 
    wire [1:0] far_3_3913_0;    relay_conn far_3_3913_0_a(.in(layer_2[771]), .out(far_3_3913_0[0]));    relay_conn far_3_3913_0_b(.in(layer_2[899]), .out(far_3_3913_0[1]));
    wire [1:0] far_3_3913_1;    relay_conn far_3_3913_1_a(.in(far_3_3913_0[0]), .out(far_3_3913_1[0]));    relay_conn far_3_3913_1_b(.in(far_3_3913_0[1]), .out(far_3_3913_1[1]));
    wire [1:0] far_3_3913_2;    relay_conn far_3_3913_2_a(.in(far_3_3913_1[0]), .out(far_3_3913_2[0]));    relay_conn far_3_3913_2_b(.in(far_3_3913_1[1]), .out(far_3_3913_2[1]));
    wire [1:0] far_3_3913_3;    relay_conn far_3_3913_3_a(.in(far_3_3913_2[0]), .out(far_3_3913_3[0]));    relay_conn far_3_3913_3_b(.in(far_3_3913_2[1]), .out(far_3_3913_3[1]));
    assign layer_3[853] = far_3_3913_3[1] & ~far_3_3913_3[0]; 
    assign layer_3[854] = layer_2[797]; 
    assign layer_3[855] = ~layer_2[588] | (layer_2[588] & layer_2[572]); 
    wire [1:0] far_3_3916_0;    relay_conn far_3_3916_0_a(.in(layer_2[827]), .out(far_3_3916_0[0]));    relay_conn far_3_3916_0_b(.in(layer_2[901]), .out(far_3_3916_0[1]));
    wire [1:0] far_3_3916_1;    relay_conn far_3_3916_1_a(.in(far_3_3916_0[0]), .out(far_3_3916_1[0]));    relay_conn far_3_3916_1_b(.in(far_3_3916_0[1]), .out(far_3_3916_1[1]));
    assign layer_3[856] = ~(far_3_3916_1[0] & far_3_3916_1[1]); 
    wire [1:0] far_3_3917_0;    relay_conn far_3_3917_0_a(.in(layer_2[783]), .out(far_3_3917_0[0]));    relay_conn far_3_3917_0_b(.in(layer_2[683]), .out(far_3_3917_0[1]));
    wire [1:0] far_3_3917_1;    relay_conn far_3_3917_1_a(.in(far_3_3917_0[0]), .out(far_3_3917_1[0]));    relay_conn far_3_3917_1_b(.in(far_3_3917_0[1]), .out(far_3_3917_1[1]));
    wire [1:0] far_3_3917_2;    relay_conn far_3_3917_2_a(.in(far_3_3917_1[0]), .out(far_3_3917_2[0]));    relay_conn far_3_3917_2_b(.in(far_3_3917_1[1]), .out(far_3_3917_2[1]));
    assign layer_3[857] = ~far_3_3917_2[0] | (far_3_3917_2[0] & far_3_3917_2[1]); 
    wire [1:0] far_3_3918_0;    relay_conn far_3_3918_0_a(.in(layer_2[79]), .out(far_3_3918_0[0]));    relay_conn far_3_3918_0_b(.in(layer_2[126]), .out(far_3_3918_0[1]));
    assign layer_3[858] = ~(far_3_3918_0[0] ^ far_3_3918_0[1]); 
    wire [1:0] far_3_3919_0;    relay_conn far_3_3919_0_a(.in(layer_2[325]), .out(far_3_3919_0[0]));    relay_conn far_3_3919_0_b(.in(layer_2[378]), .out(far_3_3919_0[1]));
    assign layer_3[859] = ~(far_3_3919_0[0] ^ far_3_3919_0[1]); 
    wire [1:0] far_3_3920_0;    relay_conn far_3_3920_0_a(.in(layer_2[768]), .out(far_3_3920_0[0]));    relay_conn far_3_3920_0_b(.in(layer_2[848]), .out(far_3_3920_0[1]));
    wire [1:0] far_3_3920_1;    relay_conn far_3_3920_1_a(.in(far_3_3920_0[0]), .out(far_3_3920_1[0]));    relay_conn far_3_3920_1_b(.in(far_3_3920_0[1]), .out(far_3_3920_1[1]));
    assign layer_3[860] = ~(far_3_3920_1[0] | far_3_3920_1[1]); 
    wire [1:0] far_3_3921_0;    relay_conn far_3_3921_0_a(.in(layer_2[553]), .out(far_3_3921_0[0]));    relay_conn far_3_3921_0_b(.in(layer_2[585]), .out(far_3_3921_0[1]));
    assign layer_3[861] = ~far_3_3921_0[1] | (far_3_3921_0[0] & far_3_3921_0[1]); 
    wire [1:0] far_3_3922_0;    relay_conn far_3_3922_0_a(.in(layer_2[244]), .out(far_3_3922_0[0]));    relay_conn far_3_3922_0_b(.in(layer_2[126]), .out(far_3_3922_0[1]));
    wire [1:0] far_3_3922_1;    relay_conn far_3_3922_1_a(.in(far_3_3922_0[0]), .out(far_3_3922_1[0]));    relay_conn far_3_3922_1_b(.in(far_3_3922_0[1]), .out(far_3_3922_1[1]));
    wire [1:0] far_3_3922_2;    relay_conn far_3_3922_2_a(.in(far_3_3922_1[0]), .out(far_3_3922_2[0]));    relay_conn far_3_3922_2_b(.in(far_3_3922_1[1]), .out(far_3_3922_2[1]));
    assign layer_3[862] = far_3_3922_2[1]; 
    assign layer_3[863] = layer_2[597]; 
    wire [1:0] far_3_3924_0;    relay_conn far_3_3924_0_a(.in(layer_2[327]), .out(far_3_3924_0[0]));    relay_conn far_3_3924_0_b(.in(layer_2[235]), .out(far_3_3924_0[1]));
    wire [1:0] far_3_3924_1;    relay_conn far_3_3924_1_a(.in(far_3_3924_0[0]), .out(far_3_3924_1[0]));    relay_conn far_3_3924_1_b(.in(far_3_3924_0[1]), .out(far_3_3924_1[1]));
    assign layer_3[864] = ~far_3_3924_1[1]; 
    wire [1:0] far_3_3925_0;    relay_conn far_3_3925_0_a(.in(layer_2[1001]), .out(far_3_3925_0[0]));    relay_conn far_3_3925_0_b(.in(layer_2[928]), .out(far_3_3925_0[1]));
    wire [1:0] far_3_3925_1;    relay_conn far_3_3925_1_a(.in(far_3_3925_0[0]), .out(far_3_3925_1[0]));    relay_conn far_3_3925_1_b(.in(far_3_3925_0[1]), .out(far_3_3925_1[1]));
    assign layer_3[865] = far_3_3925_1[1] & ~far_3_3925_1[0]; 
    wire [1:0] far_3_3926_0;    relay_conn far_3_3926_0_a(.in(layer_2[675]), .out(far_3_3926_0[0]));    relay_conn far_3_3926_0_b(.in(layer_2[725]), .out(far_3_3926_0[1]));
    assign layer_3[866] = far_3_3926_0[0]; 
    assign layer_3[867] = layer_2[467] ^ layer_2[477]; 
    wire [1:0] far_3_3928_0;    relay_conn far_3_3928_0_a(.in(layer_2[209]), .out(far_3_3928_0[0]));    relay_conn far_3_3928_0_b(.in(layer_2[335]), .out(far_3_3928_0[1]));
    wire [1:0] far_3_3928_1;    relay_conn far_3_3928_1_a(.in(far_3_3928_0[0]), .out(far_3_3928_1[0]));    relay_conn far_3_3928_1_b(.in(far_3_3928_0[1]), .out(far_3_3928_1[1]));
    wire [1:0] far_3_3928_2;    relay_conn far_3_3928_2_a(.in(far_3_3928_1[0]), .out(far_3_3928_2[0]));    relay_conn far_3_3928_2_b(.in(far_3_3928_1[1]), .out(far_3_3928_2[1]));
    assign layer_3[868] = far_3_3928_2[1] & ~far_3_3928_2[0]; 
    wire [1:0] far_3_3929_0;    relay_conn far_3_3929_0_a(.in(layer_2[248]), .out(far_3_3929_0[0]));    relay_conn far_3_3929_0_b(.in(layer_2[126]), .out(far_3_3929_0[1]));
    wire [1:0] far_3_3929_1;    relay_conn far_3_3929_1_a(.in(far_3_3929_0[0]), .out(far_3_3929_1[0]));    relay_conn far_3_3929_1_b(.in(far_3_3929_0[1]), .out(far_3_3929_1[1]));
    wire [1:0] far_3_3929_2;    relay_conn far_3_3929_2_a(.in(far_3_3929_1[0]), .out(far_3_3929_2[0]));    relay_conn far_3_3929_2_b(.in(far_3_3929_1[1]), .out(far_3_3929_2[1]));
    assign layer_3[869] = ~(far_3_3929_2[0] | far_3_3929_2[1]); 
    wire [1:0] far_3_3930_0;    relay_conn far_3_3930_0_a(.in(layer_2[746]), .out(far_3_3930_0[0]));    relay_conn far_3_3930_0_b(.in(layer_2[630]), .out(far_3_3930_0[1]));
    wire [1:0] far_3_3930_1;    relay_conn far_3_3930_1_a(.in(far_3_3930_0[0]), .out(far_3_3930_1[0]));    relay_conn far_3_3930_1_b(.in(far_3_3930_0[1]), .out(far_3_3930_1[1]));
    wire [1:0] far_3_3930_2;    relay_conn far_3_3930_2_a(.in(far_3_3930_1[0]), .out(far_3_3930_2[0]));    relay_conn far_3_3930_2_b(.in(far_3_3930_1[1]), .out(far_3_3930_2[1]));
    assign layer_3[870] = far_3_3930_2[0]; 
    wire [1:0] far_3_3931_0;    relay_conn far_3_3931_0_a(.in(layer_2[728]), .out(far_3_3931_0[0]));    relay_conn far_3_3931_0_b(.in(layer_2[666]), .out(far_3_3931_0[1]));
    assign layer_3[871] = far_3_3931_0[1]; 
    wire [1:0] far_3_3932_0;    relay_conn far_3_3932_0_a(.in(layer_2[234]), .out(far_3_3932_0[0]));    relay_conn far_3_3932_0_b(.in(layer_2[198]), .out(far_3_3932_0[1]));
    assign layer_3[872] = far_3_3932_0[1] & ~far_3_3932_0[0]; 
    assign layer_3[873] = layer_2[237] | layer_2[252]; 
    wire [1:0] far_3_3934_0;    relay_conn far_3_3934_0_a(.in(layer_2[985]), .out(far_3_3934_0[0]));    relay_conn far_3_3934_0_b(.in(layer_2[892]), .out(far_3_3934_0[1]));
    wire [1:0] far_3_3934_1;    relay_conn far_3_3934_1_a(.in(far_3_3934_0[0]), .out(far_3_3934_1[0]));    relay_conn far_3_3934_1_b(.in(far_3_3934_0[1]), .out(far_3_3934_1[1]));
    assign layer_3[874] = ~(far_3_3934_1[0] | far_3_3934_1[1]); 
    wire [1:0] far_3_3935_0;    relay_conn far_3_3935_0_a(.in(layer_2[119]), .out(far_3_3935_0[0]));    relay_conn far_3_3935_0_b(.in(layer_2[75]), .out(far_3_3935_0[1]));
    assign layer_3[875] = far_3_3935_0[0] & far_3_3935_0[1]; 
    wire [1:0] far_3_3936_0;    relay_conn far_3_3936_0_a(.in(layer_2[287]), .out(far_3_3936_0[0]));    relay_conn far_3_3936_0_b(.in(layer_2[412]), .out(far_3_3936_0[1]));
    wire [1:0] far_3_3936_1;    relay_conn far_3_3936_1_a(.in(far_3_3936_0[0]), .out(far_3_3936_1[0]));    relay_conn far_3_3936_1_b(.in(far_3_3936_0[1]), .out(far_3_3936_1[1]));
    wire [1:0] far_3_3936_2;    relay_conn far_3_3936_2_a(.in(far_3_3936_1[0]), .out(far_3_3936_2[0]));    relay_conn far_3_3936_2_b(.in(far_3_3936_1[1]), .out(far_3_3936_2[1]));
    assign layer_3[876] = far_3_3936_2[0]; 
    wire [1:0] far_3_3937_0;    relay_conn far_3_3937_0_a(.in(layer_2[262]), .out(far_3_3937_0[0]));    relay_conn far_3_3937_0_b(.in(layer_2[330]), .out(far_3_3937_0[1]));
    wire [1:0] far_3_3937_1;    relay_conn far_3_3937_1_a(.in(far_3_3937_0[0]), .out(far_3_3937_1[0]));    relay_conn far_3_3937_1_b(.in(far_3_3937_0[1]), .out(far_3_3937_1[1]));
    assign layer_3[877] = far_3_3937_1[0] ^ far_3_3937_1[1]; 
    assign layer_3[878] = ~(layer_2[101] & layer_2[102]); 
    wire [1:0] far_3_3939_0;    relay_conn far_3_3939_0_a(.in(layer_2[935]), .out(far_3_3939_0[0]));    relay_conn far_3_3939_0_b(.in(layer_2[880]), .out(far_3_3939_0[1]));
    assign layer_3[879] = ~far_3_3939_0[1] | (far_3_3939_0[0] & far_3_3939_0[1]); 
    wire [1:0] far_3_3940_0;    relay_conn far_3_3940_0_a(.in(layer_2[867]), .out(far_3_3940_0[0]));    relay_conn far_3_3940_0_b(.in(layer_2[785]), .out(far_3_3940_0[1]));
    wire [1:0] far_3_3940_1;    relay_conn far_3_3940_1_a(.in(far_3_3940_0[0]), .out(far_3_3940_1[0]));    relay_conn far_3_3940_1_b(.in(far_3_3940_0[1]), .out(far_3_3940_1[1]));
    assign layer_3[880] = ~far_3_3940_1[0]; 
    wire [1:0] far_3_3941_0;    relay_conn far_3_3941_0_a(.in(layer_2[177]), .out(far_3_3941_0[0]));    relay_conn far_3_3941_0_b(.in(layer_2[295]), .out(far_3_3941_0[1]));
    wire [1:0] far_3_3941_1;    relay_conn far_3_3941_1_a(.in(far_3_3941_0[0]), .out(far_3_3941_1[0]));    relay_conn far_3_3941_1_b(.in(far_3_3941_0[1]), .out(far_3_3941_1[1]));
    wire [1:0] far_3_3941_2;    relay_conn far_3_3941_2_a(.in(far_3_3941_1[0]), .out(far_3_3941_2[0]));    relay_conn far_3_3941_2_b(.in(far_3_3941_1[1]), .out(far_3_3941_2[1]));
    assign layer_3[881] = ~(far_3_3941_2[0] ^ far_3_3941_2[1]); 
    wire [1:0] far_3_3942_0;    relay_conn far_3_3942_0_a(.in(layer_2[447]), .out(far_3_3942_0[0]));    relay_conn far_3_3942_0_b(.in(layer_2[550]), .out(far_3_3942_0[1]));
    wire [1:0] far_3_3942_1;    relay_conn far_3_3942_1_a(.in(far_3_3942_0[0]), .out(far_3_3942_1[0]));    relay_conn far_3_3942_1_b(.in(far_3_3942_0[1]), .out(far_3_3942_1[1]));
    wire [1:0] far_3_3942_2;    relay_conn far_3_3942_2_a(.in(far_3_3942_1[0]), .out(far_3_3942_2[0]));    relay_conn far_3_3942_2_b(.in(far_3_3942_1[1]), .out(far_3_3942_2[1]));
    assign layer_3[882] = ~(far_3_3942_2[0] | far_3_3942_2[1]); 
    wire [1:0] far_3_3943_0;    relay_conn far_3_3943_0_a(.in(layer_2[198]), .out(far_3_3943_0[0]));    relay_conn far_3_3943_0_b(.in(layer_2[250]), .out(far_3_3943_0[1]));
    assign layer_3[883] = far_3_3943_0[0] & ~far_3_3943_0[1]; 
    wire [1:0] far_3_3944_0;    relay_conn far_3_3944_0_a(.in(layer_2[264]), .out(far_3_3944_0[0]));    relay_conn far_3_3944_0_b(.in(layer_2[314]), .out(far_3_3944_0[1]));
    assign layer_3[884] = ~far_3_3944_0[1] | (far_3_3944_0[0] & far_3_3944_0[1]); 
    wire [1:0] far_3_3945_0;    relay_conn far_3_3945_0_a(.in(layer_2[303]), .out(far_3_3945_0[0]));    relay_conn far_3_3945_0_b(.in(layer_2[177]), .out(far_3_3945_0[1]));
    wire [1:0] far_3_3945_1;    relay_conn far_3_3945_1_a(.in(far_3_3945_0[0]), .out(far_3_3945_1[0]));    relay_conn far_3_3945_1_b(.in(far_3_3945_0[1]), .out(far_3_3945_1[1]));
    wire [1:0] far_3_3945_2;    relay_conn far_3_3945_2_a(.in(far_3_3945_1[0]), .out(far_3_3945_2[0]));    relay_conn far_3_3945_2_b(.in(far_3_3945_1[1]), .out(far_3_3945_2[1]));
    assign layer_3[885] = far_3_3945_2[0] | far_3_3945_2[1]; 
    assign layer_3[886] = ~layer_2[498] | (layer_2[505] & layer_2[498]); 
    wire [1:0] far_3_3947_0;    relay_conn far_3_3947_0_a(.in(layer_2[835]), .out(far_3_3947_0[0]));    relay_conn far_3_3947_0_b(.in(layer_2[787]), .out(far_3_3947_0[1]));
    assign layer_3[887] = far_3_3947_0[0] | far_3_3947_0[1]; 
    wire [1:0] far_3_3948_0;    relay_conn far_3_3948_0_a(.in(layer_2[428]), .out(far_3_3948_0[0]));    relay_conn far_3_3948_0_b(.in(layer_2[505]), .out(far_3_3948_0[1]));
    wire [1:0] far_3_3948_1;    relay_conn far_3_3948_1_a(.in(far_3_3948_0[0]), .out(far_3_3948_1[0]));    relay_conn far_3_3948_1_b(.in(far_3_3948_0[1]), .out(far_3_3948_1[1]));
    assign layer_3[888] = far_3_3948_1[0] & far_3_3948_1[1]; 
    wire [1:0] far_3_3949_0;    relay_conn far_3_3949_0_a(.in(layer_2[336]), .out(far_3_3949_0[0]));    relay_conn far_3_3949_0_b(.in(layer_2[260]), .out(far_3_3949_0[1]));
    wire [1:0] far_3_3949_1;    relay_conn far_3_3949_1_a(.in(far_3_3949_0[0]), .out(far_3_3949_1[0]));    relay_conn far_3_3949_1_b(.in(far_3_3949_0[1]), .out(far_3_3949_1[1]));
    assign layer_3[889] = ~far_3_3949_1[1] | (far_3_3949_1[0] & far_3_3949_1[1]); 
    wire [1:0] far_3_3950_0;    relay_conn far_3_3950_0_a(.in(layer_2[354]), .out(far_3_3950_0[0]));    relay_conn far_3_3950_0_b(.in(layer_2[420]), .out(far_3_3950_0[1]));
    wire [1:0] far_3_3950_1;    relay_conn far_3_3950_1_a(.in(far_3_3950_0[0]), .out(far_3_3950_1[0]));    relay_conn far_3_3950_1_b(.in(far_3_3950_0[1]), .out(far_3_3950_1[1]));
    assign layer_3[890] = far_3_3950_1[0] | far_3_3950_1[1]; 
    wire [1:0] far_3_3951_0;    relay_conn far_3_3951_0_a(.in(layer_2[1011]), .out(far_3_3951_0[0]));    relay_conn far_3_3951_0_b(.in(layer_2[965]), .out(far_3_3951_0[1]));
    assign layer_3[891] = far_3_3951_0[0] | far_3_3951_0[1]; 
    wire [1:0] far_3_3952_0;    relay_conn far_3_3952_0_a(.in(layer_2[911]), .out(far_3_3952_0[0]));    relay_conn far_3_3952_0_b(.in(layer_2[835]), .out(far_3_3952_0[1]));
    wire [1:0] far_3_3952_1;    relay_conn far_3_3952_1_a(.in(far_3_3952_0[0]), .out(far_3_3952_1[0]));    relay_conn far_3_3952_1_b(.in(far_3_3952_0[1]), .out(far_3_3952_1[1]));
    assign layer_3[892] = far_3_3952_1[0]; 
    wire [1:0] far_3_3953_0;    relay_conn far_3_3953_0_a(.in(layer_2[444]), .out(far_3_3953_0[0]));    relay_conn far_3_3953_0_b(.in(layer_2[342]), .out(far_3_3953_0[1]));
    wire [1:0] far_3_3953_1;    relay_conn far_3_3953_1_a(.in(far_3_3953_0[0]), .out(far_3_3953_1[0]));    relay_conn far_3_3953_1_b(.in(far_3_3953_0[1]), .out(far_3_3953_1[1]));
    wire [1:0] far_3_3953_2;    relay_conn far_3_3953_2_a(.in(far_3_3953_1[0]), .out(far_3_3953_2[0]));    relay_conn far_3_3953_2_b(.in(far_3_3953_1[1]), .out(far_3_3953_2[1]));
    assign layer_3[893] = far_3_3953_2[1] & ~far_3_3953_2[0]; 
    assign layer_3[894] = ~layer_2[319] | (layer_2[319] & layer_2[327]); 
    wire [1:0] far_3_3955_0;    relay_conn far_3_3955_0_a(.in(layer_2[806]), .out(far_3_3955_0[0]));    relay_conn far_3_3955_0_b(.in(layer_2[913]), .out(far_3_3955_0[1]));
    wire [1:0] far_3_3955_1;    relay_conn far_3_3955_1_a(.in(far_3_3955_0[0]), .out(far_3_3955_1[0]));    relay_conn far_3_3955_1_b(.in(far_3_3955_0[1]), .out(far_3_3955_1[1]));
    wire [1:0] far_3_3955_2;    relay_conn far_3_3955_2_a(.in(far_3_3955_1[0]), .out(far_3_3955_2[0]));    relay_conn far_3_3955_2_b(.in(far_3_3955_1[1]), .out(far_3_3955_2[1]));
    assign layer_3[895] = ~(far_3_3955_2[0] | far_3_3955_2[1]); 
    wire [1:0] far_3_3956_0;    relay_conn far_3_3956_0_a(.in(layer_2[960]), .out(far_3_3956_0[0]));    relay_conn far_3_3956_0_b(.in(layer_2[842]), .out(far_3_3956_0[1]));
    wire [1:0] far_3_3956_1;    relay_conn far_3_3956_1_a(.in(far_3_3956_0[0]), .out(far_3_3956_1[0]));    relay_conn far_3_3956_1_b(.in(far_3_3956_0[1]), .out(far_3_3956_1[1]));
    wire [1:0] far_3_3956_2;    relay_conn far_3_3956_2_a(.in(far_3_3956_1[0]), .out(far_3_3956_2[0]));    relay_conn far_3_3956_2_b(.in(far_3_3956_1[1]), .out(far_3_3956_2[1]));
    assign layer_3[896] = ~(far_3_3956_2[0] ^ far_3_3956_2[1]); 
    assign layer_3[897] = layer_2[748] & ~layer_2[727]; 
    wire [1:0] far_3_3958_0;    relay_conn far_3_3958_0_a(.in(layer_2[433]), .out(far_3_3958_0[0]));    relay_conn far_3_3958_0_b(.in(layer_2[324]), .out(far_3_3958_0[1]));
    wire [1:0] far_3_3958_1;    relay_conn far_3_3958_1_a(.in(far_3_3958_0[0]), .out(far_3_3958_1[0]));    relay_conn far_3_3958_1_b(.in(far_3_3958_0[1]), .out(far_3_3958_1[1]));
    wire [1:0] far_3_3958_2;    relay_conn far_3_3958_2_a(.in(far_3_3958_1[0]), .out(far_3_3958_2[0]));    relay_conn far_3_3958_2_b(.in(far_3_3958_1[1]), .out(far_3_3958_2[1]));
    assign layer_3[898] = far_3_3958_2[1] & ~far_3_3958_2[0]; 
    wire [1:0] far_3_3959_0;    relay_conn far_3_3959_0_a(.in(layer_2[543]), .out(far_3_3959_0[0]));    relay_conn far_3_3959_0_b(.in(layer_2[626]), .out(far_3_3959_0[1]));
    wire [1:0] far_3_3959_1;    relay_conn far_3_3959_1_a(.in(far_3_3959_0[0]), .out(far_3_3959_1[0]));    relay_conn far_3_3959_1_b(.in(far_3_3959_0[1]), .out(far_3_3959_1[1]));
    assign layer_3[899] = far_3_3959_1[0]; 
    assign layer_3[900] = ~layer_2[412] | (layer_2[412] & layer_2[389]); 
    wire [1:0] far_3_3961_0;    relay_conn far_3_3961_0_a(.in(layer_2[733]), .out(far_3_3961_0[0]));    relay_conn far_3_3961_0_b(.in(layer_2[774]), .out(far_3_3961_0[1]));
    assign layer_3[901] = far_3_3961_0[0]; 
    wire [1:0] far_3_3962_0;    relay_conn far_3_3962_0_a(.in(layer_2[94]), .out(far_3_3962_0[0]));    relay_conn far_3_3962_0_b(.in(layer_2[208]), .out(far_3_3962_0[1]));
    wire [1:0] far_3_3962_1;    relay_conn far_3_3962_1_a(.in(far_3_3962_0[0]), .out(far_3_3962_1[0]));    relay_conn far_3_3962_1_b(.in(far_3_3962_0[1]), .out(far_3_3962_1[1]));
    wire [1:0] far_3_3962_2;    relay_conn far_3_3962_2_a(.in(far_3_3962_1[0]), .out(far_3_3962_2[0]));    relay_conn far_3_3962_2_b(.in(far_3_3962_1[1]), .out(far_3_3962_2[1]));
    assign layer_3[902] = ~(far_3_3962_2[0] ^ far_3_3962_2[1]); 
    assign layer_3[903] = layer_2[511] & layer_2[480]; 
    wire [1:0] far_3_3964_0;    relay_conn far_3_3964_0_a(.in(layer_2[410]), .out(far_3_3964_0[0]));    relay_conn far_3_3964_0_b(.in(layer_2[502]), .out(far_3_3964_0[1]));
    wire [1:0] far_3_3964_1;    relay_conn far_3_3964_1_a(.in(far_3_3964_0[0]), .out(far_3_3964_1[0]));    relay_conn far_3_3964_1_b(.in(far_3_3964_0[1]), .out(far_3_3964_1[1]));
    assign layer_3[904] = ~(far_3_3964_1[0] | far_3_3964_1[1]); 
    assign layer_3[905] = ~layer_2[352] | (layer_2[332] & layer_2[352]); 
    wire [1:0] far_3_3966_0;    relay_conn far_3_3966_0_a(.in(layer_2[522]), .out(far_3_3966_0[0]));    relay_conn far_3_3966_0_b(.in(layer_2[488]), .out(far_3_3966_0[1]));
    assign layer_3[906] = far_3_3966_0[0] & far_3_3966_0[1]; 
    assign layer_3[907] = layer_2[260] | layer_2[252]; 
    assign layer_3[908] = layer_2[733] & ~layer_2[726]; 
    wire [1:0] far_3_3969_0;    relay_conn far_3_3969_0_a(.in(layer_2[839]), .out(far_3_3969_0[0]));    relay_conn far_3_3969_0_b(.in(layer_2[794]), .out(far_3_3969_0[1]));
    assign layer_3[909] = far_3_3969_0[1] & ~far_3_3969_0[0]; 
    assign layer_3[910] = ~layer_2[645] | (layer_2[623] & layer_2[645]); 
    wire [1:0] far_3_3971_0;    relay_conn far_3_3971_0_a(.in(layer_2[144]), .out(far_3_3971_0[0]));    relay_conn far_3_3971_0_b(.in(layer_2[57]), .out(far_3_3971_0[1]));
    wire [1:0] far_3_3971_1;    relay_conn far_3_3971_1_a(.in(far_3_3971_0[0]), .out(far_3_3971_1[0]));    relay_conn far_3_3971_1_b(.in(far_3_3971_0[1]), .out(far_3_3971_1[1]));
    assign layer_3[911] = ~(far_3_3971_1[0] | far_3_3971_1[1]); 
    wire [1:0] far_3_3972_0;    relay_conn far_3_3972_0_a(.in(layer_2[662]), .out(far_3_3972_0[0]));    relay_conn far_3_3972_0_b(.in(layer_2[775]), .out(far_3_3972_0[1]));
    wire [1:0] far_3_3972_1;    relay_conn far_3_3972_1_a(.in(far_3_3972_0[0]), .out(far_3_3972_1[0]));    relay_conn far_3_3972_1_b(.in(far_3_3972_0[1]), .out(far_3_3972_1[1]));
    wire [1:0] far_3_3972_2;    relay_conn far_3_3972_2_a(.in(far_3_3972_1[0]), .out(far_3_3972_2[0]));    relay_conn far_3_3972_2_b(.in(far_3_3972_1[1]), .out(far_3_3972_2[1]));
    assign layer_3[912] = ~(far_3_3972_2[0] ^ far_3_3972_2[1]); 
    wire [1:0] far_3_3973_0;    relay_conn far_3_3973_0_a(.in(layer_2[289]), .out(far_3_3973_0[0]));    relay_conn far_3_3973_0_b(.in(layer_2[208]), .out(far_3_3973_0[1]));
    wire [1:0] far_3_3973_1;    relay_conn far_3_3973_1_a(.in(far_3_3973_0[0]), .out(far_3_3973_1[0]));    relay_conn far_3_3973_1_b(.in(far_3_3973_0[1]), .out(far_3_3973_1[1]));
    assign layer_3[913] = ~(far_3_3973_1[0] | far_3_3973_1[1]); 
    assign layer_3[914] = layer_2[700]; 
    wire [1:0] far_3_3975_0;    relay_conn far_3_3975_0_a(.in(layer_2[512]), .out(far_3_3975_0[0]));    relay_conn far_3_3975_0_b(.in(layer_2[466]), .out(far_3_3975_0[1]));
    assign layer_3[915] = ~far_3_3975_0[0]; 
    assign layer_3[916] = ~layer_2[560]; 
    wire [1:0] far_3_3977_0;    relay_conn far_3_3977_0_a(.in(layer_2[839]), .out(far_3_3977_0[0]));    relay_conn far_3_3977_0_b(.in(layer_2[927]), .out(far_3_3977_0[1]));
    wire [1:0] far_3_3977_1;    relay_conn far_3_3977_1_a(.in(far_3_3977_0[0]), .out(far_3_3977_1[0]));    relay_conn far_3_3977_1_b(.in(far_3_3977_0[1]), .out(far_3_3977_1[1]));
    assign layer_3[917] = far_3_3977_1[0]; 
    assign layer_3[918] = ~(layer_2[944] | layer_2[927]); 
    assign layer_3[919] = layer_2[986] | layer_2[988]; 
    wire [1:0] far_3_3980_0;    relay_conn far_3_3980_0_a(.in(layer_2[628]), .out(far_3_3980_0[0]));    relay_conn far_3_3980_0_b(.in(layer_2[520]), .out(far_3_3980_0[1]));
    wire [1:0] far_3_3980_1;    relay_conn far_3_3980_1_a(.in(far_3_3980_0[0]), .out(far_3_3980_1[0]));    relay_conn far_3_3980_1_b(.in(far_3_3980_0[1]), .out(far_3_3980_1[1]));
    wire [1:0] far_3_3980_2;    relay_conn far_3_3980_2_a(.in(far_3_3980_1[0]), .out(far_3_3980_2[0]));    relay_conn far_3_3980_2_b(.in(far_3_3980_1[1]), .out(far_3_3980_2[1]));
    assign layer_3[920] = ~far_3_3980_2[1] | (far_3_3980_2[0] & far_3_3980_2[1]); 
    wire [1:0] far_3_3981_0;    relay_conn far_3_3981_0_a(.in(layer_2[57]), .out(far_3_3981_0[0]));    relay_conn far_3_3981_0_b(.in(layer_2[144]), .out(far_3_3981_0[1]));
    wire [1:0] far_3_3981_1;    relay_conn far_3_3981_1_a(.in(far_3_3981_0[0]), .out(far_3_3981_1[0]));    relay_conn far_3_3981_1_b(.in(far_3_3981_0[1]), .out(far_3_3981_1[1]));
    assign layer_3[921] = far_3_3981_1[1] & ~far_3_3981_1[0]; 
    assign layer_3[922] = layer_2[640] ^ layer_2[654]; 
    wire [1:0] far_3_3983_0;    relay_conn far_3_3983_0_a(.in(layer_2[182]), .out(far_3_3983_0[0]));    relay_conn far_3_3983_0_b(.in(layer_2[104]), .out(far_3_3983_0[1]));
    wire [1:0] far_3_3983_1;    relay_conn far_3_3983_1_a(.in(far_3_3983_0[0]), .out(far_3_3983_1[0]));    relay_conn far_3_3983_1_b(.in(far_3_3983_0[1]), .out(far_3_3983_1[1]));
    assign layer_3[923] = ~(far_3_3983_1[0] | far_3_3983_1[1]); 
    wire [1:0] far_3_3984_0;    relay_conn far_3_3984_0_a(.in(layer_2[360]), .out(far_3_3984_0[0]));    relay_conn far_3_3984_0_b(.in(layer_2[280]), .out(far_3_3984_0[1]));
    wire [1:0] far_3_3984_1;    relay_conn far_3_3984_1_a(.in(far_3_3984_0[0]), .out(far_3_3984_1[0]));    relay_conn far_3_3984_1_b(.in(far_3_3984_0[1]), .out(far_3_3984_1[1]));
    assign layer_3[924] = ~far_3_3984_1[1]; 
    wire [1:0] far_3_3985_0;    relay_conn far_3_3985_0_a(.in(layer_2[852]), .out(far_3_3985_0[0]));    relay_conn far_3_3985_0_b(.in(layer_2[813]), .out(far_3_3985_0[1]));
    assign layer_3[925] = far_3_3985_0[0] & far_3_3985_0[1]; 
    wire [1:0] far_3_3986_0;    relay_conn far_3_3986_0_a(.in(layer_2[949]), .out(far_3_3986_0[0]));    relay_conn far_3_3986_0_b(.in(layer_2[912]), .out(far_3_3986_0[1]));
    assign layer_3[926] = far_3_3986_0[0] & ~far_3_3986_0[1]; 
    assign layer_3[927] = ~layer_2[80] | (layer_2[80] & layer_2[49]); 
    wire [1:0] far_3_3988_0;    relay_conn far_3_3988_0_a(.in(layer_2[797]), .out(far_3_3988_0[0]));    relay_conn far_3_3988_0_b(.in(layer_2[913]), .out(far_3_3988_0[1]));
    wire [1:0] far_3_3988_1;    relay_conn far_3_3988_1_a(.in(far_3_3988_0[0]), .out(far_3_3988_1[0]));    relay_conn far_3_3988_1_b(.in(far_3_3988_0[1]), .out(far_3_3988_1[1]));
    wire [1:0] far_3_3988_2;    relay_conn far_3_3988_2_a(.in(far_3_3988_1[0]), .out(far_3_3988_2[0]));    relay_conn far_3_3988_2_b(.in(far_3_3988_1[1]), .out(far_3_3988_2[1]));
    assign layer_3[928] = ~far_3_3988_2[1] | (far_3_3988_2[0] & far_3_3988_2[1]); 
    assign layer_3[929] = ~layer_2[897] | (layer_2[897] & layer_2[872]); 
    assign layer_3[930] = ~(layer_2[471] | layer_2[489]); 
    wire [1:0] far_3_3991_0;    relay_conn far_3_3991_0_a(.in(layer_2[362]), .out(far_3_3991_0[0]));    relay_conn far_3_3991_0_b(.in(layer_2[421]), .out(far_3_3991_0[1]));
    assign layer_3[931] = ~far_3_3991_0[1]; 
    wire [1:0] far_3_3992_0;    relay_conn far_3_3992_0_a(.in(layer_2[539]), .out(far_3_3992_0[0]));    relay_conn far_3_3992_0_b(.in(layer_2[429]), .out(far_3_3992_0[1]));
    wire [1:0] far_3_3992_1;    relay_conn far_3_3992_1_a(.in(far_3_3992_0[0]), .out(far_3_3992_1[0]));    relay_conn far_3_3992_1_b(.in(far_3_3992_0[1]), .out(far_3_3992_1[1]));
    wire [1:0] far_3_3992_2;    relay_conn far_3_3992_2_a(.in(far_3_3992_1[0]), .out(far_3_3992_2[0]));    relay_conn far_3_3992_2_b(.in(far_3_3992_1[1]), .out(far_3_3992_2[1]));
    assign layer_3[932] = ~far_3_3992_2[0]; 
    wire [1:0] far_3_3993_0;    relay_conn far_3_3993_0_a(.in(layer_2[170]), .out(far_3_3993_0[0]));    relay_conn far_3_3993_0_b(.in(layer_2[247]), .out(far_3_3993_0[1]));
    wire [1:0] far_3_3993_1;    relay_conn far_3_3993_1_a(.in(far_3_3993_0[0]), .out(far_3_3993_1[0]));    relay_conn far_3_3993_1_b(.in(far_3_3993_0[1]), .out(far_3_3993_1[1]));
    assign layer_3[933] = far_3_3993_1[0] & ~far_3_3993_1[1]; 
    wire [1:0] far_3_3994_0;    relay_conn far_3_3994_0_a(.in(layer_2[273]), .out(far_3_3994_0[0]));    relay_conn far_3_3994_0_b(.in(layer_2[215]), .out(far_3_3994_0[1]));
    assign layer_3[934] = ~(far_3_3994_0[0] | far_3_3994_0[1]); 
    assign layer_3[935] = layer_2[826] & ~layer_2[827]; 
    wire [1:0] far_3_3996_0;    relay_conn far_3_3996_0_a(.in(layer_2[920]), .out(far_3_3996_0[0]));    relay_conn far_3_3996_0_b(.in(layer_2[813]), .out(far_3_3996_0[1]));
    wire [1:0] far_3_3996_1;    relay_conn far_3_3996_1_a(.in(far_3_3996_0[0]), .out(far_3_3996_1[0]));    relay_conn far_3_3996_1_b(.in(far_3_3996_0[1]), .out(far_3_3996_1[1]));
    wire [1:0] far_3_3996_2;    relay_conn far_3_3996_2_a(.in(far_3_3996_1[0]), .out(far_3_3996_2[0]));    relay_conn far_3_3996_2_b(.in(far_3_3996_1[1]), .out(far_3_3996_2[1]));
    assign layer_3[936] = far_3_3996_2[0] & far_3_3996_2[1]; 
    assign layer_3[937] = layer_2[58] & ~layer_2[62]; 
    wire [1:0] far_3_3998_0;    relay_conn far_3_3998_0_a(.in(layer_2[71]), .out(far_3_3998_0[0]));    relay_conn far_3_3998_0_b(.in(layer_2[154]), .out(far_3_3998_0[1]));
    wire [1:0] far_3_3998_1;    relay_conn far_3_3998_1_a(.in(far_3_3998_0[0]), .out(far_3_3998_1[0]));    relay_conn far_3_3998_1_b(.in(far_3_3998_0[1]), .out(far_3_3998_1[1]));
    assign layer_3[938] = ~(far_3_3998_1[0] | far_3_3998_1[1]); 
    wire [1:0] far_3_3999_0;    relay_conn far_3_3999_0_a(.in(layer_2[695]), .out(far_3_3999_0[0]));    relay_conn far_3_3999_0_b(.in(layer_2[591]), .out(far_3_3999_0[1]));
    wire [1:0] far_3_3999_1;    relay_conn far_3_3999_1_a(.in(far_3_3999_0[0]), .out(far_3_3999_1[0]));    relay_conn far_3_3999_1_b(.in(far_3_3999_0[1]), .out(far_3_3999_1[1]));
    wire [1:0] far_3_3999_2;    relay_conn far_3_3999_2_a(.in(far_3_3999_1[0]), .out(far_3_3999_2[0]));    relay_conn far_3_3999_2_b(.in(far_3_3999_1[1]), .out(far_3_3999_2[1]));
    assign layer_3[939] = ~far_3_3999_2[0] | (far_3_3999_2[0] & far_3_3999_2[1]); 
    wire [1:0] far_3_4000_0;    relay_conn far_3_4000_0_a(.in(layer_2[674]), .out(far_3_4000_0[0]));    relay_conn far_3_4000_0_b(.in(layer_2[749]), .out(far_3_4000_0[1]));
    wire [1:0] far_3_4000_1;    relay_conn far_3_4000_1_a(.in(far_3_4000_0[0]), .out(far_3_4000_1[0]));    relay_conn far_3_4000_1_b(.in(far_3_4000_0[1]), .out(far_3_4000_1[1]));
    assign layer_3[940] = ~far_3_4000_1[1] | (far_3_4000_1[0] & far_3_4000_1[1]); 
    wire [1:0] far_3_4001_0;    relay_conn far_3_4001_0_a(.in(layer_2[120]), .out(far_3_4001_0[0]));    relay_conn far_3_4001_0_b(.in(layer_2[218]), .out(far_3_4001_0[1]));
    wire [1:0] far_3_4001_1;    relay_conn far_3_4001_1_a(.in(far_3_4001_0[0]), .out(far_3_4001_1[0]));    relay_conn far_3_4001_1_b(.in(far_3_4001_0[1]), .out(far_3_4001_1[1]));
    wire [1:0] far_3_4001_2;    relay_conn far_3_4001_2_a(.in(far_3_4001_1[0]), .out(far_3_4001_2[0]));    relay_conn far_3_4001_2_b(.in(far_3_4001_1[1]), .out(far_3_4001_2[1]));
    assign layer_3[941] = far_3_4001_2[0] & far_3_4001_2[1]; 
    wire [1:0] far_3_4002_0;    relay_conn far_3_4002_0_a(.in(layer_2[115]), .out(far_3_4002_0[0]));    relay_conn far_3_4002_0_b(.in(layer_2[64]), .out(far_3_4002_0[1]));
    assign layer_3[942] = far_3_4002_0[0] & far_3_4002_0[1]; 
    assign layer_3[943] = ~layer_2[483] | (layer_2[483] & layer_2[489]); 
    wire [1:0] far_3_4004_0;    relay_conn far_3_4004_0_a(.in(layer_2[155]), .out(far_3_4004_0[0]));    relay_conn far_3_4004_0_b(.in(layer_2[54]), .out(far_3_4004_0[1]));
    wire [1:0] far_3_4004_1;    relay_conn far_3_4004_1_a(.in(far_3_4004_0[0]), .out(far_3_4004_1[0]));    relay_conn far_3_4004_1_b(.in(far_3_4004_0[1]), .out(far_3_4004_1[1]));
    wire [1:0] far_3_4004_2;    relay_conn far_3_4004_2_a(.in(far_3_4004_1[0]), .out(far_3_4004_2[0]));    relay_conn far_3_4004_2_b(.in(far_3_4004_1[1]), .out(far_3_4004_2[1]));
    assign layer_3[944] = ~(far_3_4004_2[0] ^ far_3_4004_2[1]); 
    wire [1:0] far_3_4005_0;    relay_conn far_3_4005_0_a(.in(layer_2[863]), .out(far_3_4005_0[0]));    relay_conn far_3_4005_0_b(.in(layer_2[826]), .out(far_3_4005_0[1]));
    assign layer_3[945] = ~(far_3_4005_0[0] | far_3_4005_0[1]); 
    wire [1:0] far_3_4006_0;    relay_conn far_3_4006_0_a(.in(layer_2[160]), .out(far_3_4006_0[0]));    relay_conn far_3_4006_0_b(.in(layer_2[278]), .out(far_3_4006_0[1]));
    wire [1:0] far_3_4006_1;    relay_conn far_3_4006_1_a(.in(far_3_4006_0[0]), .out(far_3_4006_1[0]));    relay_conn far_3_4006_1_b(.in(far_3_4006_0[1]), .out(far_3_4006_1[1]));
    wire [1:0] far_3_4006_2;    relay_conn far_3_4006_2_a(.in(far_3_4006_1[0]), .out(far_3_4006_2[0]));    relay_conn far_3_4006_2_b(.in(far_3_4006_1[1]), .out(far_3_4006_2[1]));
    assign layer_3[946] = far_3_4006_2[0] ^ far_3_4006_2[1]; 
    wire [1:0] far_3_4007_0;    relay_conn far_3_4007_0_a(.in(layer_2[361]), .out(far_3_4007_0[0]));    relay_conn far_3_4007_0_b(.in(layer_2[404]), .out(far_3_4007_0[1]));
    assign layer_3[947] = far_3_4007_0[1] & ~far_3_4007_0[0]; 
    wire [1:0] far_3_4008_0;    relay_conn far_3_4008_0_a(.in(layer_2[487]), .out(far_3_4008_0[0]));    relay_conn far_3_4008_0_b(.in(layer_2[564]), .out(far_3_4008_0[1]));
    wire [1:0] far_3_4008_1;    relay_conn far_3_4008_1_a(.in(far_3_4008_0[0]), .out(far_3_4008_1[0]));    relay_conn far_3_4008_1_b(.in(far_3_4008_0[1]), .out(far_3_4008_1[1]));
    assign layer_3[948] = far_3_4008_1[0] & far_3_4008_1[1]; 
    wire [1:0] far_3_4009_0;    relay_conn far_3_4009_0_a(.in(layer_2[640]), .out(far_3_4009_0[0]));    relay_conn far_3_4009_0_b(.in(layer_2[674]), .out(far_3_4009_0[1]));
    assign layer_3[949] = ~far_3_4009_0[1] | (far_3_4009_0[0] & far_3_4009_0[1]); 
    wire [1:0] far_3_4010_0;    relay_conn far_3_4010_0_a(.in(layer_2[966]), .out(far_3_4010_0[0]));    relay_conn far_3_4010_0_b(.in(layer_2[1005]), .out(far_3_4010_0[1]));
    assign layer_3[950] = ~far_3_4010_0[1]; 
    wire [1:0] far_3_4011_0;    relay_conn far_3_4011_0_a(.in(layer_2[628]), .out(far_3_4011_0[0]));    relay_conn far_3_4011_0_b(.in(layer_2[747]), .out(far_3_4011_0[1]));
    wire [1:0] far_3_4011_1;    relay_conn far_3_4011_1_a(.in(far_3_4011_0[0]), .out(far_3_4011_1[0]));    relay_conn far_3_4011_1_b(.in(far_3_4011_0[1]), .out(far_3_4011_1[1]));
    wire [1:0] far_3_4011_2;    relay_conn far_3_4011_2_a(.in(far_3_4011_1[0]), .out(far_3_4011_2[0]));    relay_conn far_3_4011_2_b(.in(far_3_4011_1[1]), .out(far_3_4011_2[1]));
    assign layer_3[951] = ~(far_3_4011_2[0] & far_3_4011_2[1]); 
    wire [1:0] far_3_4012_0;    relay_conn far_3_4012_0_a(.in(layer_2[131]), .out(far_3_4012_0[0]));    relay_conn far_3_4012_0_b(.in(layer_2[223]), .out(far_3_4012_0[1]));
    wire [1:0] far_3_4012_1;    relay_conn far_3_4012_1_a(.in(far_3_4012_0[0]), .out(far_3_4012_1[0]));    relay_conn far_3_4012_1_b(.in(far_3_4012_0[1]), .out(far_3_4012_1[1]));
    assign layer_3[952] = ~(far_3_4012_1[0] | far_3_4012_1[1]); 
    wire [1:0] far_3_4013_0;    relay_conn far_3_4013_0_a(.in(layer_2[235]), .out(far_3_4013_0[0]));    relay_conn far_3_4013_0_b(.in(layer_2[309]), .out(far_3_4013_0[1]));
    wire [1:0] far_3_4013_1;    relay_conn far_3_4013_1_a(.in(far_3_4013_0[0]), .out(far_3_4013_1[0]));    relay_conn far_3_4013_1_b(.in(far_3_4013_0[1]), .out(far_3_4013_1[1]));
    assign layer_3[953] = ~far_3_4013_1[1] | (far_3_4013_1[0] & far_3_4013_1[1]); 
    wire [1:0] far_3_4014_0;    relay_conn far_3_4014_0_a(.in(layer_2[63]), .out(far_3_4014_0[0]));    relay_conn far_3_4014_0_b(.in(layer_2[8]), .out(far_3_4014_0[1]));
    assign layer_3[954] = far_3_4014_0[1]; 
    wire [1:0] far_3_4015_0;    relay_conn far_3_4015_0_a(.in(layer_2[489]), .out(far_3_4015_0[0]));    relay_conn far_3_4015_0_b(.in(layer_2[371]), .out(far_3_4015_0[1]));
    wire [1:0] far_3_4015_1;    relay_conn far_3_4015_1_a(.in(far_3_4015_0[0]), .out(far_3_4015_1[0]));    relay_conn far_3_4015_1_b(.in(far_3_4015_0[1]), .out(far_3_4015_1[1]));
    wire [1:0] far_3_4015_2;    relay_conn far_3_4015_2_a(.in(far_3_4015_1[0]), .out(far_3_4015_2[0]));    relay_conn far_3_4015_2_b(.in(far_3_4015_1[1]), .out(far_3_4015_2[1]));
    assign layer_3[955] = far_3_4015_2[0] | far_3_4015_2[1]; 
    wire [1:0] far_3_4016_0;    relay_conn far_3_4016_0_a(.in(layer_2[603]), .out(far_3_4016_0[0]));    relay_conn far_3_4016_0_b(.in(layer_2[714]), .out(far_3_4016_0[1]));
    wire [1:0] far_3_4016_1;    relay_conn far_3_4016_1_a(.in(far_3_4016_0[0]), .out(far_3_4016_1[0]));    relay_conn far_3_4016_1_b(.in(far_3_4016_0[1]), .out(far_3_4016_1[1]));
    wire [1:0] far_3_4016_2;    relay_conn far_3_4016_2_a(.in(far_3_4016_1[0]), .out(far_3_4016_2[0]));    relay_conn far_3_4016_2_b(.in(far_3_4016_1[1]), .out(far_3_4016_2[1]));
    assign layer_3[956] = ~far_3_4016_2[1] | (far_3_4016_2[0] & far_3_4016_2[1]); 
    wire [1:0] far_3_4017_0;    relay_conn far_3_4017_0_a(.in(layer_2[729]), .out(far_3_4017_0[0]));    relay_conn far_3_4017_0_b(.in(layer_2[645]), .out(far_3_4017_0[1]));
    wire [1:0] far_3_4017_1;    relay_conn far_3_4017_1_a(.in(far_3_4017_0[0]), .out(far_3_4017_1[0]));    relay_conn far_3_4017_1_b(.in(far_3_4017_0[1]), .out(far_3_4017_1[1]));
    assign layer_3[957] = far_3_4017_1[0] | far_3_4017_1[1]; 
    wire [1:0] far_3_4018_0;    relay_conn far_3_4018_0_a(.in(layer_2[710]), .out(far_3_4018_0[0]));    relay_conn far_3_4018_0_b(.in(layer_2[609]), .out(far_3_4018_0[1]));
    wire [1:0] far_3_4018_1;    relay_conn far_3_4018_1_a(.in(far_3_4018_0[0]), .out(far_3_4018_1[0]));    relay_conn far_3_4018_1_b(.in(far_3_4018_0[1]), .out(far_3_4018_1[1]));
    wire [1:0] far_3_4018_2;    relay_conn far_3_4018_2_a(.in(far_3_4018_1[0]), .out(far_3_4018_2[0]));    relay_conn far_3_4018_2_b(.in(far_3_4018_1[1]), .out(far_3_4018_2[1]));
    assign layer_3[958] = ~far_3_4018_2[1] | (far_3_4018_2[0] & far_3_4018_2[1]); 
    assign layer_3[959] = ~(layer_2[987] & layer_2[1012]); 
    wire [1:0] far_3_4020_0;    relay_conn far_3_4020_0_a(.in(layer_2[198]), .out(far_3_4020_0[0]));    relay_conn far_3_4020_0_b(.in(layer_2[126]), .out(far_3_4020_0[1]));
    wire [1:0] far_3_4020_1;    relay_conn far_3_4020_1_a(.in(far_3_4020_0[0]), .out(far_3_4020_1[0]));    relay_conn far_3_4020_1_b(.in(far_3_4020_0[1]), .out(far_3_4020_1[1]));
    assign layer_3[960] = far_3_4020_1[0] & ~far_3_4020_1[1]; 
    wire [1:0] far_3_4021_0;    relay_conn far_3_4021_0_a(.in(layer_2[783]), .out(far_3_4021_0[0]));    relay_conn far_3_4021_0_b(.in(layer_2[680]), .out(far_3_4021_0[1]));
    wire [1:0] far_3_4021_1;    relay_conn far_3_4021_1_a(.in(far_3_4021_0[0]), .out(far_3_4021_1[0]));    relay_conn far_3_4021_1_b(.in(far_3_4021_0[1]), .out(far_3_4021_1[1]));
    wire [1:0] far_3_4021_2;    relay_conn far_3_4021_2_a(.in(far_3_4021_1[0]), .out(far_3_4021_2[0]));    relay_conn far_3_4021_2_b(.in(far_3_4021_1[1]), .out(far_3_4021_2[1]));
    assign layer_3[961] = far_3_4021_2[1] & ~far_3_4021_2[0]; 
    wire [1:0] far_3_4022_0;    relay_conn far_3_4022_0_a(.in(layer_2[304]), .out(far_3_4022_0[0]));    relay_conn far_3_4022_0_b(.in(layer_2[390]), .out(far_3_4022_0[1]));
    wire [1:0] far_3_4022_1;    relay_conn far_3_4022_1_a(.in(far_3_4022_0[0]), .out(far_3_4022_1[0]));    relay_conn far_3_4022_1_b(.in(far_3_4022_0[1]), .out(far_3_4022_1[1]));
    assign layer_3[962] = far_3_4022_1[0] ^ far_3_4022_1[1]; 
    wire [1:0] far_3_4023_0;    relay_conn far_3_4023_0_a(.in(layer_2[794]), .out(far_3_4023_0[0]));    relay_conn far_3_4023_0_b(.in(layer_2[706]), .out(far_3_4023_0[1]));
    wire [1:0] far_3_4023_1;    relay_conn far_3_4023_1_a(.in(far_3_4023_0[0]), .out(far_3_4023_1[0]));    relay_conn far_3_4023_1_b(.in(far_3_4023_0[1]), .out(far_3_4023_1[1]));
    assign layer_3[963] = ~far_3_4023_1[0] | (far_3_4023_1[0] & far_3_4023_1[1]); 
    wire [1:0] far_3_4024_0;    relay_conn far_3_4024_0_a(.in(layer_2[950]), .out(far_3_4024_0[0]));    relay_conn far_3_4024_0_b(.in(layer_2[822]), .out(far_3_4024_0[1]));
    wire [1:0] far_3_4024_1;    relay_conn far_3_4024_1_a(.in(far_3_4024_0[0]), .out(far_3_4024_1[0]));    relay_conn far_3_4024_1_b(.in(far_3_4024_0[1]), .out(far_3_4024_1[1]));
    wire [1:0] far_3_4024_2;    relay_conn far_3_4024_2_a(.in(far_3_4024_1[0]), .out(far_3_4024_2[0]));    relay_conn far_3_4024_2_b(.in(far_3_4024_1[1]), .out(far_3_4024_2[1]));
    wire [1:0] far_3_4024_3;    relay_conn far_3_4024_3_a(.in(far_3_4024_2[0]), .out(far_3_4024_3[0]));    relay_conn far_3_4024_3_b(.in(far_3_4024_2[1]), .out(far_3_4024_3[1]));
    assign layer_3[964] = ~far_3_4024_3[1] | (far_3_4024_3[0] & far_3_4024_3[1]); 
    assign layer_3[965] = layer_2[700] | layer_2[712]; 
    wire [1:0] far_3_4026_0;    relay_conn far_3_4026_0_a(.in(layer_2[181]), .out(far_3_4026_0[0]));    relay_conn far_3_4026_0_b(.in(layer_2[112]), .out(far_3_4026_0[1]));
    wire [1:0] far_3_4026_1;    relay_conn far_3_4026_1_a(.in(far_3_4026_0[0]), .out(far_3_4026_1[0]));    relay_conn far_3_4026_1_b(.in(far_3_4026_0[1]), .out(far_3_4026_1[1]));
    assign layer_3[966] = far_3_4026_1[0] ^ far_3_4026_1[1]; 
    wire [1:0] far_3_4027_0;    relay_conn far_3_4027_0_a(.in(layer_2[178]), .out(far_3_4027_0[0]));    relay_conn far_3_4027_0_b(.in(layer_2[58]), .out(far_3_4027_0[1]));
    wire [1:0] far_3_4027_1;    relay_conn far_3_4027_1_a(.in(far_3_4027_0[0]), .out(far_3_4027_1[0]));    relay_conn far_3_4027_1_b(.in(far_3_4027_0[1]), .out(far_3_4027_1[1]));
    wire [1:0] far_3_4027_2;    relay_conn far_3_4027_2_a(.in(far_3_4027_1[0]), .out(far_3_4027_2[0]));    relay_conn far_3_4027_2_b(.in(far_3_4027_1[1]), .out(far_3_4027_2[1]));
    assign layer_3[967] = far_3_4027_2[1] & ~far_3_4027_2[0]; 
    assign layer_3[968] = ~(layer_2[916] | layer_2[888]); 
    wire [1:0] far_3_4029_0;    relay_conn far_3_4029_0_a(.in(layer_2[849]), .out(far_3_4029_0[0]));    relay_conn far_3_4029_0_b(.in(layer_2[813]), .out(far_3_4029_0[1]));
    assign layer_3[969] = far_3_4029_0[1] & ~far_3_4029_0[0]; 
    wire [1:0] far_3_4030_0;    relay_conn far_3_4030_0_a(.in(layer_2[324]), .out(far_3_4030_0[0]));    relay_conn far_3_4030_0_b(.in(layer_2[389]), .out(far_3_4030_0[1]));
    wire [1:0] far_3_4030_1;    relay_conn far_3_4030_1_a(.in(far_3_4030_0[0]), .out(far_3_4030_1[0]));    relay_conn far_3_4030_1_b(.in(far_3_4030_0[1]), .out(far_3_4030_1[1]));
    assign layer_3[970] = far_3_4030_1[0] & far_3_4030_1[1]; 
    wire [1:0] far_3_4031_0;    relay_conn far_3_4031_0_a(.in(layer_2[186]), .out(far_3_4031_0[0]));    relay_conn far_3_4031_0_b(.in(layer_2[151]), .out(far_3_4031_0[1]));
    assign layer_3[971] = ~(far_3_4031_0[0] | far_3_4031_0[1]); 
    wire [1:0] far_3_4032_0;    relay_conn far_3_4032_0_a(.in(layer_2[221]), .out(far_3_4032_0[0]));    relay_conn far_3_4032_0_b(.in(layer_2[120]), .out(far_3_4032_0[1]));
    wire [1:0] far_3_4032_1;    relay_conn far_3_4032_1_a(.in(far_3_4032_0[0]), .out(far_3_4032_1[0]));    relay_conn far_3_4032_1_b(.in(far_3_4032_0[1]), .out(far_3_4032_1[1]));
    wire [1:0] far_3_4032_2;    relay_conn far_3_4032_2_a(.in(far_3_4032_1[0]), .out(far_3_4032_2[0]));    relay_conn far_3_4032_2_b(.in(far_3_4032_1[1]), .out(far_3_4032_2[1]));
    assign layer_3[972] = ~far_3_4032_2[1] | (far_3_4032_2[0] & far_3_4032_2[1]); 
    wire [1:0] far_3_4033_0;    relay_conn far_3_4033_0_a(.in(layer_2[398]), .out(far_3_4033_0[0]));    relay_conn far_3_4033_0_b(.in(layer_2[292]), .out(far_3_4033_0[1]));
    wire [1:0] far_3_4033_1;    relay_conn far_3_4033_1_a(.in(far_3_4033_0[0]), .out(far_3_4033_1[0]));    relay_conn far_3_4033_1_b(.in(far_3_4033_0[1]), .out(far_3_4033_1[1]));
    wire [1:0] far_3_4033_2;    relay_conn far_3_4033_2_a(.in(far_3_4033_1[0]), .out(far_3_4033_2[0]));    relay_conn far_3_4033_2_b(.in(far_3_4033_1[1]), .out(far_3_4033_2[1]));
    assign layer_3[973] = ~far_3_4033_2[0]; 
    wire [1:0] far_3_4034_0;    relay_conn far_3_4034_0_a(.in(layer_2[957]), .out(far_3_4034_0[0]));    relay_conn far_3_4034_0_b(.in(layer_2[891]), .out(far_3_4034_0[1]));
    wire [1:0] far_3_4034_1;    relay_conn far_3_4034_1_a(.in(far_3_4034_0[0]), .out(far_3_4034_1[0]));    relay_conn far_3_4034_1_b(.in(far_3_4034_0[1]), .out(far_3_4034_1[1]));
    assign layer_3[974] = ~(far_3_4034_1[0] & far_3_4034_1[1]); 
    assign layer_3[975] = layer_2[927] | layer_2[946]; 
    assign layer_3[976] = ~(layer_2[462] & layer_2[483]); 
    wire [1:0] far_3_4037_0;    relay_conn far_3_4037_0_a(.in(layer_2[965]), .out(far_3_4037_0[0]));    relay_conn far_3_4037_0_b(.in(layer_2[839]), .out(far_3_4037_0[1]));
    wire [1:0] far_3_4037_1;    relay_conn far_3_4037_1_a(.in(far_3_4037_0[0]), .out(far_3_4037_1[0]));    relay_conn far_3_4037_1_b(.in(far_3_4037_0[1]), .out(far_3_4037_1[1]));
    wire [1:0] far_3_4037_2;    relay_conn far_3_4037_2_a(.in(far_3_4037_1[0]), .out(far_3_4037_2[0]));    relay_conn far_3_4037_2_b(.in(far_3_4037_1[1]), .out(far_3_4037_2[1]));
    assign layer_3[977] = far_3_4037_2[0]; 
    assign layer_3[978] = layer_2[370] & layer_2[343]; 
    wire [1:0] far_3_4039_0;    relay_conn far_3_4039_0_a(.in(layer_2[986]), .out(far_3_4039_0[0]));    relay_conn far_3_4039_0_b(.in(layer_2[915]), .out(far_3_4039_0[1]));
    wire [1:0] far_3_4039_1;    relay_conn far_3_4039_1_a(.in(far_3_4039_0[0]), .out(far_3_4039_1[0]));    relay_conn far_3_4039_1_b(.in(far_3_4039_0[1]), .out(far_3_4039_1[1]));
    assign layer_3[979] = far_3_4039_1[0] & ~far_3_4039_1[1]; 
    wire [1:0] far_3_4040_0;    relay_conn far_3_4040_0_a(.in(layer_2[962]), .out(far_3_4040_0[0]));    relay_conn far_3_4040_0_b(.in(layer_2[872]), .out(far_3_4040_0[1]));
    wire [1:0] far_3_4040_1;    relay_conn far_3_4040_1_a(.in(far_3_4040_0[0]), .out(far_3_4040_1[0]));    relay_conn far_3_4040_1_b(.in(far_3_4040_0[1]), .out(far_3_4040_1[1]));
    assign layer_3[980] = ~(far_3_4040_1[0] | far_3_4040_1[1]); 
    assign layer_3[981] = layer_2[206] ^ layer_2[191]; 
    wire [1:0] far_3_4042_0;    relay_conn far_3_4042_0_a(.in(layer_2[774]), .out(far_3_4042_0[0]));    relay_conn far_3_4042_0_b(.in(layer_2[821]), .out(far_3_4042_0[1]));
    assign layer_3[982] = far_3_4042_0[1]; 
    assign layer_3[983] = layer_2[43] & ~layer_2[67]; 
    wire [1:0] far_3_4044_0;    relay_conn far_3_4044_0_a(.in(layer_2[779]), .out(far_3_4044_0[0]));    relay_conn far_3_4044_0_b(.in(layer_2[735]), .out(far_3_4044_0[1]));
    assign layer_3[984] = far_3_4044_0[0] | far_3_4044_0[1]; 
    assign layer_3[985] = layer_2[989] | layer_2[965]; 
    assign layer_3[986] = layer_2[738]; 
    wire [1:0] far_3_4047_0;    relay_conn far_3_4047_0_a(.in(layer_2[218]), .out(far_3_4047_0[0]));    relay_conn far_3_4047_0_b(.in(layer_2[299]), .out(far_3_4047_0[1]));
    wire [1:0] far_3_4047_1;    relay_conn far_3_4047_1_a(.in(far_3_4047_0[0]), .out(far_3_4047_1[0]));    relay_conn far_3_4047_1_b(.in(far_3_4047_0[1]), .out(far_3_4047_1[1]));
    assign layer_3[987] = far_3_4047_1[0] | far_3_4047_1[1]; 
    wire [1:0] far_3_4048_0;    relay_conn far_3_4048_0_a(.in(layer_2[849]), .out(far_3_4048_0[0]));    relay_conn far_3_4048_0_b(.in(layer_2[907]), .out(far_3_4048_0[1]));
    assign layer_3[988] = ~far_3_4048_0[0]; 
    wire [1:0] far_3_4049_0;    relay_conn far_3_4049_0_a(.in(layer_2[661]), .out(far_3_4049_0[0]));    relay_conn far_3_4049_0_b(.in(layer_2[695]), .out(far_3_4049_0[1]));
    assign layer_3[989] = far_3_4049_0[0] | far_3_4049_0[1]; 
    wire [1:0] far_3_4050_0;    relay_conn far_3_4050_0_a(.in(layer_2[592]), .out(far_3_4050_0[0]));    relay_conn far_3_4050_0_b(.in(layer_2[674]), .out(far_3_4050_0[1]));
    wire [1:0] far_3_4050_1;    relay_conn far_3_4050_1_a(.in(far_3_4050_0[0]), .out(far_3_4050_1[0]));    relay_conn far_3_4050_1_b(.in(far_3_4050_0[1]), .out(far_3_4050_1[1]));
    assign layer_3[990] = far_3_4050_1[0] | far_3_4050_1[1]; 
    wire [1:0] far_3_4051_0;    relay_conn far_3_4051_0_a(.in(layer_2[732]), .out(far_3_4051_0[0]));    relay_conn far_3_4051_0_b(.in(layer_2[664]), .out(far_3_4051_0[1]));
    wire [1:0] far_3_4051_1;    relay_conn far_3_4051_1_a(.in(far_3_4051_0[0]), .out(far_3_4051_1[0]));    relay_conn far_3_4051_1_b(.in(far_3_4051_0[1]), .out(far_3_4051_1[1]));
    assign layer_3[991] = far_3_4051_1[1] & ~far_3_4051_1[0]; 
    wire [1:0] far_3_4052_0;    relay_conn far_3_4052_0_a(.in(layer_2[313]), .out(far_3_4052_0[0]));    relay_conn far_3_4052_0_b(.in(layer_2[265]), .out(far_3_4052_0[1]));
    assign layer_3[992] = far_3_4052_0[0] & far_3_4052_0[1]; 
    wire [1:0] far_3_4053_0;    relay_conn far_3_4053_0_a(.in(layer_2[100]), .out(far_3_4053_0[0]));    relay_conn far_3_4053_0_b(.in(layer_2[134]), .out(far_3_4053_0[1]));
    assign layer_3[993] = ~(far_3_4053_0[0] ^ far_3_4053_0[1]); 
    wire [1:0] far_3_4054_0;    relay_conn far_3_4054_0_a(.in(layer_2[306]), .out(far_3_4054_0[0]));    relay_conn far_3_4054_0_b(.in(layer_2[401]), .out(far_3_4054_0[1]));
    wire [1:0] far_3_4054_1;    relay_conn far_3_4054_1_a(.in(far_3_4054_0[0]), .out(far_3_4054_1[0]));    relay_conn far_3_4054_1_b(.in(far_3_4054_0[1]), .out(far_3_4054_1[1]));
    assign layer_3[994] = ~far_3_4054_1[1] | (far_3_4054_1[0] & far_3_4054_1[1]); 
    wire [1:0] far_3_4055_0;    relay_conn far_3_4055_0_a(.in(layer_2[903]), .out(far_3_4055_0[0]));    relay_conn far_3_4055_0_b(.in(layer_2[954]), .out(far_3_4055_0[1]));
    assign layer_3[995] = ~far_3_4055_0[0]; 
    assign layer_3[996] = ~(layer_2[854] | layer_2[880]); 
    assign layer_3[997] = ~(layer_2[247] & layer_2[265]); 
    assign layer_3[998] = ~(layer_2[57] | layer_2[58]); 
    wire [1:0] far_3_4059_0;    relay_conn far_3_4059_0_a(.in(layer_2[201]), .out(far_3_4059_0[0]));    relay_conn far_3_4059_0_b(.in(layer_2[132]), .out(far_3_4059_0[1]));
    wire [1:0] far_3_4059_1;    relay_conn far_3_4059_1_a(.in(far_3_4059_0[0]), .out(far_3_4059_1[0]));    relay_conn far_3_4059_1_b(.in(far_3_4059_0[1]), .out(far_3_4059_1[1]));
    assign layer_3[999] = ~(far_3_4059_1[0] ^ far_3_4059_1[1]); 
    wire [1:0] far_3_4060_0;    relay_conn far_3_4060_0_a(.in(layer_2[514]), .out(far_3_4060_0[0]));    relay_conn far_3_4060_0_b(.in(layer_2[435]), .out(far_3_4060_0[1]));
    wire [1:0] far_3_4060_1;    relay_conn far_3_4060_1_a(.in(far_3_4060_0[0]), .out(far_3_4060_1[0]));    relay_conn far_3_4060_1_b(.in(far_3_4060_0[1]), .out(far_3_4060_1[1]));
    assign layer_3[1000] = far_3_4060_1[0] & ~far_3_4060_1[1]; 
    wire [1:0] far_3_4061_0;    relay_conn far_3_4061_0_a(.in(layer_2[433]), .out(far_3_4061_0[0]));    relay_conn far_3_4061_0_b(.in(layer_2[546]), .out(far_3_4061_0[1]));
    wire [1:0] far_3_4061_1;    relay_conn far_3_4061_1_a(.in(far_3_4061_0[0]), .out(far_3_4061_1[0]));    relay_conn far_3_4061_1_b(.in(far_3_4061_0[1]), .out(far_3_4061_1[1]));
    wire [1:0] far_3_4061_2;    relay_conn far_3_4061_2_a(.in(far_3_4061_1[0]), .out(far_3_4061_2[0]));    relay_conn far_3_4061_2_b(.in(far_3_4061_1[1]), .out(far_3_4061_2[1]));
    assign layer_3[1001] = ~far_3_4061_2[1] | (far_3_4061_2[0] & far_3_4061_2[1]); 
    wire [1:0] far_3_4062_0;    relay_conn far_3_4062_0_a(.in(layer_2[354]), .out(far_3_4062_0[0]));    relay_conn far_3_4062_0_b(.in(layer_2[271]), .out(far_3_4062_0[1]));
    wire [1:0] far_3_4062_1;    relay_conn far_3_4062_1_a(.in(far_3_4062_0[0]), .out(far_3_4062_1[0]));    relay_conn far_3_4062_1_b(.in(far_3_4062_0[1]), .out(far_3_4062_1[1]));
    assign layer_3[1002] = far_3_4062_1[1]; 
    wire [1:0] far_3_4063_0;    relay_conn far_3_4063_0_a(.in(layer_2[327]), .out(far_3_4063_0[0]));    relay_conn far_3_4063_0_b(.in(layer_2[208]), .out(far_3_4063_0[1]));
    wire [1:0] far_3_4063_1;    relay_conn far_3_4063_1_a(.in(far_3_4063_0[0]), .out(far_3_4063_1[0]));    relay_conn far_3_4063_1_b(.in(far_3_4063_0[1]), .out(far_3_4063_1[1]));
    wire [1:0] far_3_4063_2;    relay_conn far_3_4063_2_a(.in(far_3_4063_1[0]), .out(far_3_4063_2[0]));    relay_conn far_3_4063_2_b(.in(far_3_4063_1[1]), .out(far_3_4063_2[1]));
    assign layer_3[1003] = ~(far_3_4063_2[0] | far_3_4063_2[1]); 
    assign layer_3[1004] = layer_2[1005] & ~layer_2[975]; 
    wire [1:0] far_3_4065_0;    relay_conn far_3_4065_0_a(.in(layer_2[161]), .out(far_3_4065_0[0]));    relay_conn far_3_4065_0_b(.in(layer_2[211]), .out(far_3_4065_0[1]));
    assign layer_3[1005] = far_3_4065_0[0] & ~far_3_4065_0[1]; 
    wire [1:0] far_3_4066_0;    relay_conn far_3_4066_0_a(.in(layer_2[339]), .out(far_3_4066_0[0]));    relay_conn far_3_4066_0_b(.in(layer_2[225]), .out(far_3_4066_0[1]));
    wire [1:0] far_3_4066_1;    relay_conn far_3_4066_1_a(.in(far_3_4066_0[0]), .out(far_3_4066_1[0]));    relay_conn far_3_4066_1_b(.in(far_3_4066_0[1]), .out(far_3_4066_1[1]));
    wire [1:0] far_3_4066_2;    relay_conn far_3_4066_2_a(.in(far_3_4066_1[0]), .out(far_3_4066_2[0]));    relay_conn far_3_4066_2_b(.in(far_3_4066_1[1]), .out(far_3_4066_2[1]));
    assign layer_3[1006] = far_3_4066_2[0] & far_3_4066_2[1]; 
    wire [1:0] far_3_4067_0;    relay_conn far_3_4067_0_a(.in(layer_2[178]), .out(far_3_4067_0[0]));    relay_conn far_3_4067_0_b(.in(layer_2[265]), .out(far_3_4067_0[1]));
    wire [1:0] far_3_4067_1;    relay_conn far_3_4067_1_a(.in(far_3_4067_0[0]), .out(far_3_4067_1[0]));    relay_conn far_3_4067_1_b(.in(far_3_4067_0[1]), .out(far_3_4067_1[1]));
    assign layer_3[1007] = far_3_4067_1[1] & ~far_3_4067_1[0]; 
    assign layer_3[1008] = layer_2[554] | layer_2[572]; 
    wire [1:0] far_3_4069_0;    relay_conn far_3_4069_0_a(.in(layer_2[525]), .out(far_3_4069_0[0]));    relay_conn far_3_4069_0_b(.in(layer_2[640]), .out(far_3_4069_0[1]));
    wire [1:0] far_3_4069_1;    relay_conn far_3_4069_1_a(.in(far_3_4069_0[0]), .out(far_3_4069_1[0]));    relay_conn far_3_4069_1_b(.in(far_3_4069_0[1]), .out(far_3_4069_1[1]));
    wire [1:0] far_3_4069_2;    relay_conn far_3_4069_2_a(.in(far_3_4069_1[0]), .out(far_3_4069_2[0]));    relay_conn far_3_4069_2_b(.in(far_3_4069_1[1]), .out(far_3_4069_2[1]));
    assign layer_3[1009] = ~far_3_4069_2[0]; 
    wire [1:0] far_3_4070_0;    relay_conn far_3_4070_0_a(.in(layer_2[324]), .out(far_3_4070_0[0]));    relay_conn far_3_4070_0_b(.in(layer_2[366]), .out(far_3_4070_0[1]));
    assign layer_3[1010] = ~far_3_4070_0[0]; 
    wire [1:0] far_3_4071_0;    relay_conn far_3_4071_0_a(.in(layer_2[508]), .out(far_3_4071_0[0]));    relay_conn far_3_4071_0_b(.in(layer_2[398]), .out(far_3_4071_0[1]));
    wire [1:0] far_3_4071_1;    relay_conn far_3_4071_1_a(.in(far_3_4071_0[0]), .out(far_3_4071_1[0]));    relay_conn far_3_4071_1_b(.in(far_3_4071_0[1]), .out(far_3_4071_1[1]));
    wire [1:0] far_3_4071_2;    relay_conn far_3_4071_2_a(.in(far_3_4071_1[0]), .out(far_3_4071_2[0]));    relay_conn far_3_4071_2_b(.in(far_3_4071_1[1]), .out(far_3_4071_2[1]));
    assign layer_3[1011] = ~far_3_4071_2[1] | (far_3_4071_2[0] & far_3_4071_2[1]); 
    wire [1:0] far_3_4072_0;    relay_conn far_3_4072_0_a(.in(layer_2[471]), .out(far_3_4072_0[0]));    relay_conn far_3_4072_0_b(.in(layer_2[430]), .out(far_3_4072_0[1]));
    assign layer_3[1012] = far_3_4072_0[1] & ~far_3_4072_0[0]; 
    wire [1:0] far_3_4073_0;    relay_conn far_3_4073_0_a(.in(layer_2[740]), .out(far_3_4073_0[0]));    relay_conn far_3_4073_0_b(.in(layer_2[781]), .out(far_3_4073_0[1]));
    assign layer_3[1013] = ~(far_3_4073_0[0] ^ far_3_4073_0[1]); 
    wire [1:0] far_3_4074_0;    relay_conn far_3_4074_0_a(.in(layer_2[133]), .out(far_3_4074_0[0]));    relay_conn far_3_4074_0_b(.in(layer_2[18]), .out(far_3_4074_0[1]));
    wire [1:0] far_3_4074_1;    relay_conn far_3_4074_1_a(.in(far_3_4074_0[0]), .out(far_3_4074_1[0]));    relay_conn far_3_4074_1_b(.in(far_3_4074_0[1]), .out(far_3_4074_1[1]));
    wire [1:0] far_3_4074_2;    relay_conn far_3_4074_2_a(.in(far_3_4074_1[0]), .out(far_3_4074_2[0]));    relay_conn far_3_4074_2_b(.in(far_3_4074_1[1]), .out(far_3_4074_2[1]));
    assign layer_3[1014] = ~far_3_4074_2[1]; 
    wire [1:0] far_3_4075_0;    relay_conn far_3_4075_0_a(.in(layer_2[25]), .out(far_3_4075_0[0]));    relay_conn far_3_4075_0_b(.in(layer_2[126]), .out(far_3_4075_0[1]));
    wire [1:0] far_3_4075_1;    relay_conn far_3_4075_1_a(.in(far_3_4075_0[0]), .out(far_3_4075_1[0]));    relay_conn far_3_4075_1_b(.in(far_3_4075_0[1]), .out(far_3_4075_1[1]));
    wire [1:0] far_3_4075_2;    relay_conn far_3_4075_2_a(.in(far_3_4075_1[0]), .out(far_3_4075_2[0]));    relay_conn far_3_4075_2_b(.in(far_3_4075_1[1]), .out(far_3_4075_2[1]));
    assign layer_3[1015] = ~(far_3_4075_2[0] & far_3_4075_2[1]); 
    wire [1:0] far_3_4076_0;    relay_conn far_3_4076_0_a(.in(layer_2[800]), .out(far_3_4076_0[0]));    relay_conn far_3_4076_0_b(.in(layer_2[698]), .out(far_3_4076_0[1]));
    wire [1:0] far_3_4076_1;    relay_conn far_3_4076_1_a(.in(far_3_4076_0[0]), .out(far_3_4076_1[0]));    relay_conn far_3_4076_1_b(.in(far_3_4076_0[1]), .out(far_3_4076_1[1]));
    wire [1:0] far_3_4076_2;    relay_conn far_3_4076_2_a(.in(far_3_4076_1[0]), .out(far_3_4076_2[0]));    relay_conn far_3_4076_2_b(.in(far_3_4076_1[1]), .out(far_3_4076_2[1]));
    assign layer_3[1016] = far_3_4076_2[1]; 
    wire [1:0] far_3_4077_0;    relay_conn far_3_4077_0_a(.in(layer_2[695]), .out(far_3_4077_0[0]));    relay_conn far_3_4077_0_b(.in(layer_2[575]), .out(far_3_4077_0[1]));
    wire [1:0] far_3_4077_1;    relay_conn far_3_4077_1_a(.in(far_3_4077_0[0]), .out(far_3_4077_1[0]));    relay_conn far_3_4077_1_b(.in(far_3_4077_0[1]), .out(far_3_4077_1[1]));
    wire [1:0] far_3_4077_2;    relay_conn far_3_4077_2_a(.in(far_3_4077_1[0]), .out(far_3_4077_2[0]));    relay_conn far_3_4077_2_b(.in(far_3_4077_1[1]), .out(far_3_4077_2[1]));
    assign layer_3[1017] = far_3_4077_2[0] | far_3_4077_2[1]; 
    wire [1:0] far_3_4078_0;    relay_conn far_3_4078_0_a(.in(layer_2[424]), .out(far_3_4078_0[0]));    relay_conn far_3_4078_0_b(.in(layer_2[512]), .out(far_3_4078_0[1]));
    wire [1:0] far_3_4078_1;    relay_conn far_3_4078_1_a(.in(far_3_4078_0[0]), .out(far_3_4078_1[0]));    relay_conn far_3_4078_1_b(.in(far_3_4078_0[1]), .out(far_3_4078_1[1]));
    assign layer_3[1018] = far_3_4078_1[1] & ~far_3_4078_1[0]; 
    wire [1:0] far_3_4079_0;    relay_conn far_3_4079_0_a(.in(layer_2[191]), .out(far_3_4079_0[0]));    relay_conn far_3_4079_0_b(.in(layer_2[272]), .out(far_3_4079_0[1]));
    wire [1:0] far_3_4079_1;    relay_conn far_3_4079_1_a(.in(far_3_4079_0[0]), .out(far_3_4079_1[0]));    relay_conn far_3_4079_1_b(.in(far_3_4079_0[1]), .out(far_3_4079_1[1]));
    assign layer_3[1019] = ~far_3_4079_1[0] | (far_3_4079_1[0] & far_3_4079_1[1]); 
    // Layer 4 ============================================================
    assign layer_4[0] = layer_3[21] | layer_3[52]; 
    assign layer_4[1] = ~(layer_3[860] | layer_3[834]); 
    wire [1:0] far_4_4082_0;    relay_conn far_4_4082_0_a(.in(layer_3[619]), .out(far_4_4082_0[0]));    relay_conn far_4_4082_0_b(.in(layer_3[739]), .out(far_4_4082_0[1]));
    wire [1:0] far_4_4082_1;    relay_conn far_4_4082_1_a(.in(far_4_4082_0[0]), .out(far_4_4082_1[0]));    relay_conn far_4_4082_1_b(.in(far_4_4082_0[1]), .out(far_4_4082_1[1]));
    wire [1:0] far_4_4082_2;    relay_conn far_4_4082_2_a(.in(far_4_4082_1[0]), .out(far_4_4082_2[0]));    relay_conn far_4_4082_2_b(.in(far_4_4082_1[1]), .out(far_4_4082_2[1]));
    assign layer_4[2] = ~(far_4_4082_2[0] | far_4_4082_2[1]); 
    wire [1:0] far_4_4083_0;    relay_conn far_4_4083_0_a(.in(layer_3[75]), .out(far_4_4083_0[0]));    relay_conn far_4_4083_0_b(.in(layer_3[0]), .out(far_4_4083_0[1]));
    wire [1:0] far_4_4083_1;    relay_conn far_4_4083_1_a(.in(far_4_4083_0[0]), .out(far_4_4083_1[0]));    relay_conn far_4_4083_1_b(.in(far_4_4083_0[1]), .out(far_4_4083_1[1]));
    assign layer_4[3] = ~far_4_4083_1[0] | (far_4_4083_1[0] & far_4_4083_1[1]); 
    wire [1:0] far_4_4084_0;    relay_conn far_4_4084_0_a(.in(layer_3[633]), .out(far_4_4084_0[0]));    relay_conn far_4_4084_0_b(.in(layer_3[542]), .out(far_4_4084_0[1]));
    wire [1:0] far_4_4084_1;    relay_conn far_4_4084_1_a(.in(far_4_4084_0[0]), .out(far_4_4084_1[0]));    relay_conn far_4_4084_1_b(.in(far_4_4084_0[1]), .out(far_4_4084_1[1]));
    assign layer_4[4] = ~far_4_4084_1[0] | (far_4_4084_1[0] & far_4_4084_1[1]); 
    assign layer_4[5] = layer_3[922] & ~layer_3[953]; 
    wire [1:0] far_4_4086_0;    relay_conn far_4_4086_0_a(.in(layer_3[386]), .out(far_4_4086_0[0]));    relay_conn far_4_4086_0_b(.in(layer_3[507]), .out(far_4_4086_0[1]));
    wire [1:0] far_4_4086_1;    relay_conn far_4_4086_1_a(.in(far_4_4086_0[0]), .out(far_4_4086_1[0]));    relay_conn far_4_4086_1_b(.in(far_4_4086_0[1]), .out(far_4_4086_1[1]));
    wire [1:0] far_4_4086_2;    relay_conn far_4_4086_2_a(.in(far_4_4086_1[0]), .out(far_4_4086_2[0]));    relay_conn far_4_4086_2_b(.in(far_4_4086_1[1]), .out(far_4_4086_2[1]));
    assign layer_4[6] = ~(far_4_4086_2[0] & far_4_4086_2[1]); 
    wire [1:0] far_4_4087_0;    relay_conn far_4_4087_0_a(.in(layer_3[405]), .out(far_4_4087_0[0]));    relay_conn far_4_4087_0_b(.in(layer_3[318]), .out(far_4_4087_0[1]));
    wire [1:0] far_4_4087_1;    relay_conn far_4_4087_1_a(.in(far_4_4087_0[0]), .out(far_4_4087_1[0]));    relay_conn far_4_4087_1_b(.in(far_4_4087_0[1]), .out(far_4_4087_1[1]));
    assign layer_4[7] = far_4_4087_1[0]; 
    wire [1:0] far_4_4088_0;    relay_conn far_4_4088_0_a(.in(layer_3[782]), .out(far_4_4088_0[0]));    relay_conn far_4_4088_0_b(.in(layer_3[688]), .out(far_4_4088_0[1]));
    wire [1:0] far_4_4088_1;    relay_conn far_4_4088_1_a(.in(far_4_4088_0[0]), .out(far_4_4088_1[0]));    relay_conn far_4_4088_1_b(.in(far_4_4088_0[1]), .out(far_4_4088_1[1]));
    assign layer_4[8] = far_4_4088_1[1]; 
    wire [1:0] far_4_4089_0;    relay_conn far_4_4089_0_a(.in(layer_3[220]), .out(far_4_4089_0[0]));    relay_conn far_4_4089_0_b(.in(layer_3[112]), .out(far_4_4089_0[1]));
    wire [1:0] far_4_4089_1;    relay_conn far_4_4089_1_a(.in(far_4_4089_0[0]), .out(far_4_4089_1[0]));    relay_conn far_4_4089_1_b(.in(far_4_4089_0[1]), .out(far_4_4089_1[1]));
    wire [1:0] far_4_4089_2;    relay_conn far_4_4089_2_a(.in(far_4_4089_1[0]), .out(far_4_4089_2[0]));    relay_conn far_4_4089_2_b(.in(far_4_4089_1[1]), .out(far_4_4089_2[1]));
    assign layer_4[9] = ~far_4_4089_2[0] | (far_4_4089_2[0] & far_4_4089_2[1]); 
    wire [1:0] far_4_4090_0;    relay_conn far_4_4090_0_a(.in(layer_3[65]), .out(far_4_4090_0[0]));    relay_conn far_4_4090_0_b(.in(layer_3[140]), .out(far_4_4090_0[1]));
    wire [1:0] far_4_4090_1;    relay_conn far_4_4090_1_a(.in(far_4_4090_0[0]), .out(far_4_4090_1[0]));    relay_conn far_4_4090_1_b(.in(far_4_4090_0[1]), .out(far_4_4090_1[1]));
    assign layer_4[10] = ~far_4_4090_1[1]; 
    wire [1:0] far_4_4091_0;    relay_conn far_4_4091_0_a(.in(layer_3[14]), .out(far_4_4091_0[0]));    relay_conn far_4_4091_0_b(.in(layer_3[113]), .out(far_4_4091_0[1]));
    wire [1:0] far_4_4091_1;    relay_conn far_4_4091_1_a(.in(far_4_4091_0[0]), .out(far_4_4091_1[0]));    relay_conn far_4_4091_1_b(.in(far_4_4091_0[1]), .out(far_4_4091_1[1]));
    wire [1:0] far_4_4091_2;    relay_conn far_4_4091_2_a(.in(far_4_4091_1[0]), .out(far_4_4091_2[0]));    relay_conn far_4_4091_2_b(.in(far_4_4091_1[1]), .out(far_4_4091_2[1]));
    assign layer_4[11] = far_4_4091_2[1] & ~far_4_4091_2[0]; 
    wire [1:0] far_4_4092_0;    relay_conn far_4_4092_0_a(.in(layer_3[626]), .out(far_4_4092_0[0]));    relay_conn far_4_4092_0_b(.in(layer_3[537]), .out(far_4_4092_0[1]));
    wire [1:0] far_4_4092_1;    relay_conn far_4_4092_1_a(.in(far_4_4092_0[0]), .out(far_4_4092_1[0]));    relay_conn far_4_4092_1_b(.in(far_4_4092_0[1]), .out(far_4_4092_1[1]));
    assign layer_4[12] = far_4_4092_1[0] | far_4_4092_1[1]; 
    wire [1:0] far_4_4093_0;    relay_conn far_4_4093_0_a(.in(layer_3[979]), .out(far_4_4093_0[0]));    relay_conn far_4_4093_0_b(.in(layer_3[876]), .out(far_4_4093_0[1]));
    wire [1:0] far_4_4093_1;    relay_conn far_4_4093_1_a(.in(far_4_4093_0[0]), .out(far_4_4093_1[0]));    relay_conn far_4_4093_1_b(.in(far_4_4093_0[1]), .out(far_4_4093_1[1]));
    wire [1:0] far_4_4093_2;    relay_conn far_4_4093_2_a(.in(far_4_4093_1[0]), .out(far_4_4093_2[0]));    relay_conn far_4_4093_2_b(.in(far_4_4093_1[1]), .out(far_4_4093_2[1]));
    assign layer_4[13] = far_4_4093_2[1]; 
    wire [1:0] far_4_4094_0;    relay_conn far_4_4094_0_a(.in(layer_3[597]), .out(far_4_4094_0[0]));    relay_conn far_4_4094_0_b(.in(layer_3[633]), .out(far_4_4094_0[1]));
    assign layer_4[14] = ~far_4_4094_0[1]; 
    wire [1:0] far_4_4095_0;    relay_conn far_4_4095_0_a(.in(layer_3[636]), .out(far_4_4095_0[0]));    relay_conn far_4_4095_0_b(.in(layer_3[583]), .out(far_4_4095_0[1]));
    assign layer_4[15] = ~far_4_4095_0[0] | (far_4_4095_0[0] & far_4_4095_0[1]); 
    assign layer_4[16] = layer_3[732] | layer_3[734]; 
    assign layer_4[17] = layer_3[345] & ~layer_3[318]; 
    wire [1:0] far_4_4098_0;    relay_conn far_4_4098_0_a(.in(layer_3[253]), .out(far_4_4098_0[0]));    relay_conn far_4_4098_0_b(.in(layer_3[130]), .out(far_4_4098_0[1]));
    wire [1:0] far_4_4098_1;    relay_conn far_4_4098_1_a(.in(far_4_4098_0[0]), .out(far_4_4098_1[0]));    relay_conn far_4_4098_1_b(.in(far_4_4098_0[1]), .out(far_4_4098_1[1]));
    wire [1:0] far_4_4098_2;    relay_conn far_4_4098_2_a(.in(far_4_4098_1[0]), .out(far_4_4098_2[0]));    relay_conn far_4_4098_2_b(.in(far_4_4098_1[1]), .out(far_4_4098_2[1]));
    assign layer_4[18] = far_4_4098_2[0] ^ far_4_4098_2[1]; 
    wire [1:0] far_4_4099_0;    relay_conn far_4_4099_0_a(.in(layer_3[35]), .out(far_4_4099_0[0]));    relay_conn far_4_4099_0_b(.in(layer_3[83]), .out(far_4_4099_0[1]));
    assign layer_4[19] = far_4_4099_0[1]; 
    assign layer_4[20] = ~(layer_3[586] | layer_3[570]); 
    wire [1:0] far_4_4101_0;    relay_conn far_4_4101_0_a(.in(layer_3[808]), .out(far_4_4101_0[0]));    relay_conn far_4_4101_0_b(.in(layer_3[731]), .out(far_4_4101_0[1]));
    wire [1:0] far_4_4101_1;    relay_conn far_4_4101_1_a(.in(far_4_4101_0[0]), .out(far_4_4101_1[0]));    relay_conn far_4_4101_1_b(.in(far_4_4101_0[1]), .out(far_4_4101_1[1]));
    assign layer_4[21] = far_4_4101_1[0] | far_4_4101_1[1]; 
    wire [1:0] far_4_4102_0;    relay_conn far_4_4102_0_a(.in(layer_3[312]), .out(far_4_4102_0[0]));    relay_conn far_4_4102_0_b(.in(layer_3[353]), .out(far_4_4102_0[1]));
    assign layer_4[22] = far_4_4102_0[1] & ~far_4_4102_0[0]; 
    wire [1:0] far_4_4103_0;    relay_conn far_4_4103_0_a(.in(layer_3[104]), .out(far_4_4103_0[0]));    relay_conn far_4_4103_0_b(.in(layer_3[2]), .out(far_4_4103_0[1]));
    wire [1:0] far_4_4103_1;    relay_conn far_4_4103_1_a(.in(far_4_4103_0[0]), .out(far_4_4103_1[0]));    relay_conn far_4_4103_1_b(.in(far_4_4103_0[1]), .out(far_4_4103_1[1]));
    wire [1:0] far_4_4103_2;    relay_conn far_4_4103_2_a(.in(far_4_4103_1[0]), .out(far_4_4103_2[0]));    relay_conn far_4_4103_2_b(.in(far_4_4103_1[1]), .out(far_4_4103_2[1]));
    assign layer_4[23] = far_4_4103_2[0] & ~far_4_4103_2[1]; 
    wire [1:0] far_4_4104_0;    relay_conn far_4_4104_0_a(.in(layer_3[807]), .out(far_4_4104_0[0]));    relay_conn far_4_4104_0_b(.in(layer_3[861]), .out(far_4_4104_0[1]));
    assign layer_4[24] = ~(far_4_4104_0[0] ^ far_4_4104_0[1]); 
    wire [1:0] far_4_4105_0;    relay_conn far_4_4105_0_a(.in(layer_3[840]), .out(far_4_4105_0[0]));    relay_conn far_4_4105_0_b(.in(layer_3[806]), .out(far_4_4105_0[1]));
    assign layer_4[25] = ~far_4_4105_0[1]; 
    wire [1:0] far_4_4106_0;    relay_conn far_4_4106_0_a(.in(layer_3[986]), .out(far_4_4106_0[0]));    relay_conn far_4_4106_0_b(.in(layer_3[909]), .out(far_4_4106_0[1]));
    wire [1:0] far_4_4106_1;    relay_conn far_4_4106_1_a(.in(far_4_4106_0[0]), .out(far_4_4106_1[0]));    relay_conn far_4_4106_1_b(.in(far_4_4106_0[1]), .out(far_4_4106_1[1]));
    assign layer_4[26] = far_4_4106_1[0] & far_4_4106_1[1]; 
    wire [1:0] far_4_4107_0;    relay_conn far_4_4107_0_a(.in(layer_3[466]), .out(far_4_4107_0[0]));    relay_conn far_4_4107_0_b(.in(layer_3[593]), .out(far_4_4107_0[1]));
    wire [1:0] far_4_4107_1;    relay_conn far_4_4107_1_a(.in(far_4_4107_0[0]), .out(far_4_4107_1[0]));    relay_conn far_4_4107_1_b(.in(far_4_4107_0[1]), .out(far_4_4107_1[1]));
    wire [1:0] far_4_4107_2;    relay_conn far_4_4107_2_a(.in(far_4_4107_1[0]), .out(far_4_4107_2[0]));    relay_conn far_4_4107_2_b(.in(far_4_4107_1[1]), .out(far_4_4107_2[1]));
    assign layer_4[27] = far_4_4107_2[0] ^ far_4_4107_2[1]; 
    wire [1:0] far_4_4108_0;    relay_conn far_4_4108_0_a(.in(layer_3[812]), .out(far_4_4108_0[0]));    relay_conn far_4_4108_0_b(.in(layer_3[688]), .out(far_4_4108_0[1]));
    wire [1:0] far_4_4108_1;    relay_conn far_4_4108_1_a(.in(far_4_4108_0[0]), .out(far_4_4108_1[0]));    relay_conn far_4_4108_1_b(.in(far_4_4108_0[1]), .out(far_4_4108_1[1]));
    wire [1:0] far_4_4108_2;    relay_conn far_4_4108_2_a(.in(far_4_4108_1[0]), .out(far_4_4108_2[0]));    relay_conn far_4_4108_2_b(.in(far_4_4108_1[1]), .out(far_4_4108_2[1]));
    assign layer_4[28] = far_4_4108_2[1] & ~far_4_4108_2[0]; 
    wire [1:0] far_4_4109_0;    relay_conn far_4_4109_0_a(.in(layer_3[507]), .out(far_4_4109_0[0]));    relay_conn far_4_4109_0_b(.in(layer_3[403]), .out(far_4_4109_0[1]));
    wire [1:0] far_4_4109_1;    relay_conn far_4_4109_1_a(.in(far_4_4109_0[0]), .out(far_4_4109_1[0]));    relay_conn far_4_4109_1_b(.in(far_4_4109_0[1]), .out(far_4_4109_1[1]));
    wire [1:0] far_4_4109_2;    relay_conn far_4_4109_2_a(.in(far_4_4109_1[0]), .out(far_4_4109_2[0]));    relay_conn far_4_4109_2_b(.in(far_4_4109_1[1]), .out(far_4_4109_2[1]));
    assign layer_4[29] = far_4_4109_2[0] | far_4_4109_2[1]; 
    wire [1:0] far_4_4110_0;    relay_conn far_4_4110_0_a(.in(layer_3[846]), .out(far_4_4110_0[0]));    relay_conn far_4_4110_0_b(.in(layer_3[936]), .out(far_4_4110_0[1]));
    wire [1:0] far_4_4110_1;    relay_conn far_4_4110_1_a(.in(far_4_4110_0[0]), .out(far_4_4110_1[0]));    relay_conn far_4_4110_1_b(.in(far_4_4110_0[1]), .out(far_4_4110_1[1]));
    assign layer_4[30] = ~far_4_4110_1[1] | (far_4_4110_1[0] & far_4_4110_1[1]); 
    assign layer_4[31] = ~(layer_3[47] ^ layer_3[30]); 
    assign layer_4[32] = ~(layer_3[9] ^ layer_3[32]); 
    wire [1:0] far_4_4113_0;    relay_conn far_4_4113_0_a(.in(layer_3[32]), .out(far_4_4113_0[0]));    relay_conn far_4_4113_0_b(.in(layer_3[105]), .out(far_4_4113_0[1]));
    wire [1:0] far_4_4113_1;    relay_conn far_4_4113_1_a(.in(far_4_4113_0[0]), .out(far_4_4113_1[0]));    relay_conn far_4_4113_1_b(.in(far_4_4113_0[1]), .out(far_4_4113_1[1]));
    assign layer_4[33] = far_4_4113_1[0] & far_4_4113_1[1]; 
    wire [1:0] far_4_4114_0;    relay_conn far_4_4114_0_a(.in(layer_3[13]), .out(far_4_4114_0[0]));    relay_conn far_4_4114_0_b(.in(layer_3[71]), .out(far_4_4114_0[1]));
    assign layer_4[34] = ~(far_4_4114_0[0] & far_4_4114_0[1]); 
    wire [1:0] far_4_4115_0;    relay_conn far_4_4115_0_a(.in(layer_3[1004]), .out(far_4_4115_0[0]));    relay_conn far_4_4115_0_b(.in(layer_3[957]), .out(far_4_4115_0[1]));
    assign layer_4[35] = far_4_4115_0[0] ^ far_4_4115_0[1]; 
    wire [1:0] far_4_4116_0;    relay_conn far_4_4116_0_a(.in(layer_3[958]), .out(far_4_4116_0[0]));    relay_conn far_4_4116_0_b(.in(layer_3[854]), .out(far_4_4116_0[1]));
    wire [1:0] far_4_4116_1;    relay_conn far_4_4116_1_a(.in(far_4_4116_0[0]), .out(far_4_4116_1[0]));    relay_conn far_4_4116_1_b(.in(far_4_4116_0[1]), .out(far_4_4116_1[1]));
    wire [1:0] far_4_4116_2;    relay_conn far_4_4116_2_a(.in(far_4_4116_1[0]), .out(far_4_4116_2[0]));    relay_conn far_4_4116_2_b(.in(far_4_4116_1[1]), .out(far_4_4116_2[1]));
    assign layer_4[36] = far_4_4116_2[0] & far_4_4116_2[1]; 
    assign layer_4[37] = ~(layer_3[431] & layer_3[410]); 
    wire [1:0] far_4_4118_0;    relay_conn far_4_4118_0_a(.in(layer_3[782]), .out(far_4_4118_0[0]));    relay_conn far_4_4118_0_b(.in(layer_3[878]), .out(far_4_4118_0[1]));
    wire [1:0] far_4_4118_1;    relay_conn far_4_4118_1_a(.in(far_4_4118_0[0]), .out(far_4_4118_1[0]));    relay_conn far_4_4118_1_b(.in(far_4_4118_0[1]), .out(far_4_4118_1[1]));
    wire [1:0] far_4_4118_2;    relay_conn far_4_4118_2_a(.in(far_4_4118_1[0]), .out(far_4_4118_2[0]));    relay_conn far_4_4118_2_b(.in(far_4_4118_1[1]), .out(far_4_4118_2[1]));
    assign layer_4[38] = ~far_4_4118_2[0] | (far_4_4118_2[0] & far_4_4118_2[1]); 
    assign layer_4[39] = layer_3[56] & layer_3[36]; 
    wire [1:0] far_4_4120_0;    relay_conn far_4_4120_0_a(.in(layer_3[192]), .out(far_4_4120_0[0]));    relay_conn far_4_4120_0_b(.in(layer_3[143]), .out(far_4_4120_0[1]));
    assign layer_4[40] = ~far_4_4120_0[0]; 
    wire [1:0] far_4_4121_0;    relay_conn far_4_4121_0_a(.in(layer_3[577]), .out(far_4_4121_0[0]));    relay_conn far_4_4121_0_b(.in(layer_3[543]), .out(far_4_4121_0[1]));
    assign layer_4[41] = ~far_4_4121_0[1] | (far_4_4121_0[0] & far_4_4121_0[1]); 
    assign layer_4[42] = layer_3[47] | layer_3[35]; 
    wire [1:0] far_4_4123_0;    relay_conn far_4_4123_0_a(.in(layer_3[905]), .out(far_4_4123_0[0]));    relay_conn far_4_4123_0_b(.in(layer_3[857]), .out(far_4_4123_0[1]));
    assign layer_4[43] = far_4_4123_0[0]; 
    wire [1:0] far_4_4124_0;    relay_conn far_4_4124_0_a(.in(layer_3[753]), .out(far_4_4124_0[0]));    relay_conn far_4_4124_0_b(.in(layer_3[877]), .out(far_4_4124_0[1]));
    wire [1:0] far_4_4124_1;    relay_conn far_4_4124_1_a(.in(far_4_4124_0[0]), .out(far_4_4124_1[0]));    relay_conn far_4_4124_1_b(.in(far_4_4124_0[1]), .out(far_4_4124_1[1]));
    wire [1:0] far_4_4124_2;    relay_conn far_4_4124_2_a(.in(far_4_4124_1[0]), .out(far_4_4124_2[0]));    relay_conn far_4_4124_2_b(.in(far_4_4124_1[1]), .out(far_4_4124_2[1]));
    assign layer_4[44] = ~far_4_4124_2[1]; 
    assign layer_4[45] = layer_3[854]; 
    assign layer_4[46] = layer_3[837]; 
    assign layer_4[47] = ~layer_3[419]; 
    wire [1:0] far_4_4128_0;    relay_conn far_4_4128_0_a(.in(layer_3[298]), .out(far_4_4128_0[0]));    relay_conn far_4_4128_0_b(.in(layer_3[211]), .out(far_4_4128_0[1]));
    wire [1:0] far_4_4128_1;    relay_conn far_4_4128_1_a(.in(far_4_4128_0[0]), .out(far_4_4128_1[0]));    relay_conn far_4_4128_1_b(.in(far_4_4128_0[1]), .out(far_4_4128_1[1]));
    assign layer_4[48] = far_4_4128_1[1] & ~far_4_4128_1[0]; 
    wire [1:0] far_4_4129_0;    relay_conn far_4_4129_0_a(.in(layer_3[664]), .out(far_4_4129_0[0]));    relay_conn far_4_4129_0_b(.in(layer_3[610]), .out(far_4_4129_0[1]));
    assign layer_4[49] = far_4_4129_0[0]; 
    wire [1:0] far_4_4130_0;    relay_conn far_4_4130_0_a(.in(layer_3[531]), .out(far_4_4130_0[0]));    relay_conn far_4_4130_0_b(.in(layer_3[424]), .out(far_4_4130_0[1]));
    wire [1:0] far_4_4130_1;    relay_conn far_4_4130_1_a(.in(far_4_4130_0[0]), .out(far_4_4130_1[0]));    relay_conn far_4_4130_1_b(.in(far_4_4130_0[1]), .out(far_4_4130_1[1]));
    wire [1:0] far_4_4130_2;    relay_conn far_4_4130_2_a(.in(far_4_4130_1[0]), .out(far_4_4130_2[0]));    relay_conn far_4_4130_2_b(.in(far_4_4130_1[1]), .out(far_4_4130_2[1]));
    assign layer_4[50] = ~far_4_4130_2[0]; 
    wire [1:0] far_4_4131_0;    relay_conn far_4_4131_0_a(.in(layer_3[1018]), .out(far_4_4131_0[0]));    relay_conn far_4_4131_0_b(.in(layer_3[972]), .out(far_4_4131_0[1]));
    assign layer_4[51] = ~far_4_4131_0[0] | (far_4_4131_0[0] & far_4_4131_0[1]); 
    wire [1:0] far_4_4132_0;    relay_conn far_4_4132_0_a(.in(layer_3[72]), .out(far_4_4132_0[0]));    relay_conn far_4_4132_0_b(.in(layer_3[30]), .out(far_4_4132_0[1]));
    assign layer_4[52] = far_4_4132_0[0] | far_4_4132_0[1]; 
    assign layer_4[53] = ~layer_3[455] | (layer_3[475] & layer_3[455]); 
    wire [1:0] far_4_4134_0;    relay_conn far_4_4134_0_a(.in(layer_3[5]), .out(far_4_4134_0[0]));    relay_conn far_4_4134_0_b(.in(layer_3[100]), .out(far_4_4134_0[1]));
    wire [1:0] far_4_4134_1;    relay_conn far_4_4134_1_a(.in(far_4_4134_0[0]), .out(far_4_4134_1[0]));    relay_conn far_4_4134_1_b(.in(far_4_4134_0[1]), .out(far_4_4134_1[1]));
    assign layer_4[54] = far_4_4134_1[0] | far_4_4134_1[1]; 
    wire [1:0] far_4_4135_0;    relay_conn far_4_4135_0_a(.in(layer_3[825]), .out(far_4_4135_0[0]));    relay_conn far_4_4135_0_b(.in(layer_3[731]), .out(far_4_4135_0[1]));
    wire [1:0] far_4_4135_1;    relay_conn far_4_4135_1_a(.in(far_4_4135_0[0]), .out(far_4_4135_1[0]));    relay_conn far_4_4135_1_b(.in(far_4_4135_0[1]), .out(far_4_4135_1[1]));
    assign layer_4[55] = far_4_4135_1[1]; 
    assign layer_4[56] = ~layer_3[869] | (layer_3[869] & layer_3[850]); 
    assign layer_4[57] = layer_3[969] & ~layer_3[992]; 
    wire [1:0] far_4_4138_0;    relay_conn far_4_4138_0_a(.in(layer_3[749]), .out(far_4_4138_0[0]));    relay_conn far_4_4138_0_b(.in(layer_3[843]), .out(far_4_4138_0[1]));
    wire [1:0] far_4_4138_1;    relay_conn far_4_4138_1_a(.in(far_4_4138_0[0]), .out(far_4_4138_1[0]));    relay_conn far_4_4138_1_b(.in(far_4_4138_0[1]), .out(far_4_4138_1[1]));
    assign layer_4[58] = ~far_4_4138_1[1]; 
    wire [1:0] far_4_4139_0;    relay_conn far_4_4139_0_a(.in(layer_3[402]), .out(far_4_4139_0[0]));    relay_conn far_4_4139_0_b(.in(layer_3[481]), .out(far_4_4139_0[1]));
    wire [1:0] far_4_4139_1;    relay_conn far_4_4139_1_a(.in(far_4_4139_0[0]), .out(far_4_4139_1[0]));    relay_conn far_4_4139_1_b(.in(far_4_4139_0[1]), .out(far_4_4139_1[1]));
    assign layer_4[59] = ~far_4_4139_1[1] | (far_4_4139_1[0] & far_4_4139_1[1]); 
    assign layer_4[60] = ~(layer_3[157] & layer_3[153]); 
    assign layer_4[61] = ~(layer_3[992] | layer_3[969]); 
    wire [1:0] far_4_4142_0;    relay_conn far_4_4142_0_a(.in(layer_3[34]), .out(far_4_4142_0[0]));    relay_conn far_4_4142_0_b(.in(layer_3[149]), .out(far_4_4142_0[1]));
    wire [1:0] far_4_4142_1;    relay_conn far_4_4142_1_a(.in(far_4_4142_0[0]), .out(far_4_4142_1[0]));    relay_conn far_4_4142_1_b(.in(far_4_4142_0[1]), .out(far_4_4142_1[1]));
    wire [1:0] far_4_4142_2;    relay_conn far_4_4142_2_a(.in(far_4_4142_1[0]), .out(far_4_4142_2[0]));    relay_conn far_4_4142_2_b(.in(far_4_4142_1[1]), .out(far_4_4142_2[1]));
    assign layer_4[62] = ~far_4_4142_2[1] | (far_4_4142_2[0] & far_4_4142_2[1]); 
    wire [1:0] far_4_4143_0;    relay_conn far_4_4143_0_a(.in(layer_3[816]), .out(far_4_4143_0[0]));    relay_conn far_4_4143_0_b(.in(layer_3[752]), .out(far_4_4143_0[1]));
    wire [1:0] far_4_4143_1;    relay_conn far_4_4143_1_a(.in(far_4_4143_0[0]), .out(far_4_4143_1[0]));    relay_conn far_4_4143_1_b(.in(far_4_4143_0[1]), .out(far_4_4143_1[1]));
    assign layer_4[63] = far_4_4143_1[0] & ~far_4_4143_1[1]; 
    wire [1:0] far_4_4144_0;    relay_conn far_4_4144_0_a(.in(layer_3[502]), .out(far_4_4144_0[0]));    relay_conn far_4_4144_0_b(.in(layer_3[570]), .out(far_4_4144_0[1]));
    wire [1:0] far_4_4144_1;    relay_conn far_4_4144_1_a(.in(far_4_4144_0[0]), .out(far_4_4144_1[0]));    relay_conn far_4_4144_1_b(.in(far_4_4144_0[1]), .out(far_4_4144_1[1]));
    assign layer_4[64] = far_4_4144_1[1] & ~far_4_4144_1[0]; 
    assign layer_4[65] = layer_3[312] | layer_3[288]; 
    wire [1:0] far_4_4146_0;    relay_conn far_4_4146_0_a(.in(layer_3[391]), .out(far_4_4146_0[0]));    relay_conn far_4_4146_0_b(.in(layer_3[501]), .out(far_4_4146_0[1]));
    wire [1:0] far_4_4146_1;    relay_conn far_4_4146_1_a(.in(far_4_4146_0[0]), .out(far_4_4146_1[0]));    relay_conn far_4_4146_1_b(.in(far_4_4146_0[1]), .out(far_4_4146_1[1]));
    wire [1:0] far_4_4146_2;    relay_conn far_4_4146_2_a(.in(far_4_4146_1[0]), .out(far_4_4146_2[0]));    relay_conn far_4_4146_2_b(.in(far_4_4146_1[1]), .out(far_4_4146_2[1]));
    assign layer_4[66] = far_4_4146_2[1] & ~far_4_4146_2[0]; 
    assign layer_4[67] = ~(layer_3[124] & layer_3[104]); 
    wire [1:0] far_4_4148_0;    relay_conn far_4_4148_0_a(.in(layer_3[433]), .out(far_4_4148_0[0]));    relay_conn far_4_4148_0_b(.in(layer_3[384]), .out(far_4_4148_0[1]));
    assign layer_4[68] = far_4_4148_0[0] ^ far_4_4148_0[1]; 
    wire [1:0] far_4_4149_0;    relay_conn far_4_4149_0_a(.in(layer_3[331]), .out(far_4_4149_0[0]));    relay_conn far_4_4149_0_b(.in(layer_3[418]), .out(far_4_4149_0[1]));
    wire [1:0] far_4_4149_1;    relay_conn far_4_4149_1_a(.in(far_4_4149_0[0]), .out(far_4_4149_1[0]));    relay_conn far_4_4149_1_b(.in(far_4_4149_0[1]), .out(far_4_4149_1[1]));
    assign layer_4[69] = far_4_4149_1[0] & far_4_4149_1[1]; 
    wire [1:0] far_4_4150_0;    relay_conn far_4_4150_0_a(.in(layer_3[620]), .out(far_4_4150_0[0]));    relay_conn far_4_4150_0_b(.in(layer_3[681]), .out(far_4_4150_0[1]));
    assign layer_4[70] = far_4_4150_0[1] & ~far_4_4150_0[0]; 
    wire [1:0] far_4_4151_0;    relay_conn far_4_4151_0_a(.in(layer_3[648]), .out(far_4_4151_0[0]));    relay_conn far_4_4151_0_b(.in(layer_3[744]), .out(far_4_4151_0[1]));
    wire [1:0] far_4_4151_1;    relay_conn far_4_4151_1_a(.in(far_4_4151_0[0]), .out(far_4_4151_1[0]));    relay_conn far_4_4151_1_b(.in(far_4_4151_0[1]), .out(far_4_4151_1[1]));
    wire [1:0] far_4_4151_2;    relay_conn far_4_4151_2_a(.in(far_4_4151_1[0]), .out(far_4_4151_2[0]));    relay_conn far_4_4151_2_b(.in(far_4_4151_1[1]), .out(far_4_4151_2[1]));
    assign layer_4[71] = ~far_4_4151_2[0]; 
    wire [1:0] far_4_4152_0;    relay_conn far_4_4152_0_a(.in(layer_3[907]), .out(far_4_4152_0[0]));    relay_conn far_4_4152_0_b(.in(layer_3[952]), .out(far_4_4152_0[1]));
    assign layer_4[72] = ~far_4_4152_0[1] | (far_4_4152_0[0] & far_4_4152_0[1]); 
    wire [1:0] far_4_4153_0;    relay_conn far_4_4153_0_a(.in(layer_3[334]), .out(far_4_4153_0[0]));    relay_conn far_4_4153_0_b(.in(layer_3[434]), .out(far_4_4153_0[1]));
    wire [1:0] far_4_4153_1;    relay_conn far_4_4153_1_a(.in(far_4_4153_0[0]), .out(far_4_4153_1[0]));    relay_conn far_4_4153_1_b(.in(far_4_4153_0[1]), .out(far_4_4153_1[1]));
    wire [1:0] far_4_4153_2;    relay_conn far_4_4153_2_a(.in(far_4_4153_1[0]), .out(far_4_4153_2[0]));    relay_conn far_4_4153_2_b(.in(far_4_4153_1[1]), .out(far_4_4153_2[1]));
    assign layer_4[73] = ~far_4_4153_2[0] | (far_4_4153_2[0] & far_4_4153_2[1]); 
    wire [1:0] far_4_4154_0;    relay_conn far_4_4154_0_a(.in(layer_3[879]), .out(far_4_4154_0[0]));    relay_conn far_4_4154_0_b(.in(layer_3[1004]), .out(far_4_4154_0[1]));
    wire [1:0] far_4_4154_1;    relay_conn far_4_4154_1_a(.in(far_4_4154_0[0]), .out(far_4_4154_1[0]));    relay_conn far_4_4154_1_b(.in(far_4_4154_0[1]), .out(far_4_4154_1[1]));
    wire [1:0] far_4_4154_2;    relay_conn far_4_4154_2_a(.in(far_4_4154_1[0]), .out(far_4_4154_2[0]));    relay_conn far_4_4154_2_b(.in(far_4_4154_1[1]), .out(far_4_4154_2[1]));
    assign layer_4[74] = far_4_4154_2[1]; 
    wire [1:0] far_4_4155_0;    relay_conn far_4_4155_0_a(.in(layer_3[838]), .out(far_4_4155_0[0]));    relay_conn far_4_4155_0_b(.in(layer_3[923]), .out(far_4_4155_0[1]));
    wire [1:0] far_4_4155_1;    relay_conn far_4_4155_1_a(.in(far_4_4155_0[0]), .out(far_4_4155_1[0]));    relay_conn far_4_4155_1_b(.in(far_4_4155_0[1]), .out(far_4_4155_1[1]));
    assign layer_4[75] = far_4_4155_1[0] | far_4_4155_1[1]; 
    wire [1:0] far_4_4156_0;    relay_conn far_4_4156_0_a(.in(layer_3[190]), .out(far_4_4156_0[0]));    relay_conn far_4_4156_0_b(.in(layer_3[97]), .out(far_4_4156_0[1]));
    wire [1:0] far_4_4156_1;    relay_conn far_4_4156_1_a(.in(far_4_4156_0[0]), .out(far_4_4156_1[0]));    relay_conn far_4_4156_1_b(.in(far_4_4156_0[1]), .out(far_4_4156_1[1]));
    assign layer_4[76] = ~far_4_4156_1[0]; 
    wire [1:0] far_4_4157_0;    relay_conn far_4_4157_0_a(.in(layer_3[277]), .out(far_4_4157_0[0]));    relay_conn far_4_4157_0_b(.in(layer_3[236]), .out(far_4_4157_0[1]));
    assign layer_4[77] = ~far_4_4157_0[1]; 
    wire [1:0] far_4_4158_0;    relay_conn far_4_4158_0_a(.in(layer_3[334]), .out(far_4_4158_0[0]));    relay_conn far_4_4158_0_b(.in(layer_3[440]), .out(far_4_4158_0[1]));
    wire [1:0] far_4_4158_1;    relay_conn far_4_4158_1_a(.in(far_4_4158_0[0]), .out(far_4_4158_1[0]));    relay_conn far_4_4158_1_b(.in(far_4_4158_0[1]), .out(far_4_4158_1[1]));
    wire [1:0] far_4_4158_2;    relay_conn far_4_4158_2_a(.in(far_4_4158_1[0]), .out(far_4_4158_2[0]));    relay_conn far_4_4158_2_b(.in(far_4_4158_1[1]), .out(far_4_4158_2[1]));
    assign layer_4[78] = far_4_4158_2[0]; 
    wire [1:0] far_4_4159_0;    relay_conn far_4_4159_0_a(.in(layer_3[192]), .out(far_4_4159_0[0]));    relay_conn far_4_4159_0_b(.in(layer_3[129]), .out(far_4_4159_0[1]));
    assign layer_4[79] = ~(far_4_4159_0[0] & far_4_4159_0[1]); 
    wire [1:0] far_4_4160_0;    relay_conn far_4_4160_0_a(.in(layer_3[716]), .out(far_4_4160_0[0]));    relay_conn far_4_4160_0_b(.in(layer_3[661]), .out(far_4_4160_0[1]));
    assign layer_4[80] = ~far_4_4160_0[1] | (far_4_4160_0[0] & far_4_4160_0[1]); 
    wire [1:0] far_4_4161_0;    relay_conn far_4_4161_0_a(.in(layer_3[811]), .out(far_4_4161_0[0]));    relay_conn far_4_4161_0_b(.in(layer_3[910]), .out(far_4_4161_0[1]));
    wire [1:0] far_4_4161_1;    relay_conn far_4_4161_1_a(.in(far_4_4161_0[0]), .out(far_4_4161_1[0]));    relay_conn far_4_4161_1_b(.in(far_4_4161_0[1]), .out(far_4_4161_1[1]));
    wire [1:0] far_4_4161_2;    relay_conn far_4_4161_2_a(.in(far_4_4161_1[0]), .out(far_4_4161_2[0]));    relay_conn far_4_4161_2_b(.in(far_4_4161_1[1]), .out(far_4_4161_2[1]));
    assign layer_4[81] = ~far_4_4161_2[0] | (far_4_4161_2[0] & far_4_4161_2[1]); 
    assign layer_4[82] = ~layer_3[56] | (layer_3[56] & layer_3[35]); 
    wire [1:0] far_4_4163_0;    relay_conn far_4_4163_0_a(.in(layer_3[778]), .out(far_4_4163_0[0]));    relay_conn far_4_4163_0_b(.in(layer_3[818]), .out(far_4_4163_0[1]));
    assign layer_4[83] = ~(far_4_4163_0[0] ^ far_4_4163_0[1]); 
    wire [1:0] far_4_4164_0;    relay_conn far_4_4164_0_a(.in(layer_3[630]), .out(far_4_4164_0[0]));    relay_conn far_4_4164_0_b(.in(layer_3[577]), .out(far_4_4164_0[1]));
    assign layer_4[84] = far_4_4164_0[0]; 
    assign layer_4[85] = layer_3[577]; 
    wire [1:0] far_4_4166_0;    relay_conn far_4_4166_0_a(.in(layer_3[633]), .out(far_4_4166_0[0]));    relay_conn far_4_4166_0_b(.in(layer_3[716]), .out(far_4_4166_0[1]));
    wire [1:0] far_4_4166_1;    relay_conn far_4_4166_1_a(.in(far_4_4166_0[0]), .out(far_4_4166_1[0]));    relay_conn far_4_4166_1_b(.in(far_4_4166_0[1]), .out(far_4_4166_1[1]));
    assign layer_4[86] = ~(far_4_4166_1[0] | far_4_4166_1[1]); 
    wire [1:0] far_4_4167_0;    relay_conn far_4_4167_0_a(.in(layer_3[36]), .out(far_4_4167_0[0]));    relay_conn far_4_4167_0_b(.in(layer_3[94]), .out(far_4_4167_0[1]));
    assign layer_4[87] = ~(far_4_4167_0[0] ^ far_4_4167_0[1]); 
    assign layer_4[88] = ~layer_3[630]; 
    wire [1:0] far_4_4169_0;    relay_conn far_4_4169_0_a(.in(layer_3[807]), .out(far_4_4169_0[0]));    relay_conn far_4_4169_0_b(.in(layer_3[879]), .out(far_4_4169_0[1]));
    wire [1:0] far_4_4169_1;    relay_conn far_4_4169_1_a(.in(far_4_4169_0[0]), .out(far_4_4169_1[0]));    relay_conn far_4_4169_1_b(.in(far_4_4169_0[1]), .out(far_4_4169_1[1]));
    assign layer_4[89] = far_4_4169_1[0] & far_4_4169_1[1]; 
    wire [1:0] far_4_4170_0;    relay_conn far_4_4170_0_a(.in(layer_3[823]), .out(far_4_4170_0[0]));    relay_conn far_4_4170_0_b(.in(layer_3[770]), .out(far_4_4170_0[1]));
    assign layer_4[90] = far_4_4170_0[0] & far_4_4170_0[1]; 
    wire [1:0] far_4_4171_0;    relay_conn far_4_4171_0_a(.in(layer_3[756]), .out(far_4_4171_0[0]));    relay_conn far_4_4171_0_b(.in(layer_3[662]), .out(far_4_4171_0[1]));
    wire [1:0] far_4_4171_1;    relay_conn far_4_4171_1_a(.in(far_4_4171_0[0]), .out(far_4_4171_1[0]));    relay_conn far_4_4171_1_b(.in(far_4_4171_0[1]), .out(far_4_4171_1[1]));
    assign layer_4[91] = ~far_4_4171_1[0] | (far_4_4171_1[0] & far_4_4171_1[1]); 
    wire [1:0] far_4_4172_0;    relay_conn far_4_4172_0_a(.in(layer_3[365]), .out(far_4_4172_0[0]));    relay_conn far_4_4172_0_b(.in(layer_3[242]), .out(far_4_4172_0[1]));
    wire [1:0] far_4_4172_1;    relay_conn far_4_4172_1_a(.in(far_4_4172_0[0]), .out(far_4_4172_1[0]));    relay_conn far_4_4172_1_b(.in(far_4_4172_0[1]), .out(far_4_4172_1[1]));
    wire [1:0] far_4_4172_2;    relay_conn far_4_4172_2_a(.in(far_4_4172_1[0]), .out(far_4_4172_2[0]));    relay_conn far_4_4172_2_b(.in(far_4_4172_1[1]), .out(far_4_4172_2[1]));
    assign layer_4[92] = ~far_4_4172_2[1] | (far_4_4172_2[0] & far_4_4172_2[1]); 
    wire [1:0] far_4_4173_0;    relay_conn far_4_4173_0_a(.in(layer_3[80]), .out(far_4_4173_0[0]));    relay_conn far_4_4173_0_b(.in(layer_3[136]), .out(far_4_4173_0[1]));
    assign layer_4[93] = ~(far_4_4173_0[0] & far_4_4173_0[1]); 
    wire [1:0] far_4_4174_0;    relay_conn far_4_4174_0_a(.in(layer_3[264]), .out(far_4_4174_0[0]));    relay_conn far_4_4174_0_b(.in(layer_3[184]), .out(far_4_4174_0[1]));
    wire [1:0] far_4_4174_1;    relay_conn far_4_4174_1_a(.in(far_4_4174_0[0]), .out(far_4_4174_1[0]));    relay_conn far_4_4174_1_b(.in(far_4_4174_0[1]), .out(far_4_4174_1[1]));
    assign layer_4[94] = far_4_4174_1[0] | far_4_4174_1[1]; 
    wire [1:0] far_4_4175_0;    relay_conn far_4_4175_0_a(.in(layer_3[346]), .out(far_4_4175_0[0]));    relay_conn far_4_4175_0_b(.in(layer_3[420]), .out(far_4_4175_0[1]));
    wire [1:0] far_4_4175_1;    relay_conn far_4_4175_1_a(.in(far_4_4175_0[0]), .out(far_4_4175_1[0]));    relay_conn far_4_4175_1_b(.in(far_4_4175_0[1]), .out(far_4_4175_1[1]));
    assign layer_4[95] = ~(far_4_4175_1[0] | far_4_4175_1[1]); 
    wire [1:0] far_4_4176_0;    relay_conn far_4_4176_0_a(.in(layer_3[578]), .out(far_4_4176_0[0]));    relay_conn far_4_4176_0_b(.in(layer_3[629]), .out(far_4_4176_0[1]));
    assign layer_4[96] = far_4_4176_0[0] & far_4_4176_0[1]; 
    wire [1:0] far_4_4177_0;    relay_conn far_4_4177_0_a(.in(layer_3[842]), .out(far_4_4177_0[0]));    relay_conn far_4_4177_0_b(.in(layer_3[921]), .out(far_4_4177_0[1]));
    wire [1:0] far_4_4177_1;    relay_conn far_4_4177_1_a(.in(far_4_4177_0[0]), .out(far_4_4177_1[0]));    relay_conn far_4_4177_1_b(.in(far_4_4177_0[1]), .out(far_4_4177_1[1]));
    assign layer_4[97] = ~far_4_4177_1[1] | (far_4_4177_1[0] & far_4_4177_1[1]); 
    wire [1:0] far_4_4178_0;    relay_conn far_4_4178_0_a(.in(layer_3[993]), .out(far_4_4178_0[0]));    relay_conn far_4_4178_0_b(.in(layer_3[924]), .out(far_4_4178_0[1]));
    wire [1:0] far_4_4178_1;    relay_conn far_4_4178_1_a(.in(far_4_4178_0[0]), .out(far_4_4178_1[0]));    relay_conn far_4_4178_1_b(.in(far_4_4178_0[1]), .out(far_4_4178_1[1]));
    assign layer_4[98] = ~far_4_4178_1[1] | (far_4_4178_1[0] & far_4_4178_1[1]); 
    wire [1:0] far_4_4179_0;    relay_conn far_4_4179_0_a(.in(layer_3[468]), .out(far_4_4179_0[0]));    relay_conn far_4_4179_0_b(.in(layer_3[578]), .out(far_4_4179_0[1]));
    wire [1:0] far_4_4179_1;    relay_conn far_4_4179_1_a(.in(far_4_4179_0[0]), .out(far_4_4179_1[0]));    relay_conn far_4_4179_1_b(.in(far_4_4179_0[1]), .out(far_4_4179_1[1]));
    wire [1:0] far_4_4179_2;    relay_conn far_4_4179_2_a(.in(far_4_4179_1[0]), .out(far_4_4179_2[0]));    relay_conn far_4_4179_2_b(.in(far_4_4179_1[1]), .out(far_4_4179_2[1]));
    assign layer_4[99] = far_4_4179_2[0] | far_4_4179_2[1]; 
    wire [1:0] far_4_4180_0;    relay_conn far_4_4180_0_a(.in(layer_3[433]), .out(far_4_4180_0[0]));    relay_conn far_4_4180_0_b(.in(layer_3[397]), .out(far_4_4180_0[1]));
    assign layer_4[100] = far_4_4180_0[0] | far_4_4180_0[1]; 
    wire [1:0] far_4_4181_0;    relay_conn far_4_4181_0_a(.in(layer_3[830]), .out(far_4_4181_0[0]));    relay_conn far_4_4181_0_b(.in(layer_3[775]), .out(far_4_4181_0[1]));
    assign layer_4[101] = ~(far_4_4181_0[0] ^ far_4_4181_0[1]); 
    wire [1:0] far_4_4182_0;    relay_conn far_4_4182_0_a(.in(layer_3[467]), .out(far_4_4182_0[0]));    relay_conn far_4_4182_0_b(.in(layer_3[576]), .out(far_4_4182_0[1]));
    wire [1:0] far_4_4182_1;    relay_conn far_4_4182_1_a(.in(far_4_4182_0[0]), .out(far_4_4182_1[0]));    relay_conn far_4_4182_1_b(.in(far_4_4182_0[1]), .out(far_4_4182_1[1]));
    wire [1:0] far_4_4182_2;    relay_conn far_4_4182_2_a(.in(far_4_4182_1[0]), .out(far_4_4182_2[0]));    relay_conn far_4_4182_2_b(.in(far_4_4182_1[1]), .out(far_4_4182_2[1]));
    assign layer_4[102] = far_4_4182_2[0] | far_4_4182_2[1]; 
    wire [1:0] far_4_4183_0;    relay_conn far_4_4183_0_a(.in(layer_3[576]), .out(far_4_4183_0[0]));    relay_conn far_4_4183_0_b(.in(layer_3[525]), .out(far_4_4183_0[1]));
    assign layer_4[103] = far_4_4183_0[0] & ~far_4_4183_0[1]; 
    wire [1:0] far_4_4184_0;    relay_conn far_4_4184_0_a(.in(layer_3[635]), .out(far_4_4184_0[0]));    relay_conn far_4_4184_0_b(.in(layer_3[576]), .out(far_4_4184_0[1]));
    assign layer_4[104] = ~(far_4_4184_0[0] | far_4_4184_0[1]); 
    assign layer_4[105] = layer_3[749] & ~layer_3[735]; 
    wire [1:0] far_4_4186_0;    relay_conn far_4_4186_0_a(.in(layer_3[302]), .out(far_4_4186_0[0]));    relay_conn far_4_4186_0_b(.in(layer_3[255]), .out(far_4_4186_0[1]));
    assign layer_4[106] = ~(far_4_4186_0[0] | far_4_4186_0[1]); 
    assign layer_4[107] = ~(layer_3[466] & layer_3[438]); 
    assign layer_4[108] = ~layer_3[32] | (layer_3[32] & layer_3[43]); 
    assign layer_4[109] = ~layer_3[660] | (layer_3[660] & layer_3[666]); 
    wire [1:0] far_4_4190_0;    relay_conn far_4_4190_0_a(.in(layer_3[838]), .out(far_4_4190_0[0]));    relay_conn far_4_4190_0_b(.in(layer_3[770]), .out(far_4_4190_0[1]));
    wire [1:0] far_4_4190_1;    relay_conn far_4_4190_1_a(.in(far_4_4190_0[0]), .out(far_4_4190_1[0]));    relay_conn far_4_4190_1_b(.in(far_4_4190_0[1]), .out(far_4_4190_1[1]));
    assign layer_4[110] = ~far_4_4190_1[0]; 
    wire [1:0] far_4_4191_0;    relay_conn far_4_4191_0_a(.in(layer_3[880]), .out(far_4_4191_0[0]));    relay_conn far_4_4191_0_b(.in(layer_3[834]), .out(far_4_4191_0[1]));
    assign layer_4[111] = far_4_4191_0[1]; 
    wire [1:0] far_4_4192_0;    relay_conn far_4_4192_0_a(.in(layer_3[497]), .out(far_4_4192_0[0]));    relay_conn far_4_4192_0_b(.in(layer_3[411]), .out(far_4_4192_0[1]));
    wire [1:0] far_4_4192_1;    relay_conn far_4_4192_1_a(.in(far_4_4192_0[0]), .out(far_4_4192_1[0]));    relay_conn far_4_4192_1_b(.in(far_4_4192_0[1]), .out(far_4_4192_1[1]));
    assign layer_4[112] = ~(far_4_4192_1[0] ^ far_4_4192_1[1]); 
    wire [1:0] far_4_4193_0;    relay_conn far_4_4193_0_a(.in(layer_3[935]), .out(far_4_4193_0[0]));    relay_conn far_4_4193_0_b(.in(layer_3[979]), .out(far_4_4193_0[1]));
    assign layer_4[113] = far_4_4193_0[0]; 
    wire [1:0] far_4_4194_0;    relay_conn far_4_4194_0_a(.in(layer_3[455]), .out(far_4_4194_0[0]));    relay_conn far_4_4194_0_b(.in(layer_3[507]), .out(far_4_4194_0[1]));
    assign layer_4[114] = ~far_4_4194_0[1]; 
    assign layer_4[115] = ~layer_3[952]; 
    wire [1:0] far_4_4196_0;    relay_conn far_4_4196_0_a(.in(layer_3[626]), .out(far_4_4196_0[0]));    relay_conn far_4_4196_0_b(.in(layer_3[659]), .out(far_4_4196_0[1]));
    assign layer_4[116] = far_4_4196_0[0] ^ far_4_4196_0[1]; 
    wire [1:0] far_4_4197_0;    relay_conn far_4_4197_0_a(.in(layer_3[823]), .out(far_4_4197_0[0]));    relay_conn far_4_4197_0_b(.in(layer_3[900]), .out(far_4_4197_0[1]));
    wire [1:0] far_4_4197_1;    relay_conn far_4_4197_1_a(.in(far_4_4197_0[0]), .out(far_4_4197_1[0]));    relay_conn far_4_4197_1_b(.in(far_4_4197_0[1]), .out(far_4_4197_1[1]));
    assign layer_4[117] = far_4_4197_1[1] & ~far_4_4197_1[0]; 
    wire [1:0] far_4_4198_0;    relay_conn far_4_4198_0_a(.in(layer_3[782]), .out(far_4_4198_0[0]));    relay_conn far_4_4198_0_b(.in(layer_3[901]), .out(far_4_4198_0[1]));
    wire [1:0] far_4_4198_1;    relay_conn far_4_4198_1_a(.in(far_4_4198_0[0]), .out(far_4_4198_1[0]));    relay_conn far_4_4198_1_b(.in(far_4_4198_0[1]), .out(far_4_4198_1[1]));
    wire [1:0] far_4_4198_2;    relay_conn far_4_4198_2_a(.in(far_4_4198_1[0]), .out(far_4_4198_2[0]));    relay_conn far_4_4198_2_b(.in(far_4_4198_1[1]), .out(far_4_4198_2[1]));
    assign layer_4[118] = far_4_4198_2[0] | far_4_4198_2[1]; 
    wire [1:0] far_4_4199_0;    relay_conn far_4_4199_0_a(.in(layer_3[549]), .out(far_4_4199_0[0]));    relay_conn far_4_4199_0_b(.in(layer_3[487]), .out(far_4_4199_0[1]));
    assign layer_4[119] = ~(far_4_4199_0[0] | far_4_4199_0[1]); 
    wire [1:0] far_4_4200_0;    relay_conn far_4_4200_0_a(.in(layer_3[834]), .out(far_4_4200_0[0]));    relay_conn far_4_4200_0_b(.in(layer_3[746]), .out(far_4_4200_0[1]));
    wire [1:0] far_4_4200_1;    relay_conn far_4_4200_1_a(.in(far_4_4200_0[0]), .out(far_4_4200_1[0]));    relay_conn far_4_4200_1_b(.in(far_4_4200_0[1]), .out(far_4_4200_1[1]));
    assign layer_4[120] = ~far_4_4200_1[0]; 
    wire [1:0] far_4_4201_0;    relay_conn far_4_4201_0_a(.in(layer_3[914]), .out(far_4_4201_0[0]));    relay_conn far_4_4201_0_b(.in(layer_3[868]), .out(far_4_4201_0[1]));
    assign layer_4[121] = ~far_4_4201_0[0]; 
    wire [1:0] far_4_4202_0;    relay_conn far_4_4202_0_a(.in(layer_3[589]), .out(far_4_4202_0[0]));    relay_conn far_4_4202_0_b(.in(layer_3[644]), .out(far_4_4202_0[1]));
    assign layer_4[122] = far_4_4202_0[1]; 
    assign layer_4[123] = layer_3[953] & ~layer_3[979]; 
    wire [1:0] far_4_4204_0;    relay_conn far_4_4204_0_a(.in(layer_3[793]), .out(far_4_4204_0[0]));    relay_conn far_4_4204_0_b(.in(layer_3[748]), .out(far_4_4204_0[1]));
    assign layer_4[124] = far_4_4204_0[0] & far_4_4204_0[1]; 
    assign layer_4[125] = ~layer_3[628]; 
    wire [1:0] far_4_4206_0;    relay_conn far_4_4206_0_a(.in(layer_3[332]), .out(far_4_4206_0[0]));    relay_conn far_4_4206_0_b(.in(layer_3[234]), .out(far_4_4206_0[1]));
    wire [1:0] far_4_4206_1;    relay_conn far_4_4206_1_a(.in(far_4_4206_0[0]), .out(far_4_4206_1[0]));    relay_conn far_4_4206_1_b(.in(far_4_4206_0[1]), .out(far_4_4206_1[1]));
    wire [1:0] far_4_4206_2;    relay_conn far_4_4206_2_a(.in(far_4_4206_1[0]), .out(far_4_4206_2[0]));    relay_conn far_4_4206_2_b(.in(far_4_4206_1[1]), .out(far_4_4206_2[1]));
    assign layer_4[126] = ~far_4_4206_2[1]; 
    wire [1:0] far_4_4207_0;    relay_conn far_4_4207_0_a(.in(layer_3[605]), .out(far_4_4207_0[0]));    relay_conn far_4_4207_0_b(.in(layer_3[705]), .out(far_4_4207_0[1]));
    wire [1:0] far_4_4207_1;    relay_conn far_4_4207_1_a(.in(far_4_4207_0[0]), .out(far_4_4207_1[0]));    relay_conn far_4_4207_1_b(.in(far_4_4207_0[1]), .out(far_4_4207_1[1]));
    wire [1:0] far_4_4207_2;    relay_conn far_4_4207_2_a(.in(far_4_4207_1[0]), .out(far_4_4207_2[0]));    relay_conn far_4_4207_2_b(.in(far_4_4207_1[1]), .out(far_4_4207_2[1]));
    assign layer_4[127] = ~far_4_4207_2[0]; 
    wire [1:0] far_4_4208_0;    relay_conn far_4_4208_0_a(.in(layer_3[708]), .out(far_4_4208_0[0]));    relay_conn far_4_4208_0_b(.in(layer_3[778]), .out(far_4_4208_0[1]));
    wire [1:0] far_4_4208_1;    relay_conn far_4_4208_1_a(.in(far_4_4208_0[0]), .out(far_4_4208_1[0]));    relay_conn far_4_4208_1_b(.in(far_4_4208_0[1]), .out(far_4_4208_1[1]));
    assign layer_4[128] = ~far_4_4208_1[0] | (far_4_4208_1[0] & far_4_4208_1[1]); 
    wire [1:0] far_4_4209_0;    relay_conn far_4_4209_0_a(.in(layer_3[696]), .out(far_4_4209_0[0]));    relay_conn far_4_4209_0_b(.in(layer_3[661]), .out(far_4_4209_0[1]));
    assign layer_4[129] = ~far_4_4209_0[0]; 
    wire [1:0] far_4_4210_0;    relay_conn far_4_4210_0_a(.in(layer_3[730]), .out(far_4_4210_0[0]));    relay_conn far_4_4210_0_b(.in(layer_3[634]), .out(far_4_4210_0[1]));
    wire [1:0] far_4_4210_1;    relay_conn far_4_4210_1_a(.in(far_4_4210_0[0]), .out(far_4_4210_1[0]));    relay_conn far_4_4210_1_b(.in(far_4_4210_0[1]), .out(far_4_4210_1[1]));
    wire [1:0] far_4_4210_2;    relay_conn far_4_4210_2_a(.in(far_4_4210_1[0]), .out(far_4_4210_2[0]));    relay_conn far_4_4210_2_b(.in(far_4_4210_1[1]), .out(far_4_4210_2[1]));
    assign layer_4[130] = ~far_4_4210_2[0]; 
    wire [1:0] far_4_4211_0;    relay_conn far_4_4211_0_a(.in(layer_3[466]), .out(far_4_4211_0[0]));    relay_conn far_4_4211_0_b(.in(layer_3[576]), .out(far_4_4211_0[1]));
    wire [1:0] far_4_4211_1;    relay_conn far_4_4211_1_a(.in(far_4_4211_0[0]), .out(far_4_4211_1[0]));    relay_conn far_4_4211_1_b(.in(far_4_4211_0[1]), .out(far_4_4211_1[1]));
    wire [1:0] far_4_4211_2;    relay_conn far_4_4211_2_a(.in(far_4_4211_1[0]), .out(far_4_4211_2[0]));    relay_conn far_4_4211_2_b(.in(far_4_4211_1[1]), .out(far_4_4211_2[1]));
    assign layer_4[131] = ~far_4_4211_2[0] | (far_4_4211_2[0] & far_4_4211_2[1]); 
    assign layer_4[132] = layer_3[605] | layer_3[608]; 
    wire [1:0] far_4_4213_0;    relay_conn far_4_4213_0_a(.in(layer_3[45]), .out(far_4_4213_0[0]));    relay_conn far_4_4213_0_b(.in(layer_3[113]), .out(far_4_4213_0[1]));
    wire [1:0] far_4_4213_1;    relay_conn far_4_4213_1_a(.in(far_4_4213_0[0]), .out(far_4_4213_1[0]));    relay_conn far_4_4213_1_b(.in(far_4_4213_0[1]), .out(far_4_4213_1[1]));
    assign layer_4[133] = far_4_4213_1[1] & ~far_4_4213_1[0]; 
    wire [1:0] far_4_4214_0;    relay_conn far_4_4214_0_a(.in(layer_3[900]), .out(far_4_4214_0[0]));    relay_conn far_4_4214_0_b(.in(layer_3[780]), .out(far_4_4214_0[1]));
    wire [1:0] far_4_4214_1;    relay_conn far_4_4214_1_a(.in(far_4_4214_0[0]), .out(far_4_4214_1[0]));    relay_conn far_4_4214_1_b(.in(far_4_4214_0[1]), .out(far_4_4214_1[1]));
    wire [1:0] far_4_4214_2;    relay_conn far_4_4214_2_a(.in(far_4_4214_1[0]), .out(far_4_4214_2[0]));    relay_conn far_4_4214_2_b(.in(far_4_4214_1[1]), .out(far_4_4214_2[1]));
    assign layer_4[134] = far_4_4214_2[1] & ~far_4_4214_2[0]; 
    wire [1:0] far_4_4215_0;    relay_conn far_4_4215_0_a(.in(layer_3[835]), .out(far_4_4215_0[0]));    relay_conn far_4_4215_0_b(.in(layer_3[777]), .out(far_4_4215_0[1]));
    assign layer_4[135] = ~(far_4_4215_0[0] & far_4_4215_0[1]); 
    assign layer_4[136] = ~(layer_3[507] & layer_3[486]); 
    wire [1:0] far_4_4217_0;    relay_conn far_4_4217_0_a(.in(layer_3[610]), .out(far_4_4217_0[0]));    relay_conn far_4_4217_0_b(.in(layer_3[686]), .out(far_4_4217_0[1]));
    wire [1:0] far_4_4217_1;    relay_conn far_4_4217_1_a(.in(far_4_4217_0[0]), .out(far_4_4217_1[0]));    relay_conn far_4_4217_1_b(.in(far_4_4217_0[1]), .out(far_4_4217_1[1]));
    assign layer_4[137] = far_4_4217_1[1]; 
    wire [1:0] far_4_4218_0;    relay_conn far_4_4218_0_a(.in(layer_3[898]), .out(far_4_4218_0[0]));    relay_conn far_4_4218_0_b(.in(layer_3[770]), .out(far_4_4218_0[1]));
    wire [1:0] far_4_4218_1;    relay_conn far_4_4218_1_a(.in(far_4_4218_0[0]), .out(far_4_4218_1[0]));    relay_conn far_4_4218_1_b(.in(far_4_4218_0[1]), .out(far_4_4218_1[1]));
    wire [1:0] far_4_4218_2;    relay_conn far_4_4218_2_a(.in(far_4_4218_1[0]), .out(far_4_4218_2[0]));    relay_conn far_4_4218_2_b(.in(far_4_4218_1[1]), .out(far_4_4218_2[1]));
    wire [1:0] far_4_4218_3;    relay_conn far_4_4218_3_a(.in(far_4_4218_2[0]), .out(far_4_4218_3[0]));    relay_conn far_4_4218_3_b(.in(far_4_4218_2[1]), .out(far_4_4218_3[1]));
    assign layer_4[138] = far_4_4218_3[0] ^ far_4_4218_3[1]; 
    wire [1:0] far_4_4219_0;    relay_conn far_4_4219_0_a(.in(layer_3[56]), .out(far_4_4219_0[0]));    relay_conn far_4_4219_0_b(.in(layer_3[93]), .out(far_4_4219_0[1]));
    assign layer_4[139] = far_4_4219_0[0] & far_4_4219_0[1]; 
    wire [1:0] far_4_4220_0;    relay_conn far_4_4220_0_a(.in(layer_3[599]), .out(far_4_4220_0[0]));    relay_conn far_4_4220_0_b(.in(layer_3[556]), .out(far_4_4220_0[1]));
    assign layer_4[140] = ~far_4_4220_0[1]; 
    wire [1:0] far_4_4221_0;    relay_conn far_4_4221_0_a(.in(layer_3[610]), .out(far_4_4221_0[0]));    relay_conn far_4_4221_0_b(.in(layer_3[559]), .out(far_4_4221_0[1]));
    assign layer_4[141] = far_4_4221_0[1]; 
    wire [1:0] far_4_4222_0;    relay_conn far_4_4222_0_a(.in(layer_3[846]), .out(far_4_4222_0[0]));    relay_conn far_4_4222_0_b(.in(layer_3[905]), .out(far_4_4222_0[1]));
    assign layer_4[142] = ~(far_4_4222_0[0] | far_4_4222_0[1]); 
    assign layer_4[143] = layer_3[972] & ~layer_3[979]; 
    assign layer_4[144] = layer_3[423] ^ layer_3[431]; 
    wire [1:0] far_4_4225_0;    relay_conn far_4_4225_0_a(.in(layer_3[114]), .out(far_4_4225_0[0]));    relay_conn far_4_4225_0_b(.in(layer_3[152]), .out(far_4_4225_0[1]));
    assign layer_4[145] = ~(far_4_4225_0[0] & far_4_4225_0[1]); 
    wire [1:0] far_4_4226_0;    relay_conn far_4_4226_0_a(.in(layer_3[332]), .out(far_4_4226_0[0]));    relay_conn far_4_4226_0_b(.in(layer_3[391]), .out(far_4_4226_0[1]));
    assign layer_4[146] = ~far_4_4226_0[1]; 
    wire [1:0] far_4_4227_0;    relay_conn far_4_4227_0_a(.in(layer_3[429]), .out(far_4_4227_0[0]));    relay_conn far_4_4227_0_b(.in(layer_3[511]), .out(far_4_4227_0[1]));
    wire [1:0] far_4_4227_1;    relay_conn far_4_4227_1_a(.in(far_4_4227_0[0]), .out(far_4_4227_1[0]));    relay_conn far_4_4227_1_b(.in(far_4_4227_0[1]), .out(far_4_4227_1[1]));
    assign layer_4[147] = far_4_4227_1[1] & ~far_4_4227_1[0]; 
    wire [1:0] far_4_4228_0;    relay_conn far_4_4228_0_a(.in(layer_3[807]), .out(far_4_4228_0[0]));    relay_conn far_4_4228_0_b(.in(layer_3[880]), .out(far_4_4228_0[1]));
    wire [1:0] far_4_4228_1;    relay_conn far_4_4228_1_a(.in(far_4_4228_0[0]), .out(far_4_4228_1[0]));    relay_conn far_4_4228_1_b(.in(far_4_4228_0[1]), .out(far_4_4228_1[1]));
    assign layer_4[148] = ~(far_4_4228_1[0] & far_4_4228_1[1]); 
    assign layer_4[149] = layer_3[27] & ~layer_3[41]; 
    wire [1:0] far_4_4230_0;    relay_conn far_4_4230_0_a(.in(layer_3[400]), .out(far_4_4230_0[0]));    relay_conn far_4_4230_0_b(.in(layer_3[337]), .out(far_4_4230_0[1]));
    assign layer_4[150] = ~far_4_4230_0[1]; 
    wire [1:0] far_4_4231_0;    relay_conn far_4_4231_0_a(.in(layer_3[577]), .out(far_4_4231_0[0]));    relay_conn far_4_4231_0_b(.in(layer_3[479]), .out(far_4_4231_0[1]));
    wire [1:0] far_4_4231_1;    relay_conn far_4_4231_1_a(.in(far_4_4231_0[0]), .out(far_4_4231_1[0]));    relay_conn far_4_4231_1_b(.in(far_4_4231_0[1]), .out(far_4_4231_1[1]));
    wire [1:0] far_4_4231_2;    relay_conn far_4_4231_2_a(.in(far_4_4231_1[0]), .out(far_4_4231_2[0]));    relay_conn far_4_4231_2_b(.in(far_4_4231_1[1]), .out(far_4_4231_2[1]));
    assign layer_4[151] = far_4_4231_2[0]; 
    wire [1:0] far_4_4232_0;    relay_conn far_4_4232_0_a(.in(layer_3[751]), .out(far_4_4232_0[0]));    relay_conn far_4_4232_0_b(.in(layer_3[653]), .out(far_4_4232_0[1]));
    wire [1:0] far_4_4232_1;    relay_conn far_4_4232_1_a(.in(far_4_4232_0[0]), .out(far_4_4232_1[0]));    relay_conn far_4_4232_1_b(.in(far_4_4232_0[1]), .out(far_4_4232_1[1]));
    wire [1:0] far_4_4232_2;    relay_conn far_4_4232_2_a(.in(far_4_4232_1[0]), .out(far_4_4232_2[0]));    relay_conn far_4_4232_2_b(.in(far_4_4232_1[1]), .out(far_4_4232_2[1]));
    assign layer_4[152] = ~far_4_4232_2[0] | (far_4_4232_2[0] & far_4_4232_2[1]); 
    wire [1:0] far_4_4233_0;    relay_conn far_4_4233_0_a(.in(layer_3[456]), .out(far_4_4233_0[0]));    relay_conn far_4_4233_0_b(.in(layer_3[351]), .out(far_4_4233_0[1]));
    wire [1:0] far_4_4233_1;    relay_conn far_4_4233_1_a(.in(far_4_4233_0[0]), .out(far_4_4233_1[0]));    relay_conn far_4_4233_1_b(.in(far_4_4233_0[1]), .out(far_4_4233_1[1]));
    wire [1:0] far_4_4233_2;    relay_conn far_4_4233_2_a(.in(far_4_4233_1[0]), .out(far_4_4233_2[0]));    relay_conn far_4_4233_2_b(.in(far_4_4233_1[1]), .out(far_4_4233_2[1]));
    assign layer_4[153] = ~far_4_4233_2[1]; 
    wire [1:0] far_4_4234_0;    relay_conn far_4_4234_0_a(.in(layer_3[257]), .out(far_4_4234_0[0]));    relay_conn far_4_4234_0_b(.in(layer_3[150]), .out(far_4_4234_0[1]));
    wire [1:0] far_4_4234_1;    relay_conn far_4_4234_1_a(.in(far_4_4234_0[0]), .out(far_4_4234_1[0]));    relay_conn far_4_4234_1_b(.in(far_4_4234_0[1]), .out(far_4_4234_1[1]));
    wire [1:0] far_4_4234_2;    relay_conn far_4_4234_2_a(.in(far_4_4234_1[0]), .out(far_4_4234_2[0]));    relay_conn far_4_4234_2_b(.in(far_4_4234_1[1]), .out(far_4_4234_2[1]));
    assign layer_4[154] = far_4_4234_2[1]; 
    assign layer_4[155] = ~layer_3[164] | (layer_3[165] & layer_3[164]); 
    assign layer_4[156] = ~layer_3[57] | (layer_3[57] & layer_3[72]); 
    wire [1:0] far_4_4237_0;    relay_conn far_4_4237_0_a(.in(layer_3[878]), .out(far_4_4237_0[0]));    relay_conn far_4_4237_0_b(.in(layer_3[834]), .out(far_4_4237_0[1]));
    assign layer_4[157] = far_4_4237_0[0] & far_4_4237_0[1]; 
    wire [1:0] far_4_4238_0;    relay_conn far_4_4238_0_a(.in(layer_3[576]), .out(far_4_4238_0[0]));    relay_conn far_4_4238_0_b(.in(layer_3[481]), .out(far_4_4238_0[1]));
    wire [1:0] far_4_4238_1;    relay_conn far_4_4238_1_a(.in(far_4_4238_0[0]), .out(far_4_4238_1[0]));    relay_conn far_4_4238_1_b(.in(far_4_4238_0[1]), .out(far_4_4238_1[1]));
    assign layer_4[158] = far_4_4238_1[0] & ~far_4_4238_1[1]; 
    wire [1:0] far_4_4239_0;    relay_conn far_4_4239_0_a(.in(layer_3[936]), .out(far_4_4239_0[0]));    relay_conn far_4_4239_0_b(.in(layer_3[831]), .out(far_4_4239_0[1]));
    wire [1:0] far_4_4239_1;    relay_conn far_4_4239_1_a(.in(far_4_4239_0[0]), .out(far_4_4239_1[0]));    relay_conn far_4_4239_1_b(.in(far_4_4239_0[1]), .out(far_4_4239_1[1]));
    wire [1:0] far_4_4239_2;    relay_conn far_4_4239_2_a(.in(far_4_4239_1[0]), .out(far_4_4239_2[0]));    relay_conn far_4_4239_2_b(.in(far_4_4239_1[1]), .out(far_4_4239_2[1]));
    assign layer_4[159] = far_4_4239_2[1]; 
    assign layer_4[160] = layer_3[807] & ~layer_3[779]; 
    wire [1:0] far_4_4241_0;    relay_conn far_4_4241_0_a(.in(layer_3[37]), .out(far_4_4241_0[0]));    relay_conn far_4_4241_0_b(.in(layer_3[135]), .out(far_4_4241_0[1]));
    wire [1:0] far_4_4241_1;    relay_conn far_4_4241_1_a(.in(far_4_4241_0[0]), .out(far_4_4241_1[0]));    relay_conn far_4_4241_1_b(.in(far_4_4241_0[1]), .out(far_4_4241_1[1]));
    wire [1:0] far_4_4241_2;    relay_conn far_4_4241_2_a(.in(far_4_4241_1[0]), .out(far_4_4241_2[0]));    relay_conn far_4_4241_2_b(.in(far_4_4241_1[1]), .out(far_4_4241_2[1]));
    assign layer_4[161] = ~(far_4_4241_2[0] | far_4_4241_2[1]); 
    assign layer_4[162] = layer_3[718] & ~layer_3[694]; 
    assign layer_4[163] = layer_3[116] | layer_3[134]; 
    assign layer_4[164] = layer_3[388] | layer_3[399]; 
    wire [1:0] far_4_4245_0;    relay_conn far_4_4245_0_a(.in(layer_3[255]), .out(far_4_4245_0[0]));    relay_conn far_4_4245_0_b(.in(layer_3[157]), .out(far_4_4245_0[1]));
    wire [1:0] far_4_4245_1;    relay_conn far_4_4245_1_a(.in(far_4_4245_0[0]), .out(far_4_4245_1[0]));    relay_conn far_4_4245_1_b(.in(far_4_4245_0[1]), .out(far_4_4245_1[1]));
    wire [1:0] far_4_4245_2;    relay_conn far_4_4245_2_a(.in(far_4_4245_1[0]), .out(far_4_4245_2[0]));    relay_conn far_4_4245_2_b(.in(far_4_4245_1[1]), .out(far_4_4245_2[1]));
    assign layer_4[165] = ~(far_4_4245_2[0] ^ far_4_4245_2[1]); 
    wire [1:0] far_4_4246_0;    relay_conn far_4_4246_0_a(.in(layer_3[861]), .out(far_4_4246_0[0]));    relay_conn far_4_4246_0_b(.in(layer_3[977]), .out(far_4_4246_0[1]));
    wire [1:0] far_4_4246_1;    relay_conn far_4_4246_1_a(.in(far_4_4246_0[0]), .out(far_4_4246_1[0]));    relay_conn far_4_4246_1_b(.in(far_4_4246_0[1]), .out(far_4_4246_1[1]));
    wire [1:0] far_4_4246_2;    relay_conn far_4_4246_2_a(.in(far_4_4246_1[0]), .out(far_4_4246_2[0]));    relay_conn far_4_4246_2_b(.in(far_4_4246_1[1]), .out(far_4_4246_2[1]));
    assign layer_4[166] = ~far_4_4246_2[0]; 
    wire [1:0] far_4_4247_0;    relay_conn far_4_4247_0_a(.in(layer_3[323]), .out(far_4_4247_0[0]));    relay_conn far_4_4247_0_b(.in(layer_3[281]), .out(far_4_4247_0[1]));
    assign layer_4[167] = ~far_4_4247_0[0]; 
    wire [1:0] far_4_4248_0;    relay_conn far_4_4248_0_a(.in(layer_3[110]), .out(far_4_4248_0[0]));    relay_conn far_4_4248_0_b(.in(layer_3[58]), .out(far_4_4248_0[1]));
    assign layer_4[168] = far_4_4248_0[0] | far_4_4248_0[1]; 
    wire [1:0] far_4_4249_0;    relay_conn far_4_4249_0_a(.in(layer_3[248]), .out(far_4_4249_0[0]));    relay_conn far_4_4249_0_b(.in(layer_3[137]), .out(far_4_4249_0[1]));
    wire [1:0] far_4_4249_1;    relay_conn far_4_4249_1_a(.in(far_4_4249_0[0]), .out(far_4_4249_1[0]));    relay_conn far_4_4249_1_b(.in(far_4_4249_0[1]), .out(far_4_4249_1[1]));
    wire [1:0] far_4_4249_2;    relay_conn far_4_4249_2_a(.in(far_4_4249_1[0]), .out(far_4_4249_2[0]));    relay_conn far_4_4249_2_b(.in(far_4_4249_1[1]), .out(far_4_4249_2[1]));
    assign layer_4[169] = far_4_4249_2[1] & ~far_4_4249_2[0]; 
    wire [1:0] far_4_4250_0;    relay_conn far_4_4250_0_a(.in(layer_3[686]), .out(far_4_4250_0[0]));    relay_conn far_4_4250_0_b(.in(layer_3[606]), .out(far_4_4250_0[1]));
    wire [1:0] far_4_4250_1;    relay_conn far_4_4250_1_a(.in(far_4_4250_0[0]), .out(far_4_4250_1[0]));    relay_conn far_4_4250_1_b(.in(far_4_4250_0[1]), .out(far_4_4250_1[1]));
    assign layer_4[170] = far_4_4250_1[0] & ~far_4_4250_1[1]; 
    assign layer_4[171] = ~layer_3[953] | (layer_3[953] & layer_3[958]); 
    wire [1:0] far_4_4252_0;    relay_conn far_4_4252_0_a(.in(layer_3[247]), .out(far_4_4252_0[0]));    relay_conn far_4_4252_0_b(.in(layer_3[364]), .out(far_4_4252_0[1]));
    wire [1:0] far_4_4252_1;    relay_conn far_4_4252_1_a(.in(far_4_4252_0[0]), .out(far_4_4252_1[0]));    relay_conn far_4_4252_1_b(.in(far_4_4252_0[1]), .out(far_4_4252_1[1]));
    wire [1:0] far_4_4252_2;    relay_conn far_4_4252_2_a(.in(far_4_4252_1[0]), .out(far_4_4252_2[0]));    relay_conn far_4_4252_2_b(.in(far_4_4252_1[1]), .out(far_4_4252_2[1]));
    assign layer_4[172] = far_4_4252_2[0] & far_4_4252_2[1]; 
    wire [1:0] far_4_4253_0;    relay_conn far_4_4253_0_a(.in(layer_3[149]), .out(far_4_4253_0[0]));    relay_conn far_4_4253_0_b(.in(layer_3[248]), .out(far_4_4253_0[1]));
    wire [1:0] far_4_4253_1;    relay_conn far_4_4253_1_a(.in(far_4_4253_0[0]), .out(far_4_4253_1[0]));    relay_conn far_4_4253_1_b(.in(far_4_4253_0[1]), .out(far_4_4253_1[1]));
    wire [1:0] far_4_4253_2;    relay_conn far_4_4253_2_a(.in(far_4_4253_1[0]), .out(far_4_4253_2[0]));    relay_conn far_4_4253_2_b(.in(far_4_4253_1[1]), .out(far_4_4253_2[1]));
    assign layer_4[173] = far_4_4253_2[0] & ~far_4_4253_2[1]; 
    wire [1:0] far_4_4254_0;    relay_conn far_4_4254_0_a(.in(layer_3[152]), .out(far_4_4254_0[0]));    relay_conn far_4_4254_0_b(.in(layer_3[118]), .out(far_4_4254_0[1]));
    assign layer_4[174] = far_4_4254_0[0] | far_4_4254_0[1]; 
    wire [1:0] far_4_4255_0;    relay_conn far_4_4255_0_a(.in(layer_3[253]), .out(far_4_4255_0[0]));    relay_conn far_4_4255_0_b(.in(layer_3[194]), .out(far_4_4255_0[1]));
    assign layer_4[175] = ~(far_4_4255_0[0] & far_4_4255_0[1]); 
    wire [1:0] far_4_4256_0;    relay_conn far_4_4256_0_a(.in(layer_3[787]), .out(far_4_4256_0[0]));    relay_conn far_4_4256_0_b(.in(layer_3[909]), .out(far_4_4256_0[1]));
    wire [1:0] far_4_4256_1;    relay_conn far_4_4256_1_a(.in(far_4_4256_0[0]), .out(far_4_4256_1[0]));    relay_conn far_4_4256_1_b(.in(far_4_4256_0[1]), .out(far_4_4256_1[1]));
    wire [1:0] far_4_4256_2;    relay_conn far_4_4256_2_a(.in(far_4_4256_1[0]), .out(far_4_4256_2[0]));    relay_conn far_4_4256_2_b(.in(far_4_4256_1[1]), .out(far_4_4256_2[1]));
    assign layer_4[176] = far_4_4256_2[1]; 
    wire [1:0] far_4_4257_0;    relay_conn far_4_4257_0_a(.in(layer_3[335]), .out(far_4_4257_0[0]));    relay_conn far_4_4257_0_b(.in(layer_3[375]), .out(far_4_4257_0[1]));
    assign layer_4[177] = ~(far_4_4257_0[0] | far_4_4257_0[1]); 
    wire [1:0] far_4_4258_0;    relay_conn far_4_4258_0_a(.in(layer_3[788]), .out(far_4_4258_0[0]));    relay_conn far_4_4258_0_b(.in(layer_3[734]), .out(far_4_4258_0[1]));
    assign layer_4[178] = far_4_4258_0[0] & ~far_4_4258_0[1]; 
    wire [1:0] far_4_4259_0;    relay_conn far_4_4259_0_a(.in(layer_3[83]), .out(far_4_4259_0[0]));    relay_conn far_4_4259_0_b(.in(layer_3[195]), .out(far_4_4259_0[1]));
    wire [1:0] far_4_4259_1;    relay_conn far_4_4259_1_a(.in(far_4_4259_0[0]), .out(far_4_4259_1[0]));    relay_conn far_4_4259_1_b(.in(far_4_4259_0[1]), .out(far_4_4259_1[1]));
    wire [1:0] far_4_4259_2;    relay_conn far_4_4259_2_a(.in(far_4_4259_1[0]), .out(far_4_4259_2[0]));    relay_conn far_4_4259_2_b(.in(far_4_4259_1[1]), .out(far_4_4259_2[1]));
    assign layer_4[179] = far_4_4259_2[0] & ~far_4_4259_2[1]; 
    wire [1:0] far_4_4260_0;    relay_conn far_4_4260_0_a(.in(layer_3[100]), .out(far_4_4260_0[0]));    relay_conn far_4_4260_0_b(.in(layer_3[40]), .out(far_4_4260_0[1]));
    assign layer_4[180] = ~far_4_4260_0[0] | (far_4_4260_0[0] & far_4_4260_0[1]); 
    wire [1:0] far_4_4261_0;    relay_conn far_4_4261_0_a(.in(layer_3[916]), .out(far_4_4261_0[0]));    relay_conn far_4_4261_0_b(.in(layer_3[838]), .out(far_4_4261_0[1]));
    wire [1:0] far_4_4261_1;    relay_conn far_4_4261_1_a(.in(far_4_4261_0[0]), .out(far_4_4261_1[0]));    relay_conn far_4_4261_1_b(.in(far_4_4261_0[1]), .out(far_4_4261_1[1]));
    assign layer_4[181] = ~(far_4_4261_1[0] ^ far_4_4261_1[1]); 
    wire [1:0] far_4_4262_0;    relay_conn far_4_4262_0_a(.in(layer_3[516]), .out(far_4_4262_0[0]));    relay_conn far_4_4262_0_b(.in(layer_3[559]), .out(far_4_4262_0[1]));
    assign layer_4[182] = ~far_4_4262_0[1] | (far_4_4262_0[0] & far_4_4262_0[1]); 
    assign layer_4[183] = ~layer_3[916]; 
    wire [1:0] far_4_4264_0;    relay_conn far_4_4264_0_a(.in(layer_3[686]), .out(far_4_4264_0[0]));    relay_conn far_4_4264_0_b(.in(layer_3[770]), .out(far_4_4264_0[1]));
    wire [1:0] far_4_4264_1;    relay_conn far_4_4264_1_a(.in(far_4_4264_0[0]), .out(far_4_4264_1[0]));    relay_conn far_4_4264_1_b(.in(far_4_4264_0[1]), .out(far_4_4264_1[1]));
    assign layer_4[184] = ~(far_4_4264_1[0] & far_4_4264_1[1]); 
    assign layer_4[185] = layer_3[304]; 
    wire [1:0] far_4_4266_0;    relay_conn far_4_4266_0_a(.in(layer_3[164]), .out(far_4_4266_0[0]));    relay_conn far_4_4266_0_b(.in(layer_3[274]), .out(far_4_4266_0[1]));
    wire [1:0] far_4_4266_1;    relay_conn far_4_4266_1_a(.in(far_4_4266_0[0]), .out(far_4_4266_1[0]));    relay_conn far_4_4266_1_b(.in(far_4_4266_0[1]), .out(far_4_4266_1[1]));
    wire [1:0] far_4_4266_2;    relay_conn far_4_4266_2_a(.in(far_4_4266_1[0]), .out(far_4_4266_2[0]));    relay_conn far_4_4266_2_b(.in(far_4_4266_1[1]), .out(far_4_4266_2[1]));
    assign layer_4[186] = ~(far_4_4266_2[0] & far_4_4266_2[1]); 
    wire [1:0] far_4_4267_0;    relay_conn far_4_4267_0_a(.in(layer_3[157]), .out(far_4_4267_0[0]));    relay_conn far_4_4267_0_b(.in(layer_3[57]), .out(far_4_4267_0[1]));
    wire [1:0] far_4_4267_1;    relay_conn far_4_4267_1_a(.in(far_4_4267_0[0]), .out(far_4_4267_1[0]));    relay_conn far_4_4267_1_b(.in(far_4_4267_0[1]), .out(far_4_4267_1[1]));
    wire [1:0] far_4_4267_2;    relay_conn far_4_4267_2_a(.in(far_4_4267_1[0]), .out(far_4_4267_2[0]));    relay_conn far_4_4267_2_b(.in(far_4_4267_1[1]), .out(far_4_4267_2[1]));
    assign layer_4[187] = far_4_4267_2[1]; 
    wire [1:0] far_4_4268_0;    relay_conn far_4_4268_0_a(.in(layer_3[360]), .out(far_4_4268_0[0]));    relay_conn far_4_4268_0_b(.in(layer_3[410]), .out(far_4_4268_0[1]));
    assign layer_4[188] = ~far_4_4268_0[0]; 
    assign layer_4[189] = ~layer_3[375]; 
    wire [1:0] far_4_4270_0;    relay_conn far_4_4270_0_a(.in(layer_3[648]), .out(far_4_4270_0[0]));    relay_conn far_4_4270_0_b(.in(layer_3[715]), .out(far_4_4270_0[1]));
    wire [1:0] far_4_4270_1;    relay_conn far_4_4270_1_a(.in(far_4_4270_0[0]), .out(far_4_4270_1[0]));    relay_conn far_4_4270_1_b(.in(far_4_4270_0[1]), .out(far_4_4270_1[1]));
    assign layer_4[190] = ~(far_4_4270_1[0] ^ far_4_4270_1[1]); 
    assign layer_4[191] = ~layer_3[916]; 
    wire [1:0] far_4_4272_0;    relay_conn far_4_4272_0_a(.in(layer_3[676]), .out(far_4_4272_0[0]));    relay_conn far_4_4272_0_b(.in(layer_3[791]), .out(far_4_4272_0[1]));
    wire [1:0] far_4_4272_1;    relay_conn far_4_4272_1_a(.in(far_4_4272_0[0]), .out(far_4_4272_1[0]));    relay_conn far_4_4272_1_b(.in(far_4_4272_0[1]), .out(far_4_4272_1[1]));
    wire [1:0] far_4_4272_2;    relay_conn far_4_4272_2_a(.in(far_4_4272_1[0]), .out(far_4_4272_2[0]));    relay_conn far_4_4272_2_b(.in(far_4_4272_1[1]), .out(far_4_4272_2[1]));
    assign layer_4[192] = far_4_4272_2[0] | far_4_4272_2[1]; 
    wire [1:0] far_4_4273_0;    relay_conn far_4_4273_0_a(.in(layer_3[774]), .out(far_4_4273_0[0]));    relay_conn far_4_4273_0_b(.in(layer_3[711]), .out(far_4_4273_0[1]));
    assign layer_4[193] = ~far_4_4273_0[0] | (far_4_4273_0[0] & far_4_4273_0[1]); 
    assign layer_4[194] = ~layer_3[314]; 
    assign layer_4[195] = layer_3[784] & ~layer_3[801]; 
    wire [1:0] far_4_4276_0;    relay_conn far_4_4276_0_a(.in(layer_3[154]), .out(far_4_4276_0[0]));    relay_conn far_4_4276_0_b(.in(layer_3[255]), .out(far_4_4276_0[1]));
    wire [1:0] far_4_4276_1;    relay_conn far_4_4276_1_a(.in(far_4_4276_0[0]), .out(far_4_4276_1[0]));    relay_conn far_4_4276_1_b(.in(far_4_4276_0[1]), .out(far_4_4276_1[1]));
    wire [1:0] far_4_4276_2;    relay_conn far_4_4276_2_a(.in(far_4_4276_1[0]), .out(far_4_4276_2[0]));    relay_conn far_4_4276_2_b(.in(far_4_4276_1[1]), .out(far_4_4276_2[1]));
    assign layer_4[196] = far_4_4276_2[1]; 
    assign layer_4[197] = layer_3[433] | layer_3[427]; 
    wire [1:0] far_4_4278_0;    relay_conn far_4_4278_0_a(.in(layer_3[896]), .out(far_4_4278_0[0]));    relay_conn far_4_4278_0_b(.in(layer_3[1004]), .out(far_4_4278_0[1]));
    wire [1:0] far_4_4278_1;    relay_conn far_4_4278_1_a(.in(far_4_4278_0[0]), .out(far_4_4278_1[0]));    relay_conn far_4_4278_1_b(.in(far_4_4278_0[1]), .out(far_4_4278_1[1]));
    wire [1:0] far_4_4278_2;    relay_conn far_4_4278_2_a(.in(far_4_4278_1[0]), .out(far_4_4278_2[0]));    relay_conn far_4_4278_2_b(.in(far_4_4278_1[1]), .out(far_4_4278_2[1]));
    assign layer_4[198] = far_4_4278_2[0]; 
    wire [1:0] far_4_4279_0;    relay_conn far_4_4279_0_a(.in(layer_3[171]), .out(far_4_4279_0[0]));    relay_conn far_4_4279_0_b(.in(layer_3[102]), .out(far_4_4279_0[1]));
    wire [1:0] far_4_4279_1;    relay_conn far_4_4279_1_a(.in(far_4_4279_0[0]), .out(far_4_4279_1[0]));    relay_conn far_4_4279_1_b(.in(far_4_4279_0[1]), .out(far_4_4279_1[1]));
    assign layer_4[199] = ~(far_4_4279_1[0] | far_4_4279_1[1]); 
    wire [1:0] far_4_4280_0;    relay_conn far_4_4280_0_a(.in(layer_3[879]), .out(far_4_4280_0[0]));    relay_conn far_4_4280_0_b(.in(layer_3[807]), .out(far_4_4280_0[1]));
    wire [1:0] far_4_4280_1;    relay_conn far_4_4280_1_a(.in(far_4_4280_0[0]), .out(far_4_4280_1[0]));    relay_conn far_4_4280_1_b(.in(far_4_4280_0[1]), .out(far_4_4280_1[1]));
    assign layer_4[200] = far_4_4280_1[0] & ~far_4_4280_1[1]; 
    assign layer_4[201] = layer_3[599] & ~layer_3[625]; 
    wire [1:0] far_4_4282_0;    relay_conn far_4_4282_0_a(.in(layer_3[454]), .out(far_4_4282_0[0]));    relay_conn far_4_4282_0_b(.in(layer_3[486]), .out(far_4_4282_0[1]));
    assign layer_4[202] = ~far_4_4282_0[0]; 
    wire [1:0] far_4_4283_0;    relay_conn far_4_4283_0_a(.in(layer_3[346]), .out(far_4_4283_0[0]));    relay_conn far_4_4283_0_b(.in(layer_3[455]), .out(far_4_4283_0[1]));
    wire [1:0] far_4_4283_1;    relay_conn far_4_4283_1_a(.in(far_4_4283_0[0]), .out(far_4_4283_1[0]));    relay_conn far_4_4283_1_b(.in(far_4_4283_0[1]), .out(far_4_4283_1[1]));
    wire [1:0] far_4_4283_2;    relay_conn far_4_4283_2_a(.in(far_4_4283_1[0]), .out(far_4_4283_2[0]));    relay_conn far_4_4283_2_b(.in(far_4_4283_1[1]), .out(far_4_4283_2[1]));
    assign layer_4[203] = far_4_4283_2[0] & ~far_4_4283_2[1]; 
    assign layer_4[204] = layer_3[64] ^ layer_3[37]; 
    wire [1:0] far_4_4285_0;    relay_conn far_4_4285_0_a(.in(layer_3[885]), .out(far_4_4285_0[0]));    relay_conn far_4_4285_0_b(.in(layer_3[831]), .out(far_4_4285_0[1]));
    assign layer_4[205] = ~far_4_4285_0[1] | (far_4_4285_0[0] & far_4_4285_0[1]); 
    assign layer_4[206] = ~layer_3[314]; 
    wire [1:0] far_4_4287_0;    relay_conn far_4_4287_0_a(.in(layer_3[160]), .out(far_4_4287_0[0]));    relay_conn far_4_4287_0_b(.in(layer_3[115]), .out(far_4_4287_0[1]));
    assign layer_4[207] = far_4_4287_0[1] & ~far_4_4287_0[0]; 
    wire [1:0] far_4_4288_0;    relay_conn far_4_4288_0_a(.in(layer_3[544]), .out(far_4_4288_0[0]));    relay_conn far_4_4288_0_b(.in(layer_3[446]), .out(far_4_4288_0[1]));
    wire [1:0] far_4_4288_1;    relay_conn far_4_4288_1_a(.in(far_4_4288_0[0]), .out(far_4_4288_1[0]));    relay_conn far_4_4288_1_b(.in(far_4_4288_0[1]), .out(far_4_4288_1[1]));
    wire [1:0] far_4_4288_2;    relay_conn far_4_4288_2_a(.in(far_4_4288_1[0]), .out(far_4_4288_2[0]));    relay_conn far_4_4288_2_b(.in(far_4_4288_1[1]), .out(far_4_4288_2[1]));
    assign layer_4[208] = far_4_4288_2[0] ^ far_4_4288_2[1]; 
    wire [1:0] far_4_4289_0;    relay_conn far_4_4289_0_a(.in(layer_3[138]), .out(far_4_4289_0[0]));    relay_conn far_4_4289_0_b(.in(layer_3[35]), .out(far_4_4289_0[1]));
    wire [1:0] far_4_4289_1;    relay_conn far_4_4289_1_a(.in(far_4_4289_0[0]), .out(far_4_4289_1[0]));    relay_conn far_4_4289_1_b(.in(far_4_4289_0[1]), .out(far_4_4289_1[1]));
    wire [1:0] far_4_4289_2;    relay_conn far_4_4289_2_a(.in(far_4_4289_1[0]), .out(far_4_4289_2[0]));    relay_conn far_4_4289_2_b(.in(far_4_4289_1[1]), .out(far_4_4289_2[1]));
    assign layer_4[209] = far_4_4289_2[0] & far_4_4289_2[1]; 
    wire [1:0] far_4_4290_0;    relay_conn far_4_4290_0_a(.in(layer_3[544]), .out(far_4_4290_0[0]));    relay_conn far_4_4290_0_b(.in(layer_3[664]), .out(far_4_4290_0[1]));
    wire [1:0] far_4_4290_1;    relay_conn far_4_4290_1_a(.in(far_4_4290_0[0]), .out(far_4_4290_1[0]));    relay_conn far_4_4290_1_b(.in(far_4_4290_0[1]), .out(far_4_4290_1[1]));
    wire [1:0] far_4_4290_2;    relay_conn far_4_4290_2_a(.in(far_4_4290_1[0]), .out(far_4_4290_2[0]));    relay_conn far_4_4290_2_b(.in(far_4_4290_1[1]), .out(far_4_4290_2[1]));
    assign layer_4[210] = far_4_4290_2[0] | far_4_4290_2[1]; 
    wire [1:0] far_4_4291_0;    relay_conn far_4_4291_0_a(.in(layer_3[37]), .out(far_4_4291_0[0]));    relay_conn far_4_4291_0_b(.in(layer_3[128]), .out(far_4_4291_0[1]));
    wire [1:0] far_4_4291_1;    relay_conn far_4_4291_1_a(.in(far_4_4291_0[0]), .out(far_4_4291_1[0]));    relay_conn far_4_4291_1_b(.in(far_4_4291_0[1]), .out(far_4_4291_1[1]));
    assign layer_4[211] = far_4_4291_1[0]; 
    wire [1:0] far_4_4292_0;    relay_conn far_4_4292_0_a(.in(layer_3[968]), .out(far_4_4292_0[0]));    relay_conn far_4_4292_0_b(.in(layer_3[1009]), .out(far_4_4292_0[1]));
    assign layer_4[212] = ~(far_4_4292_0[0] & far_4_4292_0[1]); 
    wire [1:0] far_4_4293_0;    relay_conn far_4_4293_0_a(.in(layer_3[488]), .out(far_4_4293_0[0]));    relay_conn far_4_4293_0_b(.in(layer_3[567]), .out(far_4_4293_0[1]));
    wire [1:0] far_4_4293_1;    relay_conn far_4_4293_1_a(.in(far_4_4293_0[0]), .out(far_4_4293_1[0]));    relay_conn far_4_4293_1_b(.in(far_4_4293_0[1]), .out(far_4_4293_1[1]));
    assign layer_4[213] = ~(far_4_4293_1[0] & far_4_4293_1[1]); 
    wire [1:0] far_4_4294_0;    relay_conn far_4_4294_0_a(.in(layer_3[41]), .out(far_4_4294_0[0]));    relay_conn far_4_4294_0_b(.in(layer_3[80]), .out(far_4_4294_0[1]));
    assign layer_4[214] = far_4_4294_0[0] | far_4_4294_0[1]; 
    wire [1:0] far_4_4295_0;    relay_conn far_4_4295_0_a(.in(layer_3[950]), .out(far_4_4295_0[0]));    relay_conn far_4_4295_0_b(.in(layer_3[898]), .out(far_4_4295_0[1]));
    assign layer_4[215] = far_4_4295_0[0]; 
    wire [1:0] far_4_4296_0;    relay_conn far_4_4296_0_a(.in(layer_3[206]), .out(far_4_4296_0[0]));    relay_conn far_4_4296_0_b(.in(layer_3[79]), .out(far_4_4296_0[1]));
    wire [1:0] far_4_4296_1;    relay_conn far_4_4296_1_a(.in(far_4_4296_0[0]), .out(far_4_4296_1[0]));    relay_conn far_4_4296_1_b(.in(far_4_4296_0[1]), .out(far_4_4296_1[1]));
    wire [1:0] far_4_4296_2;    relay_conn far_4_4296_2_a(.in(far_4_4296_1[0]), .out(far_4_4296_2[0]));    relay_conn far_4_4296_2_b(.in(far_4_4296_1[1]), .out(far_4_4296_2[1]));
    assign layer_4[216] = far_4_4296_2[0] ^ far_4_4296_2[1]; 
    wire [1:0] far_4_4297_0;    relay_conn far_4_4297_0_a(.in(layer_3[105]), .out(far_4_4297_0[0]));    relay_conn far_4_4297_0_b(.in(layer_3[153]), .out(far_4_4297_0[1]));
    assign layer_4[217] = ~(far_4_4297_0[0] & far_4_4297_0[1]); 
    wire [1:0] far_4_4298_0;    relay_conn far_4_4298_0_a(.in(layer_3[367]), .out(far_4_4298_0[0]));    relay_conn far_4_4298_0_b(.in(layer_3[271]), .out(far_4_4298_0[1]));
    wire [1:0] far_4_4298_1;    relay_conn far_4_4298_1_a(.in(far_4_4298_0[0]), .out(far_4_4298_1[0]));    relay_conn far_4_4298_1_b(.in(far_4_4298_0[1]), .out(far_4_4298_1[1]));
    wire [1:0] far_4_4298_2;    relay_conn far_4_4298_2_a(.in(far_4_4298_1[0]), .out(far_4_4298_2[0]));    relay_conn far_4_4298_2_b(.in(far_4_4298_1[1]), .out(far_4_4298_2[1]));
    assign layer_4[218] = ~far_4_4298_2[0] | (far_4_4298_2[0] & far_4_4298_2[1]); 
    assign layer_4[219] = ~layer_3[756] | (layer_3[756] & layer_3[772]); 
    wire [1:0] far_4_4300_0;    relay_conn far_4_4300_0_a(.in(layer_3[218]), .out(far_4_4300_0[0]));    relay_conn far_4_4300_0_b(.in(layer_3[336]), .out(far_4_4300_0[1]));
    wire [1:0] far_4_4300_1;    relay_conn far_4_4300_1_a(.in(far_4_4300_0[0]), .out(far_4_4300_1[0]));    relay_conn far_4_4300_1_b(.in(far_4_4300_0[1]), .out(far_4_4300_1[1]));
    wire [1:0] far_4_4300_2;    relay_conn far_4_4300_2_a(.in(far_4_4300_1[0]), .out(far_4_4300_2[0]));    relay_conn far_4_4300_2_b(.in(far_4_4300_1[1]), .out(far_4_4300_2[1]));
    assign layer_4[220] = far_4_4300_2[0] ^ far_4_4300_2[1]; 
    assign layer_4[221] = layer_3[36] | layer_3[5]; 
    wire [1:0] far_4_4302_0;    relay_conn far_4_4302_0_a(.in(layer_3[673]), .out(far_4_4302_0[0]));    relay_conn far_4_4302_0_b(.in(layer_3[734]), .out(far_4_4302_0[1]));
    assign layer_4[222] = ~far_4_4302_0[1] | (far_4_4302_0[0] & far_4_4302_0[1]); 
    assign layer_4[223] = ~layer_3[756] | (layer_3[756] & layer_3[725]); 
    wire [1:0] far_4_4304_0;    relay_conn far_4_4304_0_a(.in(layer_3[894]), .out(far_4_4304_0[0]));    relay_conn far_4_4304_0_b(.in(layer_3[950]), .out(far_4_4304_0[1]));
    assign layer_4[224] = ~far_4_4304_0[1]; 
    wire [1:0] far_4_4305_0;    relay_conn far_4_4305_0_a(.in(layer_3[332]), .out(far_4_4305_0[0]));    relay_conn far_4_4305_0_b(.in(layer_3[394]), .out(far_4_4305_0[1]));
    assign layer_4[225] = ~(far_4_4305_0[0] | far_4_4305_0[1]); 
    wire [1:0] far_4_4306_0;    relay_conn far_4_4306_0_a(.in(layer_3[555]), .out(far_4_4306_0[0]));    relay_conn far_4_4306_0_b(.in(layer_3[676]), .out(far_4_4306_0[1]));
    wire [1:0] far_4_4306_1;    relay_conn far_4_4306_1_a(.in(far_4_4306_0[0]), .out(far_4_4306_1[0]));    relay_conn far_4_4306_1_b(.in(far_4_4306_0[1]), .out(far_4_4306_1[1]));
    wire [1:0] far_4_4306_2;    relay_conn far_4_4306_2_a(.in(far_4_4306_1[0]), .out(far_4_4306_2[0]));    relay_conn far_4_4306_2_b(.in(far_4_4306_1[1]), .out(far_4_4306_2[1]));
    assign layer_4[226] = ~far_4_4306_2[1] | (far_4_4306_2[0] & far_4_4306_2[1]); 
    assign layer_4[227] = ~(layer_3[630] & layer_3[611]); 
    wire [1:0] far_4_4308_0;    relay_conn far_4_4308_0_a(.in(layer_3[507]), .out(far_4_4308_0[0]));    relay_conn far_4_4308_0_b(.in(layer_3[391]), .out(far_4_4308_0[1]));
    wire [1:0] far_4_4308_1;    relay_conn far_4_4308_1_a(.in(far_4_4308_0[0]), .out(far_4_4308_1[0]));    relay_conn far_4_4308_1_b(.in(far_4_4308_0[1]), .out(far_4_4308_1[1]));
    wire [1:0] far_4_4308_2;    relay_conn far_4_4308_2_a(.in(far_4_4308_1[0]), .out(far_4_4308_2[0]));    relay_conn far_4_4308_2_b(.in(far_4_4308_1[1]), .out(far_4_4308_2[1]));
    assign layer_4[228] = far_4_4308_2[0]; 
    assign layer_4[229] = layer_3[320] & ~layer_3[331]; 
    wire [1:0] far_4_4310_0;    relay_conn far_4_4310_0_a(.in(layer_3[903]), .out(far_4_4310_0[0]));    relay_conn far_4_4310_0_b(.in(layer_3[953]), .out(far_4_4310_0[1]));
    assign layer_4[230] = far_4_4310_0[0] ^ far_4_4310_0[1]; 
    wire [1:0] far_4_4311_0;    relay_conn far_4_4311_0_a(.in(layer_3[101]), .out(far_4_4311_0[0]));    relay_conn far_4_4311_0_b(.in(layer_3[192]), .out(far_4_4311_0[1]));
    wire [1:0] far_4_4311_1;    relay_conn far_4_4311_1_a(.in(far_4_4311_0[0]), .out(far_4_4311_1[0]));    relay_conn far_4_4311_1_b(.in(far_4_4311_0[1]), .out(far_4_4311_1[1]));
    assign layer_4[231] = far_4_4311_1[0]; 
    wire [1:0] far_4_4312_0;    relay_conn far_4_4312_0_a(.in(layer_3[831]), .out(far_4_4312_0[0]));    relay_conn far_4_4312_0_b(.in(layer_3[948]), .out(far_4_4312_0[1]));
    wire [1:0] far_4_4312_1;    relay_conn far_4_4312_1_a(.in(far_4_4312_0[0]), .out(far_4_4312_1[0]));    relay_conn far_4_4312_1_b(.in(far_4_4312_0[1]), .out(far_4_4312_1[1]));
    wire [1:0] far_4_4312_2;    relay_conn far_4_4312_2_a(.in(far_4_4312_1[0]), .out(far_4_4312_2[0]));    relay_conn far_4_4312_2_b(.in(far_4_4312_1[1]), .out(far_4_4312_2[1]));
    assign layer_4[232] = ~(far_4_4312_2[0] | far_4_4312_2[1]); 
    wire [1:0] far_4_4313_0;    relay_conn far_4_4313_0_a(.in(layer_3[321]), .out(far_4_4313_0[0]));    relay_conn far_4_4313_0_b(.in(layer_3[289]), .out(far_4_4313_0[1]));
    assign layer_4[233] = far_4_4313_0[0] & far_4_4313_0[1]; 
    wire [1:0] far_4_4314_0;    relay_conn far_4_4314_0_a(.in(layer_3[400]), .out(far_4_4314_0[0]));    relay_conn far_4_4314_0_b(.in(layer_3[317]), .out(far_4_4314_0[1]));
    wire [1:0] far_4_4314_1;    relay_conn far_4_4314_1_a(.in(far_4_4314_0[0]), .out(far_4_4314_1[0]));    relay_conn far_4_4314_1_b(.in(far_4_4314_0[1]), .out(far_4_4314_1[1]));
    assign layer_4[234] = far_4_4314_1[0] ^ far_4_4314_1[1]; 
    assign layer_4[235] = ~layer_3[681]; 
    wire [1:0] far_4_4316_0;    relay_conn far_4_4316_0_a(.in(layer_3[36]), .out(far_4_4316_0[0]));    relay_conn far_4_4316_0_b(.in(layer_3[75]), .out(far_4_4316_0[1]));
    assign layer_4[236] = far_4_4316_0[0] | far_4_4316_0[1]; 
    wire [1:0] far_4_4317_0;    relay_conn far_4_4317_0_a(.in(layer_3[323]), .out(far_4_4317_0[0]));    relay_conn far_4_4317_0_b(.in(layer_3[394]), .out(far_4_4317_0[1]));
    wire [1:0] far_4_4317_1;    relay_conn far_4_4317_1_a(.in(far_4_4317_0[0]), .out(far_4_4317_1[0]));    relay_conn far_4_4317_1_b(.in(far_4_4317_0[1]), .out(far_4_4317_1[1]));
    assign layer_4[237] = ~far_4_4317_1[1]; 
    assign layer_4[238] = layer_3[396] ^ layer_3[391]; 
    wire [1:0] far_4_4319_0;    relay_conn far_4_4319_0_a(.in(layer_3[329]), .out(far_4_4319_0[0]));    relay_conn far_4_4319_0_b(.in(layer_3[383]), .out(far_4_4319_0[1]));
    assign layer_4[239] = ~(far_4_4319_0[0] | far_4_4319_0[1]); 
    assign layer_4[240] = layer_3[440] & ~layer_3[424]; 
    assign layer_4[241] = layer_3[100] & ~layer_3[77]; 
    wire [1:0] far_4_4322_0;    relay_conn far_4_4322_0_a(.in(layer_3[2]), .out(far_4_4322_0[0]));    relay_conn far_4_4322_0_b(.in(layer_3[105]), .out(far_4_4322_0[1]));
    wire [1:0] far_4_4322_1;    relay_conn far_4_4322_1_a(.in(far_4_4322_0[0]), .out(far_4_4322_1[0]));    relay_conn far_4_4322_1_b(.in(far_4_4322_0[1]), .out(far_4_4322_1[1]));
    wire [1:0] far_4_4322_2;    relay_conn far_4_4322_2_a(.in(far_4_4322_1[0]), .out(far_4_4322_2[0]));    relay_conn far_4_4322_2_b(.in(far_4_4322_1[1]), .out(far_4_4322_2[1]));
    assign layer_4[242] = far_4_4322_2[0] & ~far_4_4322_2[1]; 
    wire [1:0] far_4_4323_0;    relay_conn far_4_4323_0_a(.in(layer_3[542]), .out(far_4_4323_0[0]));    relay_conn far_4_4323_0_b(.in(layer_3[414]), .out(far_4_4323_0[1]));
    wire [1:0] far_4_4323_1;    relay_conn far_4_4323_1_a(.in(far_4_4323_0[0]), .out(far_4_4323_1[0]));    relay_conn far_4_4323_1_b(.in(far_4_4323_0[1]), .out(far_4_4323_1[1]));
    wire [1:0] far_4_4323_2;    relay_conn far_4_4323_2_a(.in(far_4_4323_1[0]), .out(far_4_4323_2[0]));    relay_conn far_4_4323_2_b(.in(far_4_4323_1[1]), .out(far_4_4323_2[1]));
    wire [1:0] far_4_4323_3;    relay_conn far_4_4323_3_a(.in(far_4_4323_2[0]), .out(far_4_4323_3[0]));    relay_conn far_4_4323_3_b(.in(far_4_4323_2[1]), .out(far_4_4323_3[1]));
    assign layer_4[243] = far_4_4323_3[1] & ~far_4_4323_3[0]; 
    assign layer_4[244] = ~layer_3[855]; 
    wire [1:0] far_4_4325_0;    relay_conn far_4_4325_0_a(.in(layer_3[473]), .out(far_4_4325_0[0]));    relay_conn far_4_4325_0_b(.in(layer_3[400]), .out(far_4_4325_0[1]));
    wire [1:0] far_4_4325_1;    relay_conn far_4_4325_1_a(.in(far_4_4325_0[0]), .out(far_4_4325_1[0]));    relay_conn far_4_4325_1_b(.in(far_4_4325_0[1]), .out(far_4_4325_1[1]));
    assign layer_4[245] = far_4_4325_1[0] & ~far_4_4325_1[1]; 
    wire [1:0] far_4_4326_0;    relay_conn far_4_4326_0_a(.in(layer_3[529]), .out(far_4_4326_0[0]));    relay_conn far_4_4326_0_b(.in(layer_3[486]), .out(far_4_4326_0[1]));
    assign layer_4[246] = far_4_4326_0[0] & ~far_4_4326_0[1]; 
    wire [1:0] far_4_4327_0;    relay_conn far_4_4327_0_a(.in(layer_3[977]), .out(far_4_4327_0[0]));    relay_conn far_4_4327_0_b(.in(layer_3[910]), .out(far_4_4327_0[1]));
    wire [1:0] far_4_4327_1;    relay_conn far_4_4327_1_a(.in(far_4_4327_0[0]), .out(far_4_4327_1[0]));    relay_conn far_4_4327_1_b(.in(far_4_4327_0[1]), .out(far_4_4327_1[1]));
    assign layer_4[247] = far_4_4327_1[0]; 
    wire [1:0] far_4_4328_0;    relay_conn far_4_4328_0_a(.in(layer_3[92]), .out(far_4_4328_0[0]));    relay_conn far_4_4328_0_b(.in(layer_3[161]), .out(far_4_4328_0[1]));
    wire [1:0] far_4_4328_1;    relay_conn far_4_4328_1_a(.in(far_4_4328_0[0]), .out(far_4_4328_1[0]));    relay_conn far_4_4328_1_b(.in(far_4_4328_0[1]), .out(far_4_4328_1[1]));
    assign layer_4[248] = far_4_4328_1[1] & ~far_4_4328_1[0]; 
    wire [1:0] far_4_4329_0;    relay_conn far_4_4329_0_a(.in(layer_3[72]), .out(far_4_4329_0[0]));    relay_conn far_4_4329_0_b(.in(layer_3[36]), .out(far_4_4329_0[1]));
    assign layer_4[249] = ~(far_4_4329_0[0] & far_4_4329_0[1]); 
    wire [1:0] far_4_4330_0;    relay_conn far_4_4330_0_a(.in(layer_3[405]), .out(far_4_4330_0[0]));    relay_conn far_4_4330_0_b(.in(layer_3[279]), .out(far_4_4330_0[1]));
    wire [1:0] far_4_4330_1;    relay_conn far_4_4330_1_a(.in(far_4_4330_0[0]), .out(far_4_4330_1[0]));    relay_conn far_4_4330_1_b(.in(far_4_4330_0[1]), .out(far_4_4330_1[1]));
    wire [1:0] far_4_4330_2;    relay_conn far_4_4330_2_a(.in(far_4_4330_1[0]), .out(far_4_4330_2[0]));    relay_conn far_4_4330_2_b(.in(far_4_4330_1[1]), .out(far_4_4330_2[1]));
    assign layer_4[250] = far_4_4330_2[0] & far_4_4330_2[1]; 
    assign layer_4[251] = layer_3[905] & ~layer_3[935]; 
    assign layer_4[252] = ~layer_3[232]; 
    wire [1:0] far_4_4333_0;    relay_conn far_4_4333_0_a(.in(layer_3[688]), .out(far_4_4333_0[0]));    relay_conn far_4_4333_0_b(.in(layer_3[784]), .out(far_4_4333_0[1]));
    wire [1:0] far_4_4333_1;    relay_conn far_4_4333_1_a(.in(far_4_4333_0[0]), .out(far_4_4333_1[0]));    relay_conn far_4_4333_1_b(.in(far_4_4333_0[1]), .out(far_4_4333_1[1]));
    wire [1:0] far_4_4333_2;    relay_conn far_4_4333_2_a(.in(far_4_4333_1[0]), .out(far_4_4333_2[0]));    relay_conn far_4_4333_2_b(.in(far_4_4333_1[1]), .out(far_4_4333_2[1]));
    assign layer_4[253] = far_4_4333_2[0] | far_4_4333_2[1]; 
    wire [1:0] far_4_4334_0;    relay_conn far_4_4334_0_a(.in(layer_3[896]), .out(far_4_4334_0[0]));    relay_conn far_4_4334_0_b(.in(layer_3[1009]), .out(far_4_4334_0[1]));
    wire [1:0] far_4_4334_1;    relay_conn far_4_4334_1_a(.in(far_4_4334_0[0]), .out(far_4_4334_1[0]));    relay_conn far_4_4334_1_b(.in(far_4_4334_0[1]), .out(far_4_4334_1[1]));
    wire [1:0] far_4_4334_2;    relay_conn far_4_4334_2_a(.in(far_4_4334_1[0]), .out(far_4_4334_2[0]));    relay_conn far_4_4334_2_b(.in(far_4_4334_1[1]), .out(far_4_4334_2[1]));
    assign layer_4[254] = far_4_4334_2[1] & ~far_4_4334_2[0]; 
    wire [1:0] far_4_4335_0;    relay_conn far_4_4335_0_a(.in(layer_3[352]), .out(far_4_4335_0[0]));    relay_conn far_4_4335_0_b(.in(layer_3[251]), .out(far_4_4335_0[1]));
    wire [1:0] far_4_4335_1;    relay_conn far_4_4335_1_a(.in(far_4_4335_0[0]), .out(far_4_4335_1[0]));    relay_conn far_4_4335_1_b(.in(far_4_4335_0[1]), .out(far_4_4335_1[1]));
    wire [1:0] far_4_4335_2;    relay_conn far_4_4335_2_a(.in(far_4_4335_1[0]), .out(far_4_4335_2[0]));    relay_conn far_4_4335_2_b(.in(far_4_4335_1[1]), .out(far_4_4335_2[1]));
    assign layer_4[255] = far_4_4335_2[0] ^ far_4_4335_2[1]; 
    wire [1:0] far_4_4336_0;    relay_conn far_4_4336_0_a(.in(layer_3[830]), .out(far_4_4336_0[0]));    relay_conn far_4_4336_0_b(.in(layer_3[766]), .out(far_4_4336_0[1]));
    wire [1:0] far_4_4336_1;    relay_conn far_4_4336_1_a(.in(far_4_4336_0[0]), .out(far_4_4336_1[0]));    relay_conn far_4_4336_1_b(.in(far_4_4336_0[1]), .out(far_4_4336_1[1]));
    assign layer_4[256] = far_4_4336_1[0] | far_4_4336_1[1]; 
    wire [1:0] far_4_4337_0;    relay_conn far_4_4337_0_a(.in(layer_3[127]), .out(far_4_4337_0[0]));    relay_conn far_4_4337_0_b(.in(layer_3[37]), .out(far_4_4337_0[1]));
    wire [1:0] far_4_4337_1;    relay_conn far_4_4337_1_a(.in(far_4_4337_0[0]), .out(far_4_4337_1[0]));    relay_conn far_4_4337_1_b(.in(far_4_4337_0[1]), .out(far_4_4337_1[1]));
    assign layer_4[257] = far_4_4337_1[1]; 
    wire [1:0] far_4_4338_0;    relay_conn far_4_4338_0_a(.in(layer_3[985]), .out(far_4_4338_0[0]));    relay_conn far_4_4338_0_b(.in(layer_3[870]), .out(far_4_4338_0[1]));
    wire [1:0] far_4_4338_1;    relay_conn far_4_4338_1_a(.in(far_4_4338_0[0]), .out(far_4_4338_1[0]));    relay_conn far_4_4338_1_b(.in(far_4_4338_0[1]), .out(far_4_4338_1[1]));
    wire [1:0] far_4_4338_2;    relay_conn far_4_4338_2_a(.in(far_4_4338_1[0]), .out(far_4_4338_2[0]));    relay_conn far_4_4338_2_b(.in(far_4_4338_1[1]), .out(far_4_4338_2[1]));
    assign layer_4[258] = ~(far_4_4338_2[0] & far_4_4338_2[1]); 
    wire [1:0] far_4_4339_0;    relay_conn far_4_4339_0_a(.in(layer_3[495]), .out(far_4_4339_0[0]));    relay_conn far_4_4339_0_b(.in(layer_3[576]), .out(far_4_4339_0[1]));
    wire [1:0] far_4_4339_1;    relay_conn far_4_4339_1_a(.in(far_4_4339_0[0]), .out(far_4_4339_1[0]));    relay_conn far_4_4339_1_b(.in(far_4_4339_0[1]), .out(far_4_4339_1[1]));
    assign layer_4[259] = ~(far_4_4339_1[0] ^ far_4_4339_1[1]); 
    assign layer_4[260] = ~layer_3[411]; 
    wire [1:0] far_4_4341_0;    relay_conn far_4_4341_0_a(.in(layer_3[762]), .out(far_4_4341_0[0]));    relay_conn far_4_4341_0_b(.in(layer_3[880]), .out(far_4_4341_0[1]));
    wire [1:0] far_4_4341_1;    relay_conn far_4_4341_1_a(.in(far_4_4341_0[0]), .out(far_4_4341_1[0]));    relay_conn far_4_4341_1_b(.in(far_4_4341_0[1]), .out(far_4_4341_1[1]));
    wire [1:0] far_4_4341_2;    relay_conn far_4_4341_2_a(.in(far_4_4341_1[0]), .out(far_4_4341_2[0]));    relay_conn far_4_4341_2_b(.in(far_4_4341_1[1]), .out(far_4_4341_2[1]));
    assign layer_4[261] = far_4_4341_2[0]; 
    wire [1:0] far_4_4342_0;    relay_conn far_4_4342_0_a(.in(layer_3[299]), .out(far_4_4342_0[0]));    relay_conn far_4_4342_0_b(.in(layer_3[424]), .out(far_4_4342_0[1]));
    wire [1:0] far_4_4342_1;    relay_conn far_4_4342_1_a(.in(far_4_4342_0[0]), .out(far_4_4342_1[0]));    relay_conn far_4_4342_1_b(.in(far_4_4342_0[1]), .out(far_4_4342_1[1]));
    wire [1:0] far_4_4342_2;    relay_conn far_4_4342_2_a(.in(far_4_4342_1[0]), .out(far_4_4342_2[0]));    relay_conn far_4_4342_2_b(.in(far_4_4342_1[1]), .out(far_4_4342_2[1]));
    assign layer_4[262] = ~far_4_4342_2[0] | (far_4_4342_2[0] & far_4_4342_2[1]); 
    wire [1:0] far_4_4343_0;    relay_conn far_4_4343_0_a(.in(layer_3[876]), .out(far_4_4343_0[0]));    relay_conn far_4_4343_0_b(.in(layer_3[934]), .out(far_4_4343_0[1]));
    assign layer_4[263] = ~far_4_4343_0[0]; 
    wire [1:0] far_4_4344_0;    relay_conn far_4_4344_0_a(.in(layer_3[820]), .out(far_4_4344_0[0]));    relay_conn far_4_4344_0_b(.in(layer_3[869]), .out(far_4_4344_0[1]));
    assign layer_4[264] = ~far_4_4344_0[1]; 
    wire [1:0] far_4_4345_0;    relay_conn far_4_4345_0_a(.in(layer_3[638]), .out(far_4_4345_0[0]));    relay_conn far_4_4345_0_b(.in(layer_3[756]), .out(far_4_4345_0[1]));
    wire [1:0] far_4_4345_1;    relay_conn far_4_4345_1_a(.in(far_4_4345_0[0]), .out(far_4_4345_1[0]));    relay_conn far_4_4345_1_b(.in(far_4_4345_0[1]), .out(far_4_4345_1[1]));
    wire [1:0] far_4_4345_2;    relay_conn far_4_4345_2_a(.in(far_4_4345_1[0]), .out(far_4_4345_2[0]));    relay_conn far_4_4345_2_b(.in(far_4_4345_1[1]), .out(far_4_4345_2[1]));
    assign layer_4[265] = far_4_4345_2[1]; 
    wire [1:0] far_4_4346_0;    relay_conn far_4_4346_0_a(.in(layer_3[325]), .out(far_4_4346_0[0]));    relay_conn far_4_4346_0_b(.in(layer_3[222]), .out(far_4_4346_0[1]));
    wire [1:0] far_4_4346_1;    relay_conn far_4_4346_1_a(.in(far_4_4346_0[0]), .out(far_4_4346_1[0]));    relay_conn far_4_4346_1_b(.in(far_4_4346_0[1]), .out(far_4_4346_1[1]));
    wire [1:0] far_4_4346_2;    relay_conn far_4_4346_2_a(.in(far_4_4346_1[0]), .out(far_4_4346_2[0]));    relay_conn far_4_4346_2_b(.in(far_4_4346_1[1]), .out(far_4_4346_2[1]));
    assign layer_4[266] = ~far_4_4346_2[1]; 
    wire [1:0] far_4_4347_0;    relay_conn far_4_4347_0_a(.in(layer_3[191]), .out(far_4_4347_0[0]));    relay_conn far_4_4347_0_b(.in(layer_3[85]), .out(far_4_4347_0[1]));
    wire [1:0] far_4_4347_1;    relay_conn far_4_4347_1_a(.in(far_4_4347_0[0]), .out(far_4_4347_1[0]));    relay_conn far_4_4347_1_b(.in(far_4_4347_0[1]), .out(far_4_4347_1[1]));
    wire [1:0] far_4_4347_2;    relay_conn far_4_4347_2_a(.in(far_4_4347_1[0]), .out(far_4_4347_2[0]));    relay_conn far_4_4347_2_b(.in(far_4_4347_1[1]), .out(far_4_4347_2[1]));
    assign layer_4[267] = ~far_4_4347_2[0] | (far_4_4347_2[0] & far_4_4347_2[1]); 
    assign layer_4[268] = ~layer_3[140]; 
    assign layer_4[269] = ~layer_3[362]; 
    wire [1:0] far_4_4350_0;    relay_conn far_4_4350_0_a(.in(layer_3[265]), .out(far_4_4350_0[0]));    relay_conn far_4_4350_0_b(.in(layer_3[323]), .out(far_4_4350_0[1]));
    assign layer_4[270] = far_4_4350_0[0] ^ far_4_4350_0[1]; 
    wire [1:0] far_4_4351_0;    relay_conn far_4_4351_0_a(.in(layer_3[37]), .out(far_4_4351_0[0]));    relay_conn far_4_4351_0_b(.in(layer_3[100]), .out(far_4_4351_0[1]));
    assign layer_4[271] = far_4_4351_0[0]; 
    wire [1:0] far_4_4352_0;    relay_conn far_4_4352_0_a(.in(layer_3[415]), .out(far_4_4352_0[0]));    relay_conn far_4_4352_0_b(.in(layer_3[481]), .out(far_4_4352_0[1]));
    wire [1:0] far_4_4352_1;    relay_conn far_4_4352_1_a(.in(far_4_4352_0[0]), .out(far_4_4352_1[0]));    relay_conn far_4_4352_1_b(.in(far_4_4352_0[1]), .out(far_4_4352_1[1]));
    assign layer_4[272] = far_4_4352_1[1] & ~far_4_4352_1[0]; 
    wire [1:0] far_4_4353_0;    relay_conn far_4_4353_0_a(.in(layer_3[119]), .out(far_4_4353_0[0]));    relay_conn far_4_4353_0_b(.in(layer_3[175]), .out(far_4_4353_0[1]));
    assign layer_4[273] = ~far_4_4353_0[0]; 
    wire [1:0] far_4_4354_0;    relay_conn far_4_4354_0_a(.in(layer_3[124]), .out(far_4_4354_0[0]));    relay_conn far_4_4354_0_b(.in(layer_3[72]), .out(far_4_4354_0[1]));
    assign layer_4[274] = ~(far_4_4354_0[0] | far_4_4354_0[1]); 
    assign layer_4[275] = layer_3[778] & ~layer_3[756]; 
    assign layer_4[276] = layer_3[533] | layer_3[514]; 
    assign layer_4[277] = layer_3[100] & ~layer_3[73]; 
    assign layer_4[278] = layer_3[340] & ~layer_3[323]; 
    wire [1:0] far_4_4359_0;    relay_conn far_4_4359_0_a(.in(layer_3[161]), .out(far_4_4359_0[0]));    relay_conn far_4_4359_0_b(.in(layer_3[58]), .out(far_4_4359_0[1]));
    wire [1:0] far_4_4359_1;    relay_conn far_4_4359_1_a(.in(far_4_4359_0[0]), .out(far_4_4359_1[0]));    relay_conn far_4_4359_1_b(.in(far_4_4359_0[1]), .out(far_4_4359_1[1]));
    wire [1:0] far_4_4359_2;    relay_conn far_4_4359_2_a(.in(far_4_4359_1[0]), .out(far_4_4359_2[0]));    relay_conn far_4_4359_2_b(.in(far_4_4359_1[1]), .out(far_4_4359_2[1]));
    assign layer_4[279] = ~far_4_4359_2[0] | (far_4_4359_2[0] & far_4_4359_2[1]); 
    wire [1:0] far_4_4360_0;    relay_conn far_4_4360_0_a(.in(layer_3[323]), .out(far_4_4360_0[0]));    relay_conn far_4_4360_0_b(.in(layer_3[397]), .out(far_4_4360_0[1]));
    wire [1:0] far_4_4360_1;    relay_conn far_4_4360_1_a(.in(far_4_4360_0[0]), .out(far_4_4360_1[0]));    relay_conn far_4_4360_1_b(.in(far_4_4360_0[1]), .out(far_4_4360_1[1]));
    assign layer_4[280] = far_4_4360_1[0] & far_4_4360_1[1]; 
    wire [1:0] far_4_4361_0;    relay_conn far_4_4361_0_a(.in(layer_3[761]), .out(far_4_4361_0[0]));    relay_conn far_4_4361_0_b(.in(layer_3[846]), .out(far_4_4361_0[1]));
    wire [1:0] far_4_4361_1;    relay_conn far_4_4361_1_a(.in(far_4_4361_0[0]), .out(far_4_4361_1[0]));    relay_conn far_4_4361_1_b(.in(far_4_4361_0[1]), .out(far_4_4361_1[1]));
    assign layer_4[281] = far_4_4361_1[0]; 
    assign layer_4[282] = ~layer_3[318] | (layer_3[334] & layer_3[318]); 
    wire [1:0] far_4_4363_0;    relay_conn far_4_4363_0_a(.in(layer_3[66]), .out(far_4_4363_0[0]));    relay_conn far_4_4363_0_b(.in(layer_3[125]), .out(far_4_4363_0[1]));
    assign layer_4[283] = far_4_4363_0[0] | far_4_4363_0[1]; 
    wire [1:0] far_4_4364_0;    relay_conn far_4_4364_0_a(.in(layer_3[370]), .out(far_4_4364_0[0]));    relay_conn far_4_4364_0_b(.in(layer_3[473]), .out(far_4_4364_0[1]));
    wire [1:0] far_4_4364_1;    relay_conn far_4_4364_1_a(.in(far_4_4364_0[0]), .out(far_4_4364_1[0]));    relay_conn far_4_4364_1_b(.in(far_4_4364_0[1]), .out(far_4_4364_1[1]));
    wire [1:0] far_4_4364_2;    relay_conn far_4_4364_2_a(.in(far_4_4364_1[0]), .out(far_4_4364_2[0]));    relay_conn far_4_4364_2_b(.in(far_4_4364_1[1]), .out(far_4_4364_2[1]));
    assign layer_4[284] = far_4_4364_2[0] & far_4_4364_2[1]; 
    wire [1:0] far_4_4365_0;    relay_conn far_4_4365_0_a(.in(layer_3[93]), .out(far_4_4365_0[0]));    relay_conn far_4_4365_0_b(.in(layer_3[147]), .out(far_4_4365_0[1]));
    assign layer_4[285] = far_4_4365_0[0] | far_4_4365_0[1]; 
    wire [1:0] far_4_4366_0;    relay_conn far_4_4366_0_a(.in(layer_3[274]), .out(far_4_4366_0[0]));    relay_conn far_4_4366_0_b(.in(layer_3[358]), .out(far_4_4366_0[1]));
    wire [1:0] far_4_4366_1;    relay_conn far_4_4366_1_a(.in(far_4_4366_0[0]), .out(far_4_4366_1[0]));    relay_conn far_4_4366_1_b(.in(far_4_4366_0[1]), .out(far_4_4366_1[1]));
    assign layer_4[286] = ~far_4_4366_1[0] | (far_4_4366_1[0] & far_4_4366_1[1]); 
    wire [1:0] far_4_4367_0;    relay_conn far_4_4367_0_a(.in(layer_3[337]), .out(far_4_4367_0[0]));    relay_conn far_4_4367_0_b(.in(layer_3[388]), .out(far_4_4367_0[1]));
    assign layer_4[287] = ~far_4_4367_0[1]; 
    wire [1:0] far_4_4368_0;    relay_conn far_4_4368_0_a(.in(layer_3[807]), .out(far_4_4368_0[0]));    relay_conn far_4_4368_0_b(.in(layer_3[879]), .out(far_4_4368_0[1]));
    wire [1:0] far_4_4368_1;    relay_conn far_4_4368_1_a(.in(far_4_4368_0[0]), .out(far_4_4368_1[0]));    relay_conn far_4_4368_1_b(.in(far_4_4368_0[1]), .out(far_4_4368_1[1]));
    assign layer_4[288] = far_4_4368_1[0] ^ far_4_4368_1[1]; 
    wire [1:0] far_4_4369_0;    relay_conn far_4_4369_0_a(.in(layer_3[534]), .out(far_4_4369_0[0]));    relay_conn far_4_4369_0_b(.in(layer_3[605]), .out(far_4_4369_0[1]));
    wire [1:0] far_4_4369_1;    relay_conn far_4_4369_1_a(.in(far_4_4369_0[0]), .out(far_4_4369_1[0]));    relay_conn far_4_4369_1_b(.in(far_4_4369_0[1]), .out(far_4_4369_1[1]));
    assign layer_4[289] = far_4_4369_1[0] | far_4_4369_1[1]; 
    wire [1:0] far_4_4370_0;    relay_conn far_4_4370_0_a(.in(layer_3[438]), .out(far_4_4370_0[0]));    relay_conn far_4_4370_0_b(.in(layer_3[332]), .out(far_4_4370_0[1]));
    wire [1:0] far_4_4370_1;    relay_conn far_4_4370_1_a(.in(far_4_4370_0[0]), .out(far_4_4370_1[0]));    relay_conn far_4_4370_1_b(.in(far_4_4370_0[1]), .out(far_4_4370_1[1]));
    wire [1:0] far_4_4370_2;    relay_conn far_4_4370_2_a(.in(far_4_4370_1[0]), .out(far_4_4370_2[0]));    relay_conn far_4_4370_2_b(.in(far_4_4370_1[1]), .out(far_4_4370_2[1]));
    assign layer_4[290] = ~(far_4_4370_2[0] ^ far_4_4370_2[1]); 
    wire [1:0] far_4_4371_0;    relay_conn far_4_4371_0_a(.in(layer_3[958]), .out(far_4_4371_0[0]));    relay_conn far_4_4371_0_b(.in(layer_3[889]), .out(far_4_4371_0[1]));
    wire [1:0] far_4_4371_1;    relay_conn far_4_4371_1_a(.in(far_4_4371_0[0]), .out(far_4_4371_1[0]));    relay_conn far_4_4371_1_b(.in(far_4_4371_0[1]), .out(far_4_4371_1[1]));
    assign layer_4[291] = ~far_4_4371_1[0]; 
    wire [1:0] far_4_4372_0;    relay_conn far_4_4372_0_a(.in(layer_3[252]), .out(far_4_4372_0[0]));    relay_conn far_4_4372_0_b(.in(layer_3[197]), .out(far_4_4372_0[1]));
    assign layer_4[292] = ~far_4_4372_0[0] | (far_4_4372_0[0] & far_4_4372_0[1]); 
    assign layer_4[293] = layer_3[52] & ~layer_3[61]; 
    wire [1:0] far_4_4374_0;    relay_conn far_4_4374_0_a(.in(layer_3[266]), .out(far_4_4374_0[0]));    relay_conn far_4_4374_0_b(.in(layer_3[372]), .out(far_4_4374_0[1]));
    wire [1:0] far_4_4374_1;    relay_conn far_4_4374_1_a(.in(far_4_4374_0[0]), .out(far_4_4374_1[0]));    relay_conn far_4_4374_1_b(.in(far_4_4374_0[1]), .out(far_4_4374_1[1]));
    wire [1:0] far_4_4374_2;    relay_conn far_4_4374_2_a(.in(far_4_4374_1[0]), .out(far_4_4374_2[0]));    relay_conn far_4_4374_2_b(.in(far_4_4374_1[1]), .out(far_4_4374_2[1]));
    assign layer_4[294] = far_4_4374_2[0]; 
    assign layer_4[295] = layer_3[362] | layer_3[337]; 
    wire [1:0] far_4_4376_0;    relay_conn far_4_4376_0_a(.in(layer_3[47]), .out(far_4_4376_0[0]));    relay_conn far_4_4376_0_b(.in(layer_3[164]), .out(far_4_4376_0[1]));
    wire [1:0] far_4_4376_1;    relay_conn far_4_4376_1_a(.in(far_4_4376_0[0]), .out(far_4_4376_1[0]));    relay_conn far_4_4376_1_b(.in(far_4_4376_0[1]), .out(far_4_4376_1[1]));
    wire [1:0] far_4_4376_2;    relay_conn far_4_4376_2_a(.in(far_4_4376_1[0]), .out(far_4_4376_2[0]));    relay_conn far_4_4376_2_b(.in(far_4_4376_1[1]), .out(far_4_4376_2[1]));
    assign layer_4[296] = far_4_4376_2[0] | far_4_4376_2[1]; 
    wire [1:0] far_4_4377_0;    relay_conn far_4_4377_0_a(.in(layer_3[967]), .out(far_4_4377_0[0]));    relay_conn far_4_4377_0_b(.in(layer_3[846]), .out(far_4_4377_0[1]));
    wire [1:0] far_4_4377_1;    relay_conn far_4_4377_1_a(.in(far_4_4377_0[0]), .out(far_4_4377_1[0]));    relay_conn far_4_4377_1_b(.in(far_4_4377_0[1]), .out(far_4_4377_1[1]));
    wire [1:0] far_4_4377_2;    relay_conn far_4_4377_2_a(.in(far_4_4377_1[0]), .out(far_4_4377_2[0]));    relay_conn far_4_4377_2_b(.in(far_4_4377_1[1]), .out(far_4_4377_2[1]));
    assign layer_4[297] = ~far_4_4377_2[0] | (far_4_4377_2[0] & far_4_4377_2[1]); 
    assign layer_4[298] = ~layer_3[352] | (layer_3[352] & layer_3[323]); 
    wire [1:0] far_4_4379_0;    relay_conn far_4_4379_0_a(.in(layer_3[279]), .out(far_4_4379_0[0]));    relay_conn far_4_4379_0_b(.in(layer_3[178]), .out(far_4_4379_0[1]));
    wire [1:0] far_4_4379_1;    relay_conn far_4_4379_1_a(.in(far_4_4379_0[0]), .out(far_4_4379_1[0]));    relay_conn far_4_4379_1_b(.in(far_4_4379_0[1]), .out(far_4_4379_1[1]));
    wire [1:0] far_4_4379_2;    relay_conn far_4_4379_2_a(.in(far_4_4379_1[0]), .out(far_4_4379_2[0]));    relay_conn far_4_4379_2_b(.in(far_4_4379_1[1]), .out(far_4_4379_2[1]));
    assign layer_4[299] = far_4_4379_2[0] & far_4_4379_2[1]; 
    wire [1:0] far_4_4380_0;    relay_conn far_4_4380_0_a(.in(layer_3[575]), .out(far_4_4380_0[0]));    relay_conn far_4_4380_0_b(.in(layer_3[454]), .out(far_4_4380_0[1]));
    wire [1:0] far_4_4380_1;    relay_conn far_4_4380_1_a(.in(far_4_4380_0[0]), .out(far_4_4380_1[0]));    relay_conn far_4_4380_1_b(.in(far_4_4380_0[1]), .out(far_4_4380_1[1]));
    wire [1:0] far_4_4380_2;    relay_conn far_4_4380_2_a(.in(far_4_4380_1[0]), .out(far_4_4380_2[0]));    relay_conn far_4_4380_2_b(.in(far_4_4380_1[1]), .out(far_4_4380_2[1]));
    assign layer_4[300] = far_4_4380_2[1]; 
    wire [1:0] far_4_4381_0;    relay_conn far_4_4381_0_a(.in(layer_3[860]), .out(far_4_4381_0[0]));    relay_conn far_4_4381_0_b(.in(layer_3[791]), .out(far_4_4381_0[1]));
    wire [1:0] far_4_4381_1;    relay_conn far_4_4381_1_a(.in(far_4_4381_0[0]), .out(far_4_4381_1[0]));    relay_conn far_4_4381_1_b(.in(far_4_4381_0[1]), .out(far_4_4381_1[1]));
    assign layer_4[301] = ~far_4_4381_1[0]; 
    wire [1:0] far_4_4382_0;    relay_conn far_4_4382_0_a(.in(layer_3[629]), .out(far_4_4382_0[0]));    relay_conn far_4_4382_0_b(.in(layer_3[582]), .out(far_4_4382_0[1]));
    assign layer_4[302] = far_4_4382_0[0] & ~far_4_4382_0[1]; 
    assign layer_4[303] = ~(layer_3[497] & layer_3[467]); 
    wire [1:0] far_4_4384_0;    relay_conn far_4_4384_0_a(.in(layer_3[880]), .out(far_4_4384_0[0]));    relay_conn far_4_4384_0_b(.in(layer_3[923]), .out(far_4_4384_0[1]));
    assign layer_4[304] = ~far_4_4384_0[0]; 
    wire [1:0] far_4_4385_0;    relay_conn far_4_4385_0_a(.in(layer_3[67]), .out(far_4_4385_0[0]));    relay_conn far_4_4385_0_b(.in(layer_3[31]), .out(far_4_4385_0[1]));
    assign layer_4[305] = ~far_4_4385_0[1] | (far_4_4385_0[0] & far_4_4385_0[1]); 
    wire [1:0] far_4_4386_0;    relay_conn far_4_4386_0_a(.in(layer_3[770]), .out(far_4_4386_0[0]));    relay_conn far_4_4386_0_b(.in(layer_3[846]), .out(far_4_4386_0[1]));
    wire [1:0] far_4_4386_1;    relay_conn far_4_4386_1_a(.in(far_4_4386_0[0]), .out(far_4_4386_1[0]));    relay_conn far_4_4386_1_b(.in(far_4_4386_0[1]), .out(far_4_4386_1[1]));
    assign layer_4[306] = far_4_4386_1[1]; 
    wire [1:0] far_4_4387_0;    relay_conn far_4_4387_0_a(.in(layer_3[368]), .out(far_4_4387_0[0]));    relay_conn far_4_4387_0_b(.in(layer_3[436]), .out(far_4_4387_0[1]));
    wire [1:0] far_4_4387_1;    relay_conn far_4_4387_1_a(.in(far_4_4387_0[0]), .out(far_4_4387_1[0]));    relay_conn far_4_4387_1_b(.in(far_4_4387_0[1]), .out(far_4_4387_1[1]));
    assign layer_4[307] = far_4_4387_1[0] & ~far_4_4387_1[1]; 
    wire [1:0] far_4_4388_0;    relay_conn far_4_4388_0_a(.in(layer_3[125]), .out(far_4_4388_0[0]));    relay_conn far_4_4388_0_b(.in(layer_3[36]), .out(far_4_4388_0[1]));
    wire [1:0] far_4_4388_1;    relay_conn far_4_4388_1_a(.in(far_4_4388_0[0]), .out(far_4_4388_1[0]));    relay_conn far_4_4388_1_b(.in(far_4_4388_0[1]), .out(far_4_4388_1[1]));
    assign layer_4[308] = ~far_4_4388_1[1] | (far_4_4388_1[0] & far_4_4388_1[1]); 
    wire [1:0] far_4_4389_0;    relay_conn far_4_4389_0_a(.in(layer_3[901]), .out(far_4_4389_0[0]));    relay_conn far_4_4389_0_b(.in(layer_3[855]), .out(far_4_4389_0[1]));
    assign layer_4[309] = ~far_4_4389_0[0]; 
    assign layer_4[310] = ~layer_3[400] | (layer_3[372] & layer_3[400]); 
    wire [1:0] far_4_4391_0;    relay_conn far_4_4391_0_a(.in(layer_3[882]), .out(far_4_4391_0[0]));    relay_conn far_4_4391_0_b(.in(layer_3[916]), .out(far_4_4391_0[1]));
    assign layer_4[311] = far_4_4391_0[0]; 
    wire [1:0] far_4_4392_0;    relay_conn far_4_4392_0_a(.in(layer_3[718]), .out(far_4_4392_0[0]));    relay_conn far_4_4392_0_b(.in(layer_3[682]), .out(far_4_4392_0[1]));
    assign layer_4[312] = ~(far_4_4392_0[0] | far_4_4392_0[1]); 
    wire [1:0] far_4_4393_0;    relay_conn far_4_4393_0_a(.in(layer_3[697]), .out(far_4_4393_0[0]));    relay_conn far_4_4393_0_b(.in(layer_3[572]), .out(far_4_4393_0[1]));
    wire [1:0] far_4_4393_1;    relay_conn far_4_4393_1_a(.in(far_4_4393_0[0]), .out(far_4_4393_1[0]));    relay_conn far_4_4393_1_b(.in(far_4_4393_0[1]), .out(far_4_4393_1[1]));
    wire [1:0] far_4_4393_2;    relay_conn far_4_4393_2_a(.in(far_4_4393_1[0]), .out(far_4_4393_2[0]));    relay_conn far_4_4393_2_b(.in(far_4_4393_1[1]), .out(far_4_4393_2[1]));
    assign layer_4[313] = far_4_4393_2[0] | far_4_4393_2[1]; 
    wire [1:0] far_4_4394_0;    relay_conn far_4_4394_0_a(.in(layer_3[226]), .out(far_4_4394_0[0]));    relay_conn far_4_4394_0_b(.in(layer_3[124]), .out(far_4_4394_0[1]));
    wire [1:0] far_4_4394_1;    relay_conn far_4_4394_1_a(.in(far_4_4394_0[0]), .out(far_4_4394_1[0]));    relay_conn far_4_4394_1_b(.in(far_4_4394_0[1]), .out(far_4_4394_1[1]));
    wire [1:0] far_4_4394_2;    relay_conn far_4_4394_2_a(.in(far_4_4394_1[0]), .out(far_4_4394_2[0]));    relay_conn far_4_4394_2_b(.in(far_4_4394_1[1]), .out(far_4_4394_2[1]));
    assign layer_4[314] = far_4_4394_2[0] | far_4_4394_2[1]; 
    wire [1:0] far_4_4395_0;    relay_conn far_4_4395_0_a(.in(layer_3[459]), .out(far_4_4395_0[0]));    relay_conn far_4_4395_0_b(.in(layer_3[544]), .out(far_4_4395_0[1]));
    wire [1:0] far_4_4395_1;    relay_conn far_4_4395_1_a(.in(far_4_4395_0[0]), .out(far_4_4395_1[0]));    relay_conn far_4_4395_1_b(.in(far_4_4395_0[1]), .out(far_4_4395_1[1]));
    assign layer_4[315] = ~(far_4_4395_1[0] & far_4_4395_1[1]); 
    wire [1:0] far_4_4396_0;    relay_conn far_4_4396_0_a(.in(layer_3[64]), .out(far_4_4396_0[0]));    relay_conn far_4_4396_0_b(.in(layer_3[0]), .out(far_4_4396_0[1]));
    wire [1:0] far_4_4396_1;    relay_conn far_4_4396_1_a(.in(far_4_4396_0[0]), .out(far_4_4396_1[0]));    relay_conn far_4_4396_1_b(.in(far_4_4396_0[1]), .out(far_4_4396_1[1]));
    assign layer_4[316] = far_4_4396_1[0] | far_4_4396_1[1]; 
    wire [1:0] far_4_4397_0;    relay_conn far_4_4397_0_a(.in(layer_3[251]), .out(far_4_4397_0[0]));    relay_conn far_4_4397_0_b(.in(layer_3[356]), .out(far_4_4397_0[1]));
    wire [1:0] far_4_4397_1;    relay_conn far_4_4397_1_a(.in(far_4_4397_0[0]), .out(far_4_4397_1[0]));    relay_conn far_4_4397_1_b(.in(far_4_4397_0[1]), .out(far_4_4397_1[1]));
    wire [1:0] far_4_4397_2;    relay_conn far_4_4397_2_a(.in(far_4_4397_1[0]), .out(far_4_4397_2[0]));    relay_conn far_4_4397_2_b(.in(far_4_4397_1[1]), .out(far_4_4397_2[1]));
    assign layer_4[317] = far_4_4397_2[0]; 
    assign layer_4[318] = ~layer_3[364] | (layer_3[364] & layer_3[363]); 
    wire [1:0] far_4_4399_0;    relay_conn far_4_4399_0_a(.in(layer_3[134]), .out(far_4_4399_0[0]));    relay_conn far_4_4399_0_b(.in(layer_3[238]), .out(far_4_4399_0[1]));
    wire [1:0] far_4_4399_1;    relay_conn far_4_4399_1_a(.in(far_4_4399_0[0]), .out(far_4_4399_1[0]));    relay_conn far_4_4399_1_b(.in(far_4_4399_0[1]), .out(far_4_4399_1[1]));
    wire [1:0] far_4_4399_2;    relay_conn far_4_4399_2_a(.in(far_4_4399_1[0]), .out(far_4_4399_2[0]));    relay_conn far_4_4399_2_b(.in(far_4_4399_1[1]), .out(far_4_4399_2[1]));
    assign layer_4[319] = far_4_4399_2[0] | far_4_4399_2[1]; 
    wire [1:0] far_4_4400_0;    relay_conn far_4_4400_0_a(.in(layer_3[692]), .out(far_4_4400_0[0]));    relay_conn far_4_4400_0_b(.in(layer_3[605]), .out(far_4_4400_0[1]));
    wire [1:0] far_4_4400_1;    relay_conn far_4_4400_1_a(.in(far_4_4400_0[0]), .out(far_4_4400_1[0]));    relay_conn far_4_4400_1_b(.in(far_4_4400_0[1]), .out(far_4_4400_1[1]));
    assign layer_4[320] = ~(far_4_4400_1[0] ^ far_4_4400_1[1]); 
    wire [1:0] far_4_4401_0;    relay_conn far_4_4401_0_a(.in(layer_3[92]), .out(far_4_4401_0[0]));    relay_conn far_4_4401_0_b(.in(layer_3[2]), .out(far_4_4401_0[1]));
    wire [1:0] far_4_4401_1;    relay_conn far_4_4401_1_a(.in(far_4_4401_0[0]), .out(far_4_4401_1[0]));    relay_conn far_4_4401_1_b(.in(far_4_4401_0[1]), .out(far_4_4401_1[1]));
    assign layer_4[321] = far_4_4401_1[0]; 
    wire [1:0] far_4_4402_0;    relay_conn far_4_4402_0_a(.in(layer_3[353]), .out(far_4_4402_0[0]));    relay_conn far_4_4402_0_b(.in(layer_3[305]), .out(far_4_4402_0[1]));
    assign layer_4[322] = far_4_4402_0[1]; 
    wire [1:0] far_4_4403_0;    relay_conn far_4_4403_0_a(.in(layer_3[335]), .out(far_4_4403_0[0]));    relay_conn far_4_4403_0_b(.in(layer_3[426]), .out(far_4_4403_0[1]));
    wire [1:0] far_4_4403_1;    relay_conn far_4_4403_1_a(.in(far_4_4403_0[0]), .out(far_4_4403_1[0]));    relay_conn far_4_4403_1_b(.in(far_4_4403_0[1]), .out(far_4_4403_1[1]));
    assign layer_4[323] = far_4_4403_1[1]; 
    wire [1:0] far_4_4404_0;    relay_conn far_4_4404_0_a(.in(layer_3[570]), .out(far_4_4404_0[0]));    relay_conn far_4_4404_0_b(.in(layer_3[698]), .out(far_4_4404_0[1]));
    wire [1:0] far_4_4404_1;    relay_conn far_4_4404_1_a(.in(far_4_4404_0[0]), .out(far_4_4404_1[0]));    relay_conn far_4_4404_1_b(.in(far_4_4404_0[1]), .out(far_4_4404_1[1]));
    wire [1:0] far_4_4404_2;    relay_conn far_4_4404_2_a(.in(far_4_4404_1[0]), .out(far_4_4404_2[0]));    relay_conn far_4_4404_2_b(.in(far_4_4404_1[1]), .out(far_4_4404_2[1]));
    wire [1:0] far_4_4404_3;    relay_conn far_4_4404_3_a(.in(far_4_4404_2[0]), .out(far_4_4404_3[0]));    relay_conn far_4_4404_3_b(.in(far_4_4404_2[1]), .out(far_4_4404_3[1]));
    assign layer_4[324] = ~far_4_4404_3[0]; 
    wire [1:0] far_4_4405_0;    relay_conn far_4_4405_0_a(.in(layer_3[266]), .out(far_4_4405_0[0]));    relay_conn far_4_4405_0_b(.in(layer_3[352]), .out(far_4_4405_0[1]));
    wire [1:0] far_4_4405_1;    relay_conn far_4_4405_1_a(.in(far_4_4405_0[0]), .out(far_4_4405_1[0]));    relay_conn far_4_4405_1_b(.in(far_4_4405_0[1]), .out(far_4_4405_1[1]));
    assign layer_4[325] = far_4_4405_1[1] & ~far_4_4405_1[0]; 
    wire [1:0] far_4_4406_0;    relay_conn far_4_4406_0_a(.in(layer_3[576]), .out(far_4_4406_0[0]));    relay_conn far_4_4406_0_b(.in(layer_3[626]), .out(far_4_4406_0[1]));
    assign layer_4[326] = far_4_4406_0[1]; 
    assign layer_4[327] = ~(layer_3[391] & layer_3[409]); 
    wire [1:0] far_4_4408_0;    relay_conn far_4_4408_0_a(.in(layer_3[609]), .out(far_4_4408_0[0]));    relay_conn far_4_4408_0_b(.in(layer_3[553]), .out(far_4_4408_0[1]));
    assign layer_4[328] = ~far_4_4408_0[0]; 
    wire [1:0] far_4_4409_0;    relay_conn far_4_4409_0_a(.in(layer_3[784]), .out(far_4_4409_0[0]));    relay_conn far_4_4409_0_b(.in(layer_3[674]), .out(far_4_4409_0[1]));
    wire [1:0] far_4_4409_1;    relay_conn far_4_4409_1_a(.in(far_4_4409_0[0]), .out(far_4_4409_1[0]));    relay_conn far_4_4409_1_b(.in(far_4_4409_0[1]), .out(far_4_4409_1[1]));
    wire [1:0] far_4_4409_2;    relay_conn far_4_4409_2_a(.in(far_4_4409_1[0]), .out(far_4_4409_2[0]));    relay_conn far_4_4409_2_b(.in(far_4_4409_1[1]), .out(far_4_4409_2[1]));
    assign layer_4[329] = ~(far_4_4409_2[0] & far_4_4409_2[1]); 
    assign layer_4[330] = layer_3[157]; 
    assign layer_4[331] = ~layer_3[10]; 
    wire [1:0] far_4_4412_0;    relay_conn far_4_4412_0_a(.in(layer_3[398]), .out(far_4_4412_0[0]));    relay_conn far_4_4412_0_b(.in(layer_3[459]), .out(far_4_4412_0[1]));
    assign layer_4[332] = far_4_4412_0[0] & far_4_4412_0[1]; 
    wire [1:0] far_4_4413_0;    relay_conn far_4_4413_0_a(.in(layer_3[964]), .out(far_4_4413_0[0]));    relay_conn far_4_4413_0_b(.in(layer_3[882]), .out(far_4_4413_0[1]));
    wire [1:0] far_4_4413_1;    relay_conn far_4_4413_1_a(.in(far_4_4413_0[0]), .out(far_4_4413_1[0]));    relay_conn far_4_4413_1_b(.in(far_4_4413_0[1]), .out(far_4_4413_1[1]));
    assign layer_4[333] = ~far_4_4413_1[1]; 
    wire [1:0] far_4_4414_0;    relay_conn far_4_4414_0_a(.in(layer_3[102]), .out(far_4_4414_0[0]));    relay_conn far_4_4414_0_b(.in(layer_3[58]), .out(far_4_4414_0[1]));
    assign layer_4[334] = far_4_4414_0[0]; 
    wire [1:0] far_4_4415_0;    relay_conn far_4_4415_0_a(.in(layer_3[860]), .out(far_4_4415_0[0]));    relay_conn far_4_4415_0_b(.in(layer_3[801]), .out(far_4_4415_0[1]));
    assign layer_4[335] = far_4_4415_0[0] | far_4_4415_0[1]; 
    wire [1:0] far_4_4416_0;    relay_conn far_4_4416_0_a(.in(layer_3[100]), .out(far_4_4416_0[0]));    relay_conn far_4_4416_0_b(.in(layer_3[164]), .out(far_4_4416_0[1]));
    wire [1:0] far_4_4416_1;    relay_conn far_4_4416_1_a(.in(far_4_4416_0[0]), .out(far_4_4416_1[0]));    relay_conn far_4_4416_1_b(.in(far_4_4416_0[1]), .out(far_4_4416_1[1]));
    assign layer_4[336] = far_4_4416_1[0] & ~far_4_4416_1[1]; 
    wire [1:0] far_4_4417_0;    relay_conn far_4_4417_0_a(.in(layer_3[878]), .out(far_4_4417_0[0]));    relay_conn far_4_4417_0_b(.in(layer_3[834]), .out(far_4_4417_0[1]));
    assign layer_4[337] = ~far_4_4417_0[1]; 
    wire [1:0] far_4_4418_0;    relay_conn far_4_4418_0_a(.in(layer_3[353]), .out(far_4_4418_0[0]));    relay_conn far_4_4418_0_b(.in(layer_3[473]), .out(far_4_4418_0[1]));
    wire [1:0] far_4_4418_1;    relay_conn far_4_4418_1_a(.in(far_4_4418_0[0]), .out(far_4_4418_1[0]));    relay_conn far_4_4418_1_b(.in(far_4_4418_0[1]), .out(far_4_4418_1[1]));
    wire [1:0] far_4_4418_2;    relay_conn far_4_4418_2_a(.in(far_4_4418_1[0]), .out(far_4_4418_2[0]));    relay_conn far_4_4418_2_b(.in(far_4_4418_1[1]), .out(far_4_4418_2[1]));
    assign layer_4[338] = ~far_4_4418_2[0]; 
    wire [1:0] far_4_4419_0;    relay_conn far_4_4419_0_a(.in(layer_3[669]), .out(far_4_4419_0[0]));    relay_conn far_4_4419_0_b(.in(layer_3[633]), .out(far_4_4419_0[1]));
    assign layer_4[339] = far_4_4419_0[0] | far_4_4419_0[1]; 
    wire [1:0] far_4_4420_0;    relay_conn far_4_4420_0_a(.in(layer_3[143]), .out(far_4_4420_0[0]));    relay_conn far_4_4420_0_b(.in(layer_3[56]), .out(far_4_4420_0[1]));
    wire [1:0] far_4_4420_1;    relay_conn far_4_4420_1_a(.in(far_4_4420_0[0]), .out(far_4_4420_1[0]));    relay_conn far_4_4420_1_b(.in(far_4_4420_0[1]), .out(far_4_4420_1[1]));
    assign layer_4[340] = far_4_4420_1[0]; 
    assign layer_4[341] = ~layer_3[459]; 
    assign layer_4[342] = layer_3[1018]; 
    wire [1:0] far_4_4423_0;    relay_conn far_4_4423_0_a(.in(layer_3[112]), .out(far_4_4423_0[0]));    relay_conn far_4_4423_0_b(.in(layer_3[154]), .out(far_4_4423_0[1]));
    assign layer_4[343] = far_4_4423_0[0] & ~far_4_4423_0[1]; 
    assign layer_4[344] = ~(layer_3[642] ^ layer_3[634]); 
    assign layer_4[345] = layer_3[314] | layer_3[332]; 
    assign layer_4[346] = layer_3[936] & ~layer_3[964]; 
    wire [1:0] far_4_4427_0;    relay_conn far_4_4427_0_a(.in(layer_3[834]), .out(far_4_4427_0[0]));    relay_conn far_4_4427_0_b(.in(layer_3[898]), .out(far_4_4427_0[1]));
    wire [1:0] far_4_4427_1;    relay_conn far_4_4427_1_a(.in(far_4_4427_0[0]), .out(far_4_4427_1[0]));    relay_conn far_4_4427_1_b(.in(far_4_4427_0[1]), .out(far_4_4427_1[1]));
    assign layer_4[347] = far_4_4427_1[0]; 
    wire [1:0] far_4_4428_0;    relay_conn far_4_4428_0_a(.in(layer_3[715]), .out(far_4_4428_0[0]));    relay_conn far_4_4428_0_b(.in(layer_3[653]), .out(far_4_4428_0[1]));
    assign layer_4[348] = ~far_4_4428_0[0] | (far_4_4428_0[0] & far_4_4428_0[1]); 
    wire [1:0] far_4_4429_0;    relay_conn far_4_4429_0_a(.in(layer_3[279]), .out(far_4_4429_0[0]));    relay_conn far_4_4429_0_b(.in(layer_3[402]), .out(far_4_4429_0[1]));
    wire [1:0] far_4_4429_1;    relay_conn far_4_4429_1_a(.in(far_4_4429_0[0]), .out(far_4_4429_1[0]));    relay_conn far_4_4429_1_b(.in(far_4_4429_0[1]), .out(far_4_4429_1[1]));
    wire [1:0] far_4_4429_2;    relay_conn far_4_4429_2_a(.in(far_4_4429_1[0]), .out(far_4_4429_2[0]));    relay_conn far_4_4429_2_b(.in(far_4_4429_1[1]), .out(far_4_4429_2[1]));
    assign layer_4[349] = far_4_4429_2[0] & far_4_4429_2[1]; 
    wire [1:0] far_4_4430_0;    relay_conn far_4_4430_0_a(.in(layer_3[318]), .out(far_4_4430_0[0]));    relay_conn far_4_4430_0_b(.in(layer_3[434]), .out(far_4_4430_0[1]));
    wire [1:0] far_4_4430_1;    relay_conn far_4_4430_1_a(.in(far_4_4430_0[0]), .out(far_4_4430_1[0]));    relay_conn far_4_4430_1_b(.in(far_4_4430_0[1]), .out(far_4_4430_1[1]));
    wire [1:0] far_4_4430_2;    relay_conn far_4_4430_2_a(.in(far_4_4430_1[0]), .out(far_4_4430_2[0]));    relay_conn far_4_4430_2_b(.in(far_4_4430_1[1]), .out(far_4_4430_2[1]));
    assign layer_4[350] = ~(far_4_4430_2[0] & far_4_4430_2[1]); 
    wire [1:0] far_4_4431_0;    relay_conn far_4_4431_0_a(.in(layer_3[605]), .out(far_4_4431_0[0]));    relay_conn far_4_4431_0_b(.in(layer_3[709]), .out(far_4_4431_0[1]));
    wire [1:0] far_4_4431_1;    relay_conn far_4_4431_1_a(.in(far_4_4431_0[0]), .out(far_4_4431_1[0]));    relay_conn far_4_4431_1_b(.in(far_4_4431_0[1]), .out(far_4_4431_1[1]));
    wire [1:0] far_4_4431_2;    relay_conn far_4_4431_2_a(.in(far_4_4431_1[0]), .out(far_4_4431_2[0]));    relay_conn far_4_4431_2_b(.in(far_4_4431_1[1]), .out(far_4_4431_2[1]));
    assign layer_4[351] = ~far_4_4431_2[0] | (far_4_4431_2[0] & far_4_4431_2[1]); 
    wire [1:0] far_4_4432_0;    relay_conn far_4_4432_0_a(.in(layer_3[991]), .out(far_4_4432_0[0]));    relay_conn far_4_4432_0_b(.in(layer_3[909]), .out(far_4_4432_0[1]));
    wire [1:0] far_4_4432_1;    relay_conn far_4_4432_1_a(.in(far_4_4432_0[0]), .out(far_4_4432_1[0]));    relay_conn far_4_4432_1_b(.in(far_4_4432_0[1]), .out(far_4_4432_1[1]));
    assign layer_4[352] = far_4_4432_1[1] & ~far_4_4432_1[0]; 
    wire [1:0] far_4_4433_0;    relay_conn far_4_4433_0_a(.in(layer_3[768]), .out(far_4_4433_0[0]));    relay_conn far_4_4433_0_b(.in(layer_3[672]), .out(far_4_4433_0[1]));
    wire [1:0] far_4_4433_1;    relay_conn far_4_4433_1_a(.in(far_4_4433_0[0]), .out(far_4_4433_1[0]));    relay_conn far_4_4433_1_b(.in(far_4_4433_0[1]), .out(far_4_4433_1[1]));
    wire [1:0] far_4_4433_2;    relay_conn far_4_4433_2_a(.in(far_4_4433_1[0]), .out(far_4_4433_2[0]));    relay_conn far_4_4433_2_b(.in(far_4_4433_1[1]), .out(far_4_4433_2[1]));
    assign layer_4[353] = ~far_4_4433_2[0] | (far_4_4433_2[0] & far_4_4433_2[1]); 
    wire [1:0] far_4_4434_0;    relay_conn far_4_4434_0_a(.in(layer_3[218]), .out(far_4_4434_0[0]));    relay_conn far_4_4434_0_b(.in(layer_3[94]), .out(far_4_4434_0[1]));
    wire [1:0] far_4_4434_1;    relay_conn far_4_4434_1_a(.in(far_4_4434_0[0]), .out(far_4_4434_1[0]));    relay_conn far_4_4434_1_b(.in(far_4_4434_0[1]), .out(far_4_4434_1[1]));
    wire [1:0] far_4_4434_2;    relay_conn far_4_4434_2_a(.in(far_4_4434_1[0]), .out(far_4_4434_2[0]));    relay_conn far_4_4434_2_b(.in(far_4_4434_1[1]), .out(far_4_4434_2[1]));
    assign layer_4[354] = ~far_4_4434_2[1] | (far_4_4434_2[0] & far_4_4434_2[1]); 
    wire [1:0] far_4_4435_0;    relay_conn far_4_4435_0_a(.in(layer_3[903]), .out(far_4_4435_0[0]));    relay_conn far_4_4435_0_b(.in(layer_3[991]), .out(far_4_4435_0[1]));
    wire [1:0] far_4_4435_1;    relay_conn far_4_4435_1_a(.in(far_4_4435_0[0]), .out(far_4_4435_1[0]));    relay_conn far_4_4435_1_b(.in(far_4_4435_0[1]), .out(far_4_4435_1[1]));
    assign layer_4[355] = far_4_4435_1[0] | far_4_4435_1[1]; 
    wire [1:0] far_4_4436_0;    relay_conn far_4_4436_0_a(.in(layer_3[707]), .out(far_4_4436_0[0]));    relay_conn far_4_4436_0_b(.in(layer_3[740]), .out(far_4_4436_0[1]));
    assign layer_4[356] = ~far_4_4436_0[1] | (far_4_4436_0[0] & far_4_4436_0[1]); 
    wire [1:0] far_4_4437_0;    relay_conn far_4_4437_0_a(.in(layer_3[116]), .out(far_4_4437_0[0]));    relay_conn far_4_4437_0_b(.in(layer_3[63]), .out(far_4_4437_0[1]));
    assign layer_4[357] = ~far_4_4437_0[1]; 
    wire [1:0] far_4_4438_0;    relay_conn far_4_4438_0_a(.in(layer_3[350]), .out(far_4_4438_0[0]));    relay_conn far_4_4438_0_b(.in(layer_3[285]), .out(far_4_4438_0[1]));
    wire [1:0] far_4_4438_1;    relay_conn far_4_4438_1_a(.in(far_4_4438_0[0]), .out(far_4_4438_1[0]));    relay_conn far_4_4438_1_b(.in(far_4_4438_0[1]), .out(far_4_4438_1[1]));
    assign layer_4[358] = far_4_4438_1[0] & far_4_4438_1[1]; 
    wire [1:0] far_4_4439_0;    relay_conn far_4_4439_0_a(.in(layer_3[416]), .out(far_4_4439_0[0]));    relay_conn far_4_4439_0_b(.in(layer_3[375]), .out(far_4_4439_0[1]));
    assign layer_4[359] = far_4_4439_0[1]; 
    wire [1:0] far_4_4440_0;    relay_conn far_4_4440_0_a(.in(layer_3[977]), .out(far_4_4440_0[0]));    relay_conn far_4_4440_0_b(.in(layer_3[896]), .out(far_4_4440_0[1]));
    wire [1:0] far_4_4440_1;    relay_conn far_4_4440_1_a(.in(far_4_4440_0[0]), .out(far_4_4440_1[0]));    relay_conn far_4_4440_1_b(.in(far_4_4440_0[1]), .out(far_4_4440_1[1]));
    assign layer_4[360] = ~(far_4_4440_1[0] | far_4_4440_1[1]); 
    wire [1:0] far_4_4441_0;    relay_conn far_4_4441_0_a(.in(layer_3[50]), .out(far_4_4441_0[0]));    relay_conn far_4_4441_0_b(.in(layer_3[1]), .out(far_4_4441_0[1]));
    assign layer_4[361] = ~far_4_4441_0[0]; 
    wire [1:0] far_4_4442_0;    relay_conn far_4_4442_0_a(.in(layer_3[368]), .out(far_4_4442_0[0]));    relay_conn far_4_4442_0_b(.in(layer_3[467]), .out(far_4_4442_0[1]));
    wire [1:0] far_4_4442_1;    relay_conn far_4_4442_1_a(.in(far_4_4442_0[0]), .out(far_4_4442_1[0]));    relay_conn far_4_4442_1_b(.in(far_4_4442_0[1]), .out(far_4_4442_1[1]));
    wire [1:0] far_4_4442_2;    relay_conn far_4_4442_2_a(.in(far_4_4442_1[0]), .out(far_4_4442_2[0]));    relay_conn far_4_4442_2_b(.in(far_4_4442_1[1]), .out(far_4_4442_2[1]));
    assign layer_4[362] = ~(far_4_4442_2[0] & far_4_4442_2[1]); 
    wire [1:0] far_4_4443_0;    relay_conn far_4_4443_0_a(.in(layer_3[149]), .out(far_4_4443_0[0]));    relay_conn far_4_4443_0_b(.in(layer_3[199]), .out(far_4_4443_0[1]));
    assign layer_4[363] = ~far_4_4443_0[0] | (far_4_4443_0[0] & far_4_4443_0[1]); 
    wire [1:0] far_4_4444_0;    relay_conn far_4_4444_0_a(.in(layer_3[63]), .out(far_4_4444_0[0]));    relay_conn far_4_4444_0_b(.in(layer_3[149]), .out(far_4_4444_0[1]));
    wire [1:0] far_4_4444_1;    relay_conn far_4_4444_1_a(.in(far_4_4444_0[0]), .out(far_4_4444_1[0]));    relay_conn far_4_4444_1_b(.in(far_4_4444_0[1]), .out(far_4_4444_1[1]));
    assign layer_4[364] = far_4_4444_1[0] & far_4_4444_1[1]; 
    wire [1:0] far_4_4445_0;    relay_conn far_4_4445_0_a(.in(layer_3[990]), .out(far_4_4445_0[0]));    relay_conn far_4_4445_0_b(.in(layer_3[886]), .out(far_4_4445_0[1]));
    wire [1:0] far_4_4445_1;    relay_conn far_4_4445_1_a(.in(far_4_4445_0[0]), .out(far_4_4445_1[0]));    relay_conn far_4_4445_1_b(.in(far_4_4445_0[1]), .out(far_4_4445_1[1]));
    wire [1:0] far_4_4445_2;    relay_conn far_4_4445_2_a(.in(far_4_4445_1[0]), .out(far_4_4445_2[0]));    relay_conn far_4_4445_2_b(.in(far_4_4445_1[1]), .out(far_4_4445_2[1]));
    assign layer_4[365] = far_4_4445_2[0] | far_4_4445_2[1]; 
    assign layer_4[366] = ~layer_3[512] | (layer_3[512] & layer_3[481]); 
    assign layer_4[367] = ~layer_3[950] | (layer_3[950] & layer_3[953]); 
    wire [1:0] far_4_4448_0;    relay_conn far_4_4448_0_a(.in(layer_3[949]), .out(far_4_4448_0[0]));    relay_conn far_4_4448_0_b(.in(layer_3[913]), .out(far_4_4448_0[1]));
    assign layer_4[368] = far_4_4448_0[0] | far_4_4448_0[1]; 
    wire [1:0] far_4_4449_0;    relay_conn far_4_4449_0_a(.in(layer_3[756]), .out(far_4_4449_0[0]));    relay_conn far_4_4449_0_b(.in(layer_3[831]), .out(far_4_4449_0[1]));
    wire [1:0] far_4_4449_1;    relay_conn far_4_4449_1_a(.in(far_4_4449_0[0]), .out(far_4_4449_1[0]));    relay_conn far_4_4449_1_b(.in(far_4_4449_0[1]), .out(far_4_4449_1[1]));
    assign layer_4[369] = ~(far_4_4449_1[0] & far_4_4449_1[1]); 
    wire [1:0] far_4_4450_0;    relay_conn far_4_4450_0_a(.in(layer_3[265]), .out(far_4_4450_0[0]));    relay_conn far_4_4450_0_b(.in(layer_3[160]), .out(far_4_4450_0[1]));
    wire [1:0] far_4_4450_1;    relay_conn far_4_4450_1_a(.in(far_4_4450_0[0]), .out(far_4_4450_1[0]));    relay_conn far_4_4450_1_b(.in(far_4_4450_0[1]), .out(far_4_4450_1[1]));
    wire [1:0] far_4_4450_2;    relay_conn far_4_4450_2_a(.in(far_4_4450_1[0]), .out(far_4_4450_2[0]));    relay_conn far_4_4450_2_b(.in(far_4_4450_1[1]), .out(far_4_4450_2[1]));
    assign layer_4[370] = ~far_4_4450_2[0] | (far_4_4450_2[0] & far_4_4450_2[1]); 
    assign layer_4[371] = layer_3[352] ^ layer_3[321]; 
    wire [1:0] far_4_4452_0;    relay_conn far_4_4452_0_a(.in(layer_3[511]), .out(far_4_4452_0[0]));    relay_conn far_4_4452_0_b(.in(layer_3[438]), .out(far_4_4452_0[1]));
    wire [1:0] far_4_4452_1;    relay_conn far_4_4452_1_a(.in(far_4_4452_0[0]), .out(far_4_4452_1[0]));    relay_conn far_4_4452_1_b(.in(far_4_4452_0[1]), .out(far_4_4452_1[1]));
    assign layer_4[372] = ~(far_4_4452_1[0] | far_4_4452_1[1]); 
    wire [1:0] far_4_4453_0;    relay_conn far_4_4453_0_a(.in(layer_3[199]), .out(far_4_4453_0[0]));    relay_conn far_4_4453_0_b(.in(layer_3[275]), .out(far_4_4453_0[1]));
    wire [1:0] far_4_4453_1;    relay_conn far_4_4453_1_a(.in(far_4_4453_0[0]), .out(far_4_4453_1[0]));    relay_conn far_4_4453_1_b(.in(far_4_4453_0[1]), .out(far_4_4453_1[1]));
    assign layer_4[373] = far_4_4453_1[0] ^ far_4_4453_1[1]; 
    assign layer_4[374] = ~layer_3[37]; 
    wire [1:0] far_4_4455_0;    relay_conn far_4_4455_0_a(.in(layer_3[581]), .out(far_4_4455_0[0]));    relay_conn far_4_4455_0_b(.in(layer_3[490]), .out(far_4_4455_0[1]));
    wire [1:0] far_4_4455_1;    relay_conn far_4_4455_1_a(.in(far_4_4455_0[0]), .out(far_4_4455_1[0]));    relay_conn far_4_4455_1_b(.in(far_4_4455_0[1]), .out(far_4_4455_1[1]));
    assign layer_4[375] = ~far_4_4455_1[1] | (far_4_4455_1[0] & far_4_4455_1[1]); 
    wire [1:0] far_4_4456_0;    relay_conn far_4_4456_0_a(.in(layer_3[207]), .out(far_4_4456_0[0]));    relay_conn far_4_4456_0_b(.in(layer_3[165]), .out(far_4_4456_0[1]));
    assign layer_4[376] = ~far_4_4456_0[0] | (far_4_4456_0[0] & far_4_4456_0[1]); 
    wire [1:0] far_4_4457_0;    relay_conn far_4_4457_0_a(.in(layer_3[104]), .out(far_4_4457_0[0]));    relay_conn far_4_4457_0_b(.in(layer_3[147]), .out(far_4_4457_0[1]));
    assign layer_4[377] = ~far_4_4457_0[0] | (far_4_4457_0[0] & far_4_4457_0[1]); 
    wire [1:0] far_4_4458_0;    relay_conn far_4_4458_0_a(.in(layer_3[467]), .out(far_4_4458_0[0]));    relay_conn far_4_4458_0_b(.in(layer_3[570]), .out(far_4_4458_0[1]));
    wire [1:0] far_4_4458_1;    relay_conn far_4_4458_1_a(.in(far_4_4458_0[0]), .out(far_4_4458_1[0]));    relay_conn far_4_4458_1_b(.in(far_4_4458_0[1]), .out(far_4_4458_1[1]));
    wire [1:0] far_4_4458_2;    relay_conn far_4_4458_2_a(.in(far_4_4458_1[0]), .out(far_4_4458_2[0]));    relay_conn far_4_4458_2_b(.in(far_4_4458_1[1]), .out(far_4_4458_2[1]));
    assign layer_4[378] = ~(far_4_4458_2[0] | far_4_4458_2[1]); 
    wire [1:0] far_4_4459_0;    relay_conn far_4_4459_0_a(.in(layer_3[524]), .out(far_4_4459_0[0]));    relay_conn far_4_4459_0_b(.in(layer_3[422]), .out(far_4_4459_0[1]));
    wire [1:0] far_4_4459_1;    relay_conn far_4_4459_1_a(.in(far_4_4459_0[0]), .out(far_4_4459_1[0]));    relay_conn far_4_4459_1_b(.in(far_4_4459_0[1]), .out(far_4_4459_1[1]));
    wire [1:0] far_4_4459_2;    relay_conn far_4_4459_2_a(.in(far_4_4459_1[0]), .out(far_4_4459_2[0]));    relay_conn far_4_4459_2_b(.in(far_4_4459_1[1]), .out(far_4_4459_2[1]));
    assign layer_4[379] = ~(far_4_4459_2[0] | far_4_4459_2[1]); 
    assign layer_4[380] = ~layer_3[909]; 
    assign layer_4[381] = ~layer_3[711] | (layer_3[685] & layer_3[711]); 
    wire [1:0] far_4_4462_0;    relay_conn far_4_4462_0_a(.in(layer_3[676]), .out(far_4_4462_0[0]));    relay_conn far_4_4462_0_b(.in(layer_3[565]), .out(far_4_4462_0[1]));
    wire [1:0] far_4_4462_1;    relay_conn far_4_4462_1_a(.in(far_4_4462_0[0]), .out(far_4_4462_1[0]));    relay_conn far_4_4462_1_b(.in(far_4_4462_0[1]), .out(far_4_4462_1[1]));
    wire [1:0] far_4_4462_2;    relay_conn far_4_4462_2_a(.in(far_4_4462_1[0]), .out(far_4_4462_2[0]));    relay_conn far_4_4462_2_b(.in(far_4_4462_1[1]), .out(far_4_4462_2[1]));
    assign layer_4[382] = ~far_4_4462_2[1] | (far_4_4462_2[0] & far_4_4462_2[1]); 
    assign layer_4[383] = ~layer_3[175] | (layer_3[175] & layer_3[196]); 
    wire [1:0] far_4_4464_0;    relay_conn far_4_4464_0_a(.in(layer_3[175]), .out(far_4_4464_0[0]));    relay_conn far_4_4464_0_b(.in(layer_3[279]), .out(far_4_4464_0[1]));
    wire [1:0] far_4_4464_1;    relay_conn far_4_4464_1_a(.in(far_4_4464_0[0]), .out(far_4_4464_1[0]));    relay_conn far_4_4464_1_b(.in(far_4_4464_0[1]), .out(far_4_4464_1[1]));
    wire [1:0] far_4_4464_2;    relay_conn far_4_4464_2_a(.in(far_4_4464_1[0]), .out(far_4_4464_2[0]));    relay_conn far_4_4464_2_b(.in(far_4_4464_1[1]), .out(far_4_4464_2[1]));
    assign layer_4[384] = ~far_4_4464_2[0] | (far_4_4464_2[0] & far_4_4464_2[1]); 
    wire [1:0] far_4_4465_0;    relay_conn far_4_4465_0_a(.in(layer_3[932]), .out(far_4_4465_0[0]));    relay_conn far_4_4465_0_b(.in(layer_3[848]), .out(far_4_4465_0[1]));
    wire [1:0] far_4_4465_1;    relay_conn far_4_4465_1_a(.in(far_4_4465_0[0]), .out(far_4_4465_1[0]));    relay_conn far_4_4465_1_b(.in(far_4_4465_0[1]), .out(far_4_4465_1[1]));
    assign layer_4[385] = far_4_4465_1[0] ^ far_4_4465_1[1]; 
    wire [1:0] far_4_4466_0;    relay_conn far_4_4466_0_a(.in(layer_3[507]), .out(far_4_4466_0[0]));    relay_conn far_4_4466_0_b(.in(layer_3[428]), .out(far_4_4466_0[1]));
    wire [1:0] far_4_4466_1;    relay_conn far_4_4466_1_a(.in(far_4_4466_0[0]), .out(far_4_4466_1[0]));    relay_conn far_4_4466_1_b(.in(far_4_4466_0[1]), .out(far_4_4466_1[1]));
    assign layer_4[386] = far_4_4466_1[1]; 
    assign layer_4[387] = ~layer_3[47]; 
    wire [1:0] far_4_4468_0;    relay_conn far_4_4468_0_a(.in(layer_3[692]), .out(far_4_4468_0[0]));    relay_conn far_4_4468_0_b(.in(layer_3[598]), .out(far_4_4468_0[1]));
    wire [1:0] far_4_4468_1;    relay_conn far_4_4468_1_a(.in(far_4_4468_0[0]), .out(far_4_4468_1[0]));    relay_conn far_4_4468_1_b(.in(far_4_4468_0[1]), .out(far_4_4468_1[1]));
    assign layer_4[388] = ~far_4_4468_1[0] | (far_4_4468_1[0] & far_4_4468_1[1]); 
    wire [1:0] far_4_4469_0;    relay_conn far_4_4469_0_a(.in(layer_3[47]), .out(far_4_4469_0[0]));    relay_conn far_4_4469_0_b(.in(layer_3[148]), .out(far_4_4469_0[1]));
    wire [1:0] far_4_4469_1;    relay_conn far_4_4469_1_a(.in(far_4_4469_0[0]), .out(far_4_4469_1[0]));    relay_conn far_4_4469_1_b(.in(far_4_4469_0[1]), .out(far_4_4469_1[1]));
    wire [1:0] far_4_4469_2;    relay_conn far_4_4469_2_a(.in(far_4_4469_1[0]), .out(far_4_4469_2[0]));    relay_conn far_4_4469_2_b(.in(far_4_4469_1[1]), .out(far_4_4469_2[1]));
    assign layer_4[389] = ~far_4_4469_2[0] | (far_4_4469_2[0] & far_4_4469_2[1]); 
    wire [1:0] far_4_4470_0;    relay_conn far_4_4470_0_a(.in(layer_3[337]), .out(far_4_4470_0[0]));    relay_conn far_4_4470_0_b(.in(layer_3[253]), .out(far_4_4470_0[1]));
    wire [1:0] far_4_4470_1;    relay_conn far_4_4470_1_a(.in(far_4_4470_0[0]), .out(far_4_4470_1[0]));    relay_conn far_4_4470_1_b(.in(far_4_4470_0[1]), .out(far_4_4470_1[1]));
    assign layer_4[390] = far_4_4470_1[0] ^ far_4_4470_1[1]; 
    wire [1:0] far_4_4471_0;    relay_conn far_4_4471_0_a(.in(layer_3[546]), .out(far_4_4471_0[0]));    relay_conn far_4_4471_0_b(.in(layer_3[426]), .out(far_4_4471_0[1]));
    wire [1:0] far_4_4471_1;    relay_conn far_4_4471_1_a(.in(far_4_4471_0[0]), .out(far_4_4471_1[0]));    relay_conn far_4_4471_1_b(.in(far_4_4471_0[1]), .out(far_4_4471_1[1]));
    wire [1:0] far_4_4471_2;    relay_conn far_4_4471_2_a(.in(far_4_4471_1[0]), .out(far_4_4471_2[0]));    relay_conn far_4_4471_2_b(.in(far_4_4471_1[1]), .out(far_4_4471_2[1]));
    assign layer_4[391] = far_4_4471_2[1]; 
    wire [1:0] far_4_4472_0;    relay_conn far_4_4472_0_a(.in(layer_3[864]), .out(far_4_4472_0[0]));    relay_conn far_4_4472_0_b(.in(layer_3[799]), .out(far_4_4472_0[1]));
    wire [1:0] far_4_4472_1;    relay_conn far_4_4472_1_a(.in(far_4_4472_0[0]), .out(far_4_4472_1[0]));    relay_conn far_4_4472_1_b(.in(far_4_4472_0[1]), .out(far_4_4472_1[1]));
    assign layer_4[392] = ~(far_4_4472_1[0] & far_4_4472_1[1]); 
    assign layer_4[393] = layer_3[90] | layer_3[114]; 
    wire [1:0] far_4_4474_0;    relay_conn far_4_4474_0_a(.in(layer_3[895]), .out(far_4_4474_0[0]));    relay_conn far_4_4474_0_b(.in(layer_3[861]), .out(far_4_4474_0[1]));
    assign layer_4[394] = far_4_4474_0[0] & ~far_4_4474_0[1]; 
    assign layer_4[395] = ~layer_3[164]; 
    assign layer_4[396] = layer_3[556] & ~layer_3[577]; 
    assign layer_4[397] = layer_3[353] & ~layer_3[323]; 
    assign layer_4[398] = ~(layer_3[760] & layer_3[738]); 
    assign layer_4[399] = ~layer_3[805] | (layer_3[781] & layer_3[805]); 
    wire [1:0] far_4_4480_0;    relay_conn far_4_4480_0_a(.in(layer_3[682]), .out(far_4_4480_0[0]));    relay_conn far_4_4480_0_b(.in(layer_3[634]), .out(far_4_4480_0[1]));
    assign layer_4[400] = ~far_4_4480_0[0] | (far_4_4480_0[0] & far_4_4480_0[1]); 
    wire [1:0] far_4_4481_0;    relay_conn far_4_4481_0_a(.in(layer_3[725]), .out(far_4_4481_0[0]));    relay_conn far_4_4481_0_b(.in(layer_3[782]), .out(far_4_4481_0[1]));
    assign layer_4[401] = ~far_4_4481_0[1]; 
    wire [1:0] far_4_4482_0;    relay_conn far_4_4482_0_a(.in(layer_3[336]), .out(far_4_4482_0[0]));    relay_conn far_4_4482_0_b(.in(layer_3[300]), .out(far_4_4482_0[1]));
    assign layer_4[402] = ~(far_4_4482_0[0] | far_4_4482_0[1]); 
    wire [1:0] far_4_4483_0;    relay_conn far_4_4483_0_a(.in(layer_3[154]), .out(far_4_4483_0[0]));    relay_conn far_4_4483_0_b(.in(layer_3[202]), .out(far_4_4483_0[1]));
    assign layer_4[403] = ~far_4_4483_0[0]; 
    wire [1:0] far_4_4484_0;    relay_conn far_4_4484_0_a(.in(layer_3[424]), .out(far_4_4484_0[0]));    relay_conn far_4_4484_0_b(.in(layer_3[362]), .out(far_4_4484_0[1]));
    assign layer_4[404] = ~far_4_4484_0[0] | (far_4_4484_0[0] & far_4_4484_0[1]); 
    wire [1:0] far_4_4485_0;    relay_conn far_4_4485_0_a(.in(layer_3[711]), .out(far_4_4485_0[0]));    relay_conn far_4_4485_0_b(.in(layer_3[632]), .out(far_4_4485_0[1]));
    wire [1:0] far_4_4485_1;    relay_conn far_4_4485_1_a(.in(far_4_4485_0[0]), .out(far_4_4485_1[0]));    relay_conn far_4_4485_1_b(.in(far_4_4485_0[1]), .out(far_4_4485_1[1]));
    assign layer_4[405] = ~(far_4_4485_1[0] | far_4_4485_1[1]); 
    wire [1:0] far_4_4486_0;    relay_conn far_4_4486_0_a(.in(layer_3[818]), .out(far_4_4486_0[0]));    relay_conn far_4_4486_0_b(.in(layer_3[782]), .out(far_4_4486_0[1]));
    assign layer_4[406] = far_4_4486_0[0] & far_4_4486_0[1]; 
    wire [1:0] far_4_4487_0;    relay_conn far_4_4487_0_a(.in(layer_3[883]), .out(far_4_4487_0[0]));    relay_conn far_4_4487_0_b(.in(layer_3[846]), .out(far_4_4487_0[1]));
    assign layer_4[407] = far_4_4487_0[0] & far_4_4487_0[1]; 
    wire [1:0] far_4_4488_0;    relay_conn far_4_4488_0_a(.in(layer_3[610]), .out(far_4_4488_0[0]));    relay_conn far_4_4488_0_b(.in(layer_3[733]), .out(far_4_4488_0[1]));
    wire [1:0] far_4_4488_1;    relay_conn far_4_4488_1_a(.in(far_4_4488_0[0]), .out(far_4_4488_1[0]));    relay_conn far_4_4488_1_b(.in(far_4_4488_0[1]), .out(far_4_4488_1[1]));
    wire [1:0] far_4_4488_2;    relay_conn far_4_4488_2_a(.in(far_4_4488_1[0]), .out(far_4_4488_2[0]));    relay_conn far_4_4488_2_b(.in(far_4_4488_1[1]), .out(far_4_4488_2[1]));
    assign layer_4[408] = ~far_4_4488_2[0] | (far_4_4488_2[0] & far_4_4488_2[1]); 
    wire [1:0] far_4_4489_0;    relay_conn far_4_4489_0_a(.in(layer_3[297]), .out(far_4_4489_0[0]));    relay_conn far_4_4489_0_b(.in(layer_3[346]), .out(far_4_4489_0[1]));
    assign layer_4[409] = ~far_4_4489_0[1] | (far_4_4489_0[0] & far_4_4489_0[1]); 
    wire [1:0] far_4_4490_0;    relay_conn far_4_4490_0_a(.in(layer_3[117]), .out(far_4_4490_0[0]));    relay_conn far_4_4490_0_b(.in(layer_3[75]), .out(far_4_4490_0[1]));
    assign layer_4[410] = ~far_4_4490_0[1] | (far_4_4490_0[0] & far_4_4490_0[1]); 
    wire [1:0] far_4_4491_0;    relay_conn far_4_4491_0_a(.in(layer_3[551]), .out(far_4_4491_0[0]));    relay_conn far_4_4491_0_b(.in(layer_3[468]), .out(far_4_4491_0[1]));
    wire [1:0] far_4_4491_1;    relay_conn far_4_4491_1_a(.in(far_4_4491_0[0]), .out(far_4_4491_1[0]));    relay_conn far_4_4491_1_b(.in(far_4_4491_0[1]), .out(far_4_4491_1[1]));
    assign layer_4[411] = ~(far_4_4491_1[0] ^ far_4_4491_1[1]); 
    assign layer_4[412] = layer_3[393]; 
    assign layer_4[413] = layer_3[908]; 
    wire [1:0] far_4_4494_0;    relay_conn far_4_4494_0_a(.in(layer_3[104]), .out(far_4_4494_0[0]));    relay_conn far_4_4494_0_b(.in(layer_3[217]), .out(far_4_4494_0[1]));
    wire [1:0] far_4_4494_1;    relay_conn far_4_4494_1_a(.in(far_4_4494_0[0]), .out(far_4_4494_1[0]));    relay_conn far_4_4494_1_b(.in(far_4_4494_0[1]), .out(far_4_4494_1[1]));
    wire [1:0] far_4_4494_2;    relay_conn far_4_4494_2_a(.in(far_4_4494_1[0]), .out(far_4_4494_2[0]));    relay_conn far_4_4494_2_b(.in(far_4_4494_1[1]), .out(far_4_4494_2[1]));
    assign layer_4[414] = far_4_4494_2[0] ^ far_4_4494_2[1]; 
    wire [1:0] far_4_4495_0;    relay_conn far_4_4495_0_a(.in(layer_3[21]), .out(far_4_4495_0[0]));    relay_conn far_4_4495_0_b(.in(layer_3[100]), .out(far_4_4495_0[1]));
    wire [1:0] far_4_4495_1;    relay_conn far_4_4495_1_a(.in(far_4_4495_0[0]), .out(far_4_4495_1[0]));    relay_conn far_4_4495_1_b(.in(far_4_4495_0[1]), .out(far_4_4495_1[1]));
    assign layer_4[415] = far_4_4495_1[1]; 
    assign layer_4[416] = layer_3[402]; 
    assign layer_4[417] = layer_3[400] | layer_3[408]; 
    wire [1:0] far_4_4498_0;    relay_conn far_4_4498_0_a(.in(layer_3[323]), .out(far_4_4498_0[0]));    relay_conn far_4_4498_0_b(.in(layer_3[386]), .out(far_4_4498_0[1]));
    assign layer_4[418] = ~(far_4_4498_0[0] | far_4_4498_0[1]); 
    wire [1:0] far_4_4499_0;    relay_conn far_4_4499_0_a(.in(layer_3[459]), .out(far_4_4499_0[0]));    relay_conn far_4_4499_0_b(.in(layer_3[368]), .out(far_4_4499_0[1]));
    wire [1:0] far_4_4499_1;    relay_conn far_4_4499_1_a(.in(far_4_4499_0[0]), .out(far_4_4499_1[0]));    relay_conn far_4_4499_1_b(.in(far_4_4499_0[1]), .out(far_4_4499_1[1]));
    assign layer_4[419] = far_4_4499_1[0]; 
    wire [1:0] far_4_4500_0;    relay_conn far_4_4500_0_a(.in(layer_3[667]), .out(far_4_4500_0[0]));    relay_conn far_4_4500_0_b(.in(layer_3[770]), .out(far_4_4500_0[1]));
    wire [1:0] far_4_4500_1;    relay_conn far_4_4500_1_a(.in(far_4_4500_0[0]), .out(far_4_4500_1[0]));    relay_conn far_4_4500_1_b(.in(far_4_4500_0[1]), .out(far_4_4500_1[1]));
    wire [1:0] far_4_4500_2;    relay_conn far_4_4500_2_a(.in(far_4_4500_1[0]), .out(far_4_4500_2[0]));    relay_conn far_4_4500_2_b(.in(far_4_4500_1[1]), .out(far_4_4500_2[1]));
    assign layer_4[420] = ~(far_4_4500_2[0] | far_4_4500_2[1]); 
    wire [1:0] far_4_4501_0;    relay_conn far_4_4501_0_a(.in(layer_3[586]), .out(far_4_4501_0[0]));    relay_conn far_4_4501_0_b(.in(layer_3[483]), .out(far_4_4501_0[1]));
    wire [1:0] far_4_4501_1;    relay_conn far_4_4501_1_a(.in(far_4_4501_0[0]), .out(far_4_4501_1[0]));    relay_conn far_4_4501_1_b(.in(far_4_4501_0[1]), .out(far_4_4501_1[1]));
    wire [1:0] far_4_4501_2;    relay_conn far_4_4501_2_a(.in(far_4_4501_1[0]), .out(far_4_4501_2[0]));    relay_conn far_4_4501_2_b(.in(far_4_4501_1[1]), .out(far_4_4501_2[1]));
    assign layer_4[421] = far_4_4501_2[0] & far_4_4501_2[1]; 
    wire [1:0] far_4_4502_0;    relay_conn far_4_4502_0_a(.in(layer_3[268]), .out(far_4_4502_0[0]));    relay_conn far_4_4502_0_b(.in(layer_3[392]), .out(far_4_4502_0[1]));
    wire [1:0] far_4_4502_1;    relay_conn far_4_4502_1_a(.in(far_4_4502_0[0]), .out(far_4_4502_1[0]));    relay_conn far_4_4502_1_b(.in(far_4_4502_0[1]), .out(far_4_4502_1[1]));
    wire [1:0] far_4_4502_2;    relay_conn far_4_4502_2_a(.in(far_4_4502_1[0]), .out(far_4_4502_2[0]));    relay_conn far_4_4502_2_b(.in(far_4_4502_1[1]), .out(far_4_4502_2[1]));
    assign layer_4[422] = far_4_4502_2[1] & ~far_4_4502_2[0]; 
    wire [1:0] far_4_4503_0;    relay_conn far_4_4503_0_a(.in(layer_3[517]), .out(far_4_4503_0[0]));    relay_conn far_4_4503_0_b(.in(layer_3[578]), .out(far_4_4503_0[1]));
    assign layer_4[423] = ~far_4_4503_0[0] | (far_4_4503_0[0] & far_4_4503_0[1]); 
    wire [1:0] far_4_4504_0;    relay_conn far_4_4504_0_a(.in(layer_3[722]), .out(far_4_4504_0[0]));    relay_conn far_4_4504_0_b(.in(layer_3[633]), .out(far_4_4504_0[1]));
    wire [1:0] far_4_4504_1;    relay_conn far_4_4504_1_a(.in(far_4_4504_0[0]), .out(far_4_4504_1[0]));    relay_conn far_4_4504_1_b(.in(far_4_4504_0[1]), .out(far_4_4504_1[1]));
    assign layer_4[424] = ~far_4_4504_1[1] | (far_4_4504_1[0] & far_4_4504_1[1]); 
    wire [1:0] far_4_4505_0;    relay_conn far_4_4505_0_a(.in(layer_3[164]), .out(far_4_4505_0[0]));    relay_conn far_4_4505_0_b(.in(layer_3[222]), .out(far_4_4505_0[1]));
    assign layer_4[425] = far_4_4505_0[1]; 
    wire [1:0] far_4_4506_0;    relay_conn far_4_4506_0_a(.in(layer_3[682]), .out(far_4_4506_0[0]));    relay_conn far_4_4506_0_b(.in(layer_3[734]), .out(far_4_4506_0[1]));
    assign layer_4[426] = far_4_4506_0[0] | far_4_4506_0[1]; 
    assign layer_4[427] = layer_3[661]; 
    wire [1:0] far_4_4508_0;    relay_conn far_4_4508_0_a(.in(layer_3[924]), .out(far_4_4508_0[0]));    relay_conn far_4_4508_0_b(.in(layer_3[821]), .out(far_4_4508_0[1]));
    wire [1:0] far_4_4508_1;    relay_conn far_4_4508_1_a(.in(far_4_4508_0[0]), .out(far_4_4508_1[0]));    relay_conn far_4_4508_1_b(.in(far_4_4508_0[1]), .out(far_4_4508_1[1]));
    wire [1:0] far_4_4508_2;    relay_conn far_4_4508_2_a(.in(far_4_4508_1[0]), .out(far_4_4508_2[0]));    relay_conn far_4_4508_2_b(.in(far_4_4508_1[1]), .out(far_4_4508_2[1]));
    assign layer_4[428] = far_4_4508_2[0] | far_4_4508_2[1]; 
    wire [1:0] far_4_4509_0;    relay_conn far_4_4509_0_a(.in(layer_3[162]), .out(far_4_4509_0[0]));    relay_conn far_4_4509_0_b(.in(layer_3[73]), .out(far_4_4509_0[1]));
    wire [1:0] far_4_4509_1;    relay_conn far_4_4509_1_a(.in(far_4_4509_0[0]), .out(far_4_4509_1[0]));    relay_conn far_4_4509_1_b(.in(far_4_4509_0[1]), .out(far_4_4509_1[1]));
    assign layer_4[429] = ~(far_4_4509_1[0] & far_4_4509_1[1]); 
    wire [1:0] far_4_4510_0;    relay_conn far_4_4510_0_a(.in(layer_3[80]), .out(far_4_4510_0[0]));    relay_conn far_4_4510_0_b(.in(layer_3[7]), .out(far_4_4510_0[1]));
    wire [1:0] far_4_4510_1;    relay_conn far_4_4510_1_a(.in(far_4_4510_0[0]), .out(far_4_4510_1[0]));    relay_conn far_4_4510_1_b(.in(far_4_4510_0[1]), .out(far_4_4510_1[1]));
    assign layer_4[430] = ~(far_4_4510_1[0] & far_4_4510_1[1]); 
    assign layer_4[431] = ~layer_3[927] | (layer_3[927] & layer_3[932]); 
    wire [1:0] far_4_4512_0;    relay_conn far_4_4512_0_a(.in(layer_3[35]), .out(far_4_4512_0[0]));    relay_conn far_4_4512_0_b(.in(layer_3[100]), .out(far_4_4512_0[1]));
    wire [1:0] far_4_4512_1;    relay_conn far_4_4512_1_a(.in(far_4_4512_0[0]), .out(far_4_4512_1[0]));    relay_conn far_4_4512_1_b(.in(far_4_4512_0[1]), .out(far_4_4512_1[1]));
    assign layer_4[432] = ~(far_4_4512_1[0] | far_4_4512_1[1]); 
    assign layer_4[433] = ~layer_3[979] | (layer_3[959] & layer_3[979]); 
    wire [1:0] far_4_4514_0;    relay_conn far_4_4514_0_a(.in(layer_3[775]), .out(far_4_4514_0[0]));    relay_conn far_4_4514_0_b(.in(layer_3[674]), .out(far_4_4514_0[1]));
    wire [1:0] far_4_4514_1;    relay_conn far_4_4514_1_a(.in(far_4_4514_0[0]), .out(far_4_4514_1[0]));    relay_conn far_4_4514_1_b(.in(far_4_4514_0[1]), .out(far_4_4514_1[1]));
    wire [1:0] far_4_4514_2;    relay_conn far_4_4514_2_a(.in(far_4_4514_1[0]), .out(far_4_4514_2[0]));    relay_conn far_4_4514_2_b(.in(far_4_4514_1[1]), .out(far_4_4514_2[1]));
    assign layer_4[434] = far_4_4514_2[0]; 
    wire [1:0] far_4_4515_0;    relay_conn far_4_4515_0_a(.in(layer_3[801]), .out(far_4_4515_0[0]));    relay_conn far_4_4515_0_b(.in(layer_3[688]), .out(far_4_4515_0[1]));
    wire [1:0] far_4_4515_1;    relay_conn far_4_4515_1_a(.in(far_4_4515_0[0]), .out(far_4_4515_1[0]));    relay_conn far_4_4515_1_b(.in(far_4_4515_0[1]), .out(far_4_4515_1[1]));
    wire [1:0] far_4_4515_2;    relay_conn far_4_4515_2_a(.in(far_4_4515_1[0]), .out(far_4_4515_2[0]));    relay_conn far_4_4515_2_b(.in(far_4_4515_1[1]), .out(far_4_4515_2[1]));
    assign layer_4[435] = far_4_4515_2[0] | far_4_4515_2[1]; 
    wire [1:0] far_4_4516_0;    relay_conn far_4_4516_0_a(.in(layer_3[149]), .out(far_4_4516_0[0]));    relay_conn far_4_4516_0_b(.in(layer_3[100]), .out(far_4_4516_0[1]));
    assign layer_4[436] = ~far_4_4516_0[1]; 
    assign layer_4[437] = ~layer_3[790] | (layer_3[780] & layer_3[790]); 
    assign layer_4[438] = ~layer_3[221] | (layer_3[192] & layer_3[221]); 
    assign layer_4[439] = ~layer_3[562] | (layer_3[562] & layer_3[535]); 
    assign layer_4[440] = layer_3[546] & ~layer_3[542]; 
    assign layer_4[441] = ~(layer_3[1003] ^ layer_3[1000]); 
    wire [1:0] far_4_4522_0;    relay_conn far_4_4522_0_a(.in(layer_3[244]), .out(far_4_4522_0[0]));    relay_conn far_4_4522_0_b(.in(layer_3[345]), .out(far_4_4522_0[1]));
    wire [1:0] far_4_4522_1;    relay_conn far_4_4522_1_a(.in(far_4_4522_0[0]), .out(far_4_4522_1[0]));    relay_conn far_4_4522_1_b(.in(far_4_4522_0[1]), .out(far_4_4522_1[1]));
    wire [1:0] far_4_4522_2;    relay_conn far_4_4522_2_a(.in(far_4_4522_1[0]), .out(far_4_4522_2[0]));    relay_conn far_4_4522_2_b(.in(far_4_4522_1[1]), .out(far_4_4522_2[1]));
    assign layer_4[442] = far_4_4522_2[1]; 
    wire [1:0] far_4_4523_0;    relay_conn far_4_4523_0_a(.in(layer_3[629]), .out(far_4_4523_0[0]));    relay_conn far_4_4523_0_b(.in(layer_3[532]), .out(far_4_4523_0[1]));
    wire [1:0] far_4_4523_1;    relay_conn far_4_4523_1_a(.in(far_4_4523_0[0]), .out(far_4_4523_1[0]));    relay_conn far_4_4523_1_b(.in(far_4_4523_0[1]), .out(far_4_4523_1[1]));
    wire [1:0] far_4_4523_2;    relay_conn far_4_4523_2_a(.in(far_4_4523_1[0]), .out(far_4_4523_2[0]));    relay_conn far_4_4523_2_b(.in(far_4_4523_1[1]), .out(far_4_4523_2[1]));
    assign layer_4[443] = ~far_4_4523_2[1] | (far_4_4523_2[0] & far_4_4523_2[1]); 
    wire [1:0] far_4_4524_0;    relay_conn far_4_4524_0_a(.in(layer_3[414]), .out(far_4_4524_0[0]));    relay_conn far_4_4524_0_b(.in(layer_3[352]), .out(far_4_4524_0[1]));
    assign layer_4[444] = far_4_4524_0[0] & ~far_4_4524_0[1]; 
    wire [1:0] far_4_4525_0;    relay_conn far_4_4525_0_a(.in(layer_3[146]), .out(far_4_4525_0[0]));    relay_conn far_4_4525_0_b(.in(layer_3[35]), .out(far_4_4525_0[1]));
    wire [1:0] far_4_4525_1;    relay_conn far_4_4525_1_a(.in(far_4_4525_0[0]), .out(far_4_4525_1[0]));    relay_conn far_4_4525_1_b(.in(far_4_4525_0[1]), .out(far_4_4525_1[1]));
    wire [1:0] far_4_4525_2;    relay_conn far_4_4525_2_a(.in(far_4_4525_1[0]), .out(far_4_4525_2[0]));    relay_conn far_4_4525_2_b(.in(far_4_4525_1[1]), .out(far_4_4525_2[1]));
    assign layer_4[445] = far_4_4525_2[0] & ~far_4_4525_2[1]; 
    wire [1:0] far_4_4526_0;    relay_conn far_4_4526_0_a(.in(layer_3[656]), .out(far_4_4526_0[0]));    relay_conn far_4_4526_0_b(.in(layer_3[702]), .out(far_4_4526_0[1]));
    assign layer_4[446] = ~(far_4_4526_0[0] | far_4_4526_0[1]); 
    wire [1:0] far_4_4527_0;    relay_conn far_4_4527_0_a(.in(layer_3[935]), .out(far_4_4527_0[0]));    relay_conn far_4_4527_0_b(.in(layer_3[884]), .out(far_4_4527_0[1]));
    assign layer_4[447] = far_4_4527_0[0] & far_4_4527_0[1]; 
    assign layer_4[448] = ~(layer_3[512] & layer_3[507]); 
    wire [1:0] far_4_4529_0;    relay_conn far_4_4529_0_a(.in(layer_3[142]), .out(far_4_4529_0[0]));    relay_conn far_4_4529_0_b(.in(layer_3[36]), .out(far_4_4529_0[1]));
    wire [1:0] far_4_4529_1;    relay_conn far_4_4529_1_a(.in(far_4_4529_0[0]), .out(far_4_4529_1[0]));    relay_conn far_4_4529_1_b(.in(far_4_4529_0[1]), .out(far_4_4529_1[1]));
    wire [1:0] far_4_4529_2;    relay_conn far_4_4529_2_a(.in(far_4_4529_1[0]), .out(far_4_4529_2[0]));    relay_conn far_4_4529_2_b(.in(far_4_4529_1[1]), .out(far_4_4529_2[1]));
    assign layer_4[449] = ~(far_4_4529_2[0] | far_4_4529_2[1]); 
    wire [1:0] far_4_4530_0;    relay_conn far_4_4530_0_a(.in(layer_3[318]), .out(far_4_4530_0[0]));    relay_conn far_4_4530_0_b(.in(layer_3[400]), .out(far_4_4530_0[1]));
    wire [1:0] far_4_4530_1;    relay_conn far_4_4530_1_a(.in(far_4_4530_0[0]), .out(far_4_4530_1[0]));    relay_conn far_4_4530_1_b(.in(far_4_4530_0[1]), .out(far_4_4530_1[1]));
    assign layer_4[450] = ~(far_4_4530_1[0] | far_4_4530_1[1]); 
    assign layer_4[451] = ~(layer_3[576] | layer_3[569]); 
    wire [1:0] far_4_4532_0;    relay_conn far_4_4532_0_a(.in(layer_3[935]), .out(far_4_4532_0[0]));    relay_conn far_4_4532_0_b(.in(layer_3[1000]), .out(far_4_4532_0[1]));
    wire [1:0] far_4_4532_1;    relay_conn far_4_4532_1_a(.in(far_4_4532_0[0]), .out(far_4_4532_1[0]));    relay_conn far_4_4532_1_b(.in(far_4_4532_0[1]), .out(far_4_4532_1[1]));
    assign layer_4[452] = ~(far_4_4532_1[0] & far_4_4532_1[1]); 
    wire [1:0] far_4_4533_0;    relay_conn far_4_4533_0_a(.in(layer_3[835]), .out(far_4_4533_0[0]));    relay_conn far_4_4533_0_b(.in(layer_3[903]), .out(far_4_4533_0[1]));
    wire [1:0] far_4_4533_1;    relay_conn far_4_4533_1_a(.in(far_4_4533_0[0]), .out(far_4_4533_1[0]));    relay_conn far_4_4533_1_b(.in(far_4_4533_0[1]), .out(far_4_4533_1[1]));
    assign layer_4[453] = far_4_4533_1[1] & ~far_4_4533_1[0]; 
    wire [1:0] far_4_4534_0;    relay_conn far_4_4534_0_a(.in(layer_3[758]), .out(far_4_4534_0[0]));    relay_conn far_4_4534_0_b(.in(layer_3[682]), .out(far_4_4534_0[1]));
    wire [1:0] far_4_4534_1;    relay_conn far_4_4534_1_a(.in(far_4_4534_0[0]), .out(far_4_4534_1[0]));    relay_conn far_4_4534_1_b(.in(far_4_4534_0[1]), .out(far_4_4534_1[1]));
    assign layer_4[454] = far_4_4534_1[0]; 
    wire [1:0] far_4_4535_0;    relay_conn far_4_4535_0_a(.in(layer_3[251]), .out(far_4_4535_0[0]));    relay_conn far_4_4535_0_b(.in(layer_3[215]), .out(far_4_4535_0[1]));
    assign layer_4[455] = ~far_4_4535_0[0]; 
    wire [1:0] far_4_4536_0;    relay_conn far_4_4536_0_a(.in(layer_3[312]), .out(far_4_4536_0[0]));    relay_conn far_4_4536_0_b(.in(layer_3[348]), .out(far_4_4536_0[1]));
    assign layer_4[456] = far_4_4536_0[0] & far_4_4536_0[1]; 
    assign layer_4[457] = layer_3[158] | layer_3[168]; 
    wire [1:0] far_4_4538_0;    relay_conn far_4_4538_0_a(.in(layer_3[512]), .out(far_4_4538_0[0]));    relay_conn far_4_4538_0_b(.in(layer_3[410]), .out(far_4_4538_0[1]));
    wire [1:0] far_4_4538_1;    relay_conn far_4_4538_1_a(.in(far_4_4538_0[0]), .out(far_4_4538_1[0]));    relay_conn far_4_4538_1_b(.in(far_4_4538_0[1]), .out(far_4_4538_1[1]));
    wire [1:0] far_4_4538_2;    relay_conn far_4_4538_2_a(.in(far_4_4538_1[0]), .out(far_4_4538_2[0]));    relay_conn far_4_4538_2_b(.in(far_4_4538_1[1]), .out(far_4_4538_2[1]));
    assign layer_4[458] = ~(far_4_4538_2[0] & far_4_4538_2[1]); 
    assign layer_4[459] = layer_3[854] | layer_3[831]; 
    assign layer_4[460] = layer_3[154] ^ layer_3[179]; 
    assign layer_4[461] = ~layer_3[192]; 
    wire [1:0] far_4_4542_0;    relay_conn far_4_4542_0_a(.in(layer_3[785]), .out(far_4_4542_0[0]));    relay_conn far_4_4542_0_b(.in(layer_3[700]), .out(far_4_4542_0[1]));
    wire [1:0] far_4_4542_1;    relay_conn far_4_4542_1_a(.in(far_4_4542_0[0]), .out(far_4_4542_1[0]));    relay_conn far_4_4542_1_b(.in(far_4_4542_0[1]), .out(far_4_4542_1[1]));
    assign layer_4[462] = ~(far_4_4542_1[0] & far_4_4542_1[1]); 
    assign layer_4[463] = layer_3[948] & ~layer_3[977]; 
    wire [1:0] far_4_4544_0;    relay_conn far_4_4544_0_a(.in(layer_3[714]), .out(far_4_4544_0[0]));    relay_conn far_4_4544_0_b(.in(layer_3[648]), .out(far_4_4544_0[1]));
    wire [1:0] far_4_4544_1;    relay_conn far_4_4544_1_a(.in(far_4_4544_0[0]), .out(far_4_4544_1[0]));    relay_conn far_4_4544_1_b(.in(far_4_4544_0[1]), .out(far_4_4544_1[1]));
    assign layer_4[464] = far_4_4544_1[0] | far_4_4544_1[1]; 
    wire [1:0] far_4_4545_0;    relay_conn far_4_4545_0_a(.in(layer_3[834]), .out(far_4_4545_0[0]));    relay_conn far_4_4545_0_b(.in(layer_3[916]), .out(far_4_4545_0[1]));
    wire [1:0] far_4_4545_1;    relay_conn far_4_4545_1_a(.in(far_4_4545_0[0]), .out(far_4_4545_1[0]));    relay_conn far_4_4545_1_b(.in(far_4_4545_0[1]), .out(far_4_4545_1[1]));
    assign layer_4[465] = ~far_4_4545_1[1]; 
    wire [1:0] far_4_4546_0;    relay_conn far_4_4546_0_a(.in(layer_3[386]), .out(far_4_4546_0[0]));    relay_conn far_4_4546_0_b(.in(layer_3[331]), .out(far_4_4546_0[1]));
    assign layer_4[466] = ~far_4_4546_0[1]; 
    wire [1:0] far_4_4547_0;    relay_conn far_4_4547_0_a(.in(layer_3[278]), .out(far_4_4547_0[0]));    relay_conn far_4_4547_0_b(.in(layer_3[365]), .out(far_4_4547_0[1]));
    wire [1:0] far_4_4547_1;    relay_conn far_4_4547_1_a(.in(far_4_4547_0[0]), .out(far_4_4547_1[0]));    relay_conn far_4_4547_1_b(.in(far_4_4547_0[1]), .out(far_4_4547_1[1]));
    assign layer_4[467] = far_4_4547_1[0] ^ far_4_4547_1[1]; 
    wire [1:0] far_4_4548_0;    relay_conn far_4_4548_0_a(.in(layer_3[275]), .out(far_4_4548_0[0]));    relay_conn far_4_4548_0_b(.in(layer_3[337]), .out(far_4_4548_0[1]));
    assign layer_4[468] = ~far_4_4548_0[0] | (far_4_4548_0[0] & far_4_4548_0[1]); 
    assign layer_4[469] = layer_3[741] & ~layer_3[746]; 
    assign layer_4[470] = layer_3[400] | layer_3[414]; 
    wire [1:0] far_4_4551_0;    relay_conn far_4_4551_0_a(.in(layer_3[675]), .out(far_4_4551_0[0]));    relay_conn far_4_4551_0_b(.in(layer_3[596]), .out(far_4_4551_0[1]));
    wire [1:0] far_4_4551_1;    relay_conn far_4_4551_1_a(.in(far_4_4551_0[0]), .out(far_4_4551_1[0]));    relay_conn far_4_4551_1_b(.in(far_4_4551_0[1]), .out(far_4_4551_1[1]));
    assign layer_4[471] = ~far_4_4551_1[1]; 
    wire [1:0] far_4_4552_0;    relay_conn far_4_4552_0_a(.in(layer_3[197]), .out(far_4_4552_0[0]));    relay_conn far_4_4552_0_b(.in(layer_3[113]), .out(far_4_4552_0[1]));
    wire [1:0] far_4_4552_1;    relay_conn far_4_4552_1_a(.in(far_4_4552_0[0]), .out(far_4_4552_1[0]));    relay_conn far_4_4552_1_b(.in(far_4_4552_0[1]), .out(far_4_4552_1[1]));
    assign layer_4[472] = far_4_4552_1[1]; 
    assign layer_4[473] = ~layer_3[788]; 
    wire [1:0] far_4_4554_0;    relay_conn far_4_4554_0_a(.in(layer_3[884]), .out(far_4_4554_0[0]));    relay_conn far_4_4554_0_b(.in(layer_3[846]), .out(far_4_4554_0[1]));
    assign layer_4[474] = ~(far_4_4554_0[0] & far_4_4554_0[1]); 
    wire [1:0] far_4_4555_0;    relay_conn far_4_4555_0_a(.in(layer_3[164]), .out(far_4_4555_0[0]));    relay_conn far_4_4555_0_b(.in(layer_3[282]), .out(far_4_4555_0[1]));
    wire [1:0] far_4_4555_1;    relay_conn far_4_4555_1_a(.in(far_4_4555_0[0]), .out(far_4_4555_1[0]));    relay_conn far_4_4555_1_b(.in(far_4_4555_0[1]), .out(far_4_4555_1[1]));
    wire [1:0] far_4_4555_2;    relay_conn far_4_4555_2_a(.in(far_4_4555_1[0]), .out(far_4_4555_2[0]));    relay_conn far_4_4555_2_b(.in(far_4_4555_1[1]), .out(far_4_4555_2[1]));
    assign layer_4[475] = far_4_4555_2[1] & ~far_4_4555_2[0]; 
    wire [1:0] far_4_4556_0;    relay_conn far_4_4556_0_a(.in(layer_3[927]), .out(far_4_4556_0[0]));    relay_conn far_4_4556_0_b(.in(layer_3[835]), .out(far_4_4556_0[1]));
    wire [1:0] far_4_4556_1;    relay_conn far_4_4556_1_a(.in(far_4_4556_0[0]), .out(far_4_4556_1[0]));    relay_conn far_4_4556_1_b(.in(far_4_4556_0[1]), .out(far_4_4556_1[1]));
    assign layer_4[476] = far_4_4556_1[0]; 
    wire [1:0] far_4_4557_0;    relay_conn far_4_4557_0_a(.in(layer_3[503]), .out(far_4_4557_0[0]));    relay_conn far_4_4557_0_b(.in(layer_3[403]), .out(far_4_4557_0[1]));
    wire [1:0] far_4_4557_1;    relay_conn far_4_4557_1_a(.in(far_4_4557_0[0]), .out(far_4_4557_1[0]));    relay_conn far_4_4557_1_b(.in(far_4_4557_0[1]), .out(far_4_4557_1[1]));
    wire [1:0] far_4_4557_2;    relay_conn far_4_4557_2_a(.in(far_4_4557_1[0]), .out(far_4_4557_2[0]));    relay_conn far_4_4557_2_b(.in(far_4_4557_1[1]), .out(far_4_4557_2[1]));
    assign layer_4[477] = ~far_4_4557_2[1]; 
    wire [1:0] far_4_4558_0;    relay_conn far_4_4558_0_a(.in(layer_3[0]), .out(far_4_4558_0[0]));    relay_conn far_4_4558_0_b(.in(layer_3[113]), .out(far_4_4558_0[1]));
    wire [1:0] far_4_4558_1;    relay_conn far_4_4558_1_a(.in(far_4_4558_0[0]), .out(far_4_4558_1[0]));    relay_conn far_4_4558_1_b(.in(far_4_4558_0[1]), .out(far_4_4558_1[1]));
    wire [1:0] far_4_4558_2;    relay_conn far_4_4558_2_a(.in(far_4_4558_1[0]), .out(far_4_4558_2[0]));    relay_conn far_4_4558_2_b(.in(far_4_4558_1[1]), .out(far_4_4558_2[1]));
    assign layer_4[478] = far_4_4558_2[1]; 
    wire [1:0] far_4_4559_0;    relay_conn far_4_4559_0_a(.in(layer_3[68]), .out(far_4_4559_0[0]));    relay_conn far_4_4559_0_b(.in(layer_3[113]), .out(far_4_4559_0[1]));
    assign layer_4[479] = far_4_4559_0[1]; 
    wire [1:0] far_4_4560_0;    relay_conn far_4_4560_0_a(.in(layer_3[596]), .out(far_4_4560_0[0]));    relay_conn far_4_4560_0_b(.in(layer_3[564]), .out(far_4_4560_0[1]));
    assign layer_4[480] = far_4_4560_0[1] & ~far_4_4560_0[0]; 
    wire [1:0] far_4_4561_0;    relay_conn far_4_4561_0_a(.in(layer_3[769]), .out(far_4_4561_0[0]));    relay_conn far_4_4561_0_b(.in(layer_3[705]), .out(far_4_4561_0[1]));
    wire [1:0] far_4_4561_1;    relay_conn far_4_4561_1_a(.in(far_4_4561_0[0]), .out(far_4_4561_1[0]));    relay_conn far_4_4561_1_b(.in(far_4_4561_0[1]), .out(far_4_4561_1[1]));
    assign layer_4[481] = ~(far_4_4561_1[0] | far_4_4561_1[1]); 
    wire [1:0] far_4_4562_0;    relay_conn far_4_4562_0_a(.in(layer_3[654]), .out(far_4_4562_0[0]));    relay_conn far_4_4562_0_b(.in(layer_3[756]), .out(far_4_4562_0[1]));
    wire [1:0] far_4_4562_1;    relay_conn far_4_4562_1_a(.in(far_4_4562_0[0]), .out(far_4_4562_1[0]));    relay_conn far_4_4562_1_b(.in(far_4_4562_0[1]), .out(far_4_4562_1[1]));
    wire [1:0] far_4_4562_2;    relay_conn far_4_4562_2_a(.in(far_4_4562_1[0]), .out(far_4_4562_2[0]));    relay_conn far_4_4562_2_b(.in(far_4_4562_1[1]), .out(far_4_4562_2[1]));
    assign layer_4[482] = far_4_4562_2[0] & ~far_4_4562_2[1]; 
    wire [1:0] far_4_4563_0;    relay_conn far_4_4563_0_a(.in(layer_3[932]), .out(far_4_4563_0[0]));    relay_conn far_4_4563_0_b(.in(layer_3[809]), .out(far_4_4563_0[1]));
    wire [1:0] far_4_4563_1;    relay_conn far_4_4563_1_a(.in(far_4_4563_0[0]), .out(far_4_4563_1[0]));    relay_conn far_4_4563_1_b(.in(far_4_4563_0[1]), .out(far_4_4563_1[1]));
    wire [1:0] far_4_4563_2;    relay_conn far_4_4563_2_a(.in(far_4_4563_1[0]), .out(far_4_4563_2[0]));    relay_conn far_4_4563_2_b(.in(far_4_4563_1[1]), .out(far_4_4563_2[1]));
    assign layer_4[483] = ~far_4_4563_2[0]; 
    wire [1:0] far_4_4564_0;    relay_conn far_4_4564_0_a(.in(layer_3[157]), .out(far_4_4564_0[0]));    relay_conn far_4_4564_0_b(.in(layer_3[242]), .out(far_4_4564_0[1]));
    wire [1:0] far_4_4564_1;    relay_conn far_4_4564_1_a(.in(far_4_4564_0[0]), .out(far_4_4564_1[0]));    relay_conn far_4_4564_1_b(.in(far_4_4564_0[1]), .out(far_4_4564_1[1]));
    assign layer_4[484] = ~(far_4_4564_1[0] ^ far_4_4564_1[1]); 
    assign layer_4[485] = layer_3[165] & ~layer_3[140]; 
    wire [1:0] far_4_4566_0;    relay_conn far_4_4566_0_a(.in(layer_3[755]), .out(far_4_4566_0[0]));    relay_conn far_4_4566_0_b(.in(layer_3[865]), .out(far_4_4566_0[1]));
    wire [1:0] far_4_4566_1;    relay_conn far_4_4566_1_a(.in(far_4_4566_0[0]), .out(far_4_4566_1[0]));    relay_conn far_4_4566_1_b(.in(far_4_4566_0[1]), .out(far_4_4566_1[1]));
    wire [1:0] far_4_4566_2;    relay_conn far_4_4566_2_a(.in(far_4_4566_1[0]), .out(far_4_4566_2[0]));    relay_conn far_4_4566_2_b(.in(far_4_4566_1[1]), .out(far_4_4566_2[1]));
    assign layer_4[486] = far_4_4566_2[0] & far_4_4566_2[1]; 
    wire [1:0] far_4_4567_0;    relay_conn far_4_4567_0_a(.in(layer_3[625]), .out(far_4_4567_0[0]));    relay_conn far_4_4567_0_b(.in(layer_3[681]), .out(far_4_4567_0[1]));
    assign layer_4[487] = far_4_4567_0[1]; 
    assign layer_4[488] = ~layer_3[958]; 
    assign layer_4[489] = layer_3[56] & ~layer_3[52]; 
    wire [1:0] far_4_4570_0;    relay_conn far_4_4570_0_a(.in(layer_3[923]), .out(far_4_4570_0[0]));    relay_conn far_4_4570_0_b(.in(layer_3[958]), .out(far_4_4570_0[1]));
    assign layer_4[490] = far_4_4570_0[0] & ~far_4_4570_0[1]; 
    wire [1:0] far_4_4571_0;    relay_conn far_4_4571_0_a(.in(layer_3[975]), .out(far_4_4571_0[0]));    relay_conn far_4_4571_0_b(.in(layer_3[866]), .out(far_4_4571_0[1]));
    wire [1:0] far_4_4571_1;    relay_conn far_4_4571_1_a(.in(far_4_4571_0[0]), .out(far_4_4571_1[0]));    relay_conn far_4_4571_1_b(.in(far_4_4571_0[1]), .out(far_4_4571_1[1]));
    wire [1:0] far_4_4571_2;    relay_conn far_4_4571_2_a(.in(far_4_4571_1[0]), .out(far_4_4571_2[0]));    relay_conn far_4_4571_2_b(.in(far_4_4571_1[1]), .out(far_4_4571_2[1]));
    assign layer_4[491] = ~(far_4_4571_2[0] ^ far_4_4571_2[1]); 
    assign layer_4[492] = layer_3[883] ^ layer_3[868]; 
    wire [1:0] far_4_4573_0;    relay_conn far_4_4573_0_a(.in(layer_3[16]), .out(far_4_4573_0[0]));    relay_conn far_4_4573_0_b(.in(layer_3[101]), .out(far_4_4573_0[1]));
    wire [1:0] far_4_4573_1;    relay_conn far_4_4573_1_a(.in(far_4_4573_0[0]), .out(far_4_4573_1[0]));    relay_conn far_4_4573_1_b(.in(far_4_4573_0[1]), .out(far_4_4573_1[1]));
    assign layer_4[493] = ~far_4_4573_1[0] | (far_4_4573_1[0] & far_4_4573_1[1]); 
    wire [1:0] far_4_4574_0;    relay_conn far_4_4574_0_a(.in(layer_3[837]), .out(far_4_4574_0[0]));    relay_conn far_4_4574_0_b(.in(layer_3[885]), .out(far_4_4574_0[1]));
    assign layer_4[494] = ~far_4_4574_0[1]; 
    wire [1:0] far_4_4575_0;    relay_conn far_4_4575_0_a(.in(layer_3[72]), .out(far_4_4575_0[0]));    relay_conn far_4_4575_0_b(.in(layer_3[115]), .out(far_4_4575_0[1]));
    assign layer_4[495] = far_4_4575_0[1] & ~far_4_4575_0[0]; 
    wire [1:0] far_4_4576_0;    relay_conn far_4_4576_0_a(.in(layer_3[284]), .out(far_4_4576_0[0]));    relay_conn far_4_4576_0_b(.in(layer_3[182]), .out(far_4_4576_0[1]));
    wire [1:0] far_4_4576_1;    relay_conn far_4_4576_1_a(.in(far_4_4576_0[0]), .out(far_4_4576_1[0]));    relay_conn far_4_4576_1_b(.in(far_4_4576_0[1]), .out(far_4_4576_1[1]));
    wire [1:0] far_4_4576_2;    relay_conn far_4_4576_2_a(.in(far_4_4576_1[0]), .out(far_4_4576_2[0]));    relay_conn far_4_4576_2_b(.in(far_4_4576_1[1]), .out(far_4_4576_2[1]));
    assign layer_4[496] = ~(far_4_4576_2[0] | far_4_4576_2[1]); 
    assign layer_4[497] = ~layer_3[839] | (layer_3[839] & layer_3[849]); 
    wire [1:0] far_4_4578_0;    relay_conn far_4_4578_0_a(.in(layer_3[793]), .out(far_4_4578_0[0]));    relay_conn far_4_4578_0_b(.in(layer_3[746]), .out(far_4_4578_0[1]));
    assign layer_4[498] = far_4_4578_0[1] & ~far_4_4578_0[0]; 
    assign layer_4[499] = layer_3[475] | layer_3[484]; 
    assign layer_4[500] = layer_3[113]; 
    wire [1:0] far_4_4581_0;    relay_conn far_4_4581_0_a(.in(layer_3[749]), .out(far_4_4581_0[0]));    relay_conn far_4_4581_0_b(.in(layer_3[623]), .out(far_4_4581_0[1]));
    wire [1:0] far_4_4581_1;    relay_conn far_4_4581_1_a(.in(far_4_4581_0[0]), .out(far_4_4581_1[0]));    relay_conn far_4_4581_1_b(.in(far_4_4581_0[1]), .out(far_4_4581_1[1]));
    wire [1:0] far_4_4581_2;    relay_conn far_4_4581_2_a(.in(far_4_4581_1[0]), .out(far_4_4581_2[0]));    relay_conn far_4_4581_2_b(.in(far_4_4581_1[1]), .out(far_4_4581_2[1]));
    assign layer_4[501] = ~(far_4_4581_2[0] ^ far_4_4581_2[1]); 
    wire [1:0] far_4_4582_0;    relay_conn far_4_4582_0_a(.in(layer_3[503]), .out(far_4_4582_0[0]));    relay_conn far_4_4582_0_b(.in(layer_3[403]), .out(far_4_4582_0[1]));
    wire [1:0] far_4_4582_1;    relay_conn far_4_4582_1_a(.in(far_4_4582_0[0]), .out(far_4_4582_1[0]));    relay_conn far_4_4582_1_b(.in(far_4_4582_0[1]), .out(far_4_4582_1[1]));
    wire [1:0] far_4_4582_2;    relay_conn far_4_4582_2_a(.in(far_4_4582_1[0]), .out(far_4_4582_2[0]));    relay_conn far_4_4582_2_b(.in(far_4_4582_1[1]), .out(far_4_4582_2[1]));
    assign layer_4[502] = far_4_4582_2[0] & far_4_4582_2[1]; 
    wire [1:0] far_4_4583_0;    relay_conn far_4_4583_0_a(.in(layer_3[847]), .out(far_4_4583_0[0]));    relay_conn far_4_4583_0_b(.in(layer_3[921]), .out(far_4_4583_0[1]));
    wire [1:0] far_4_4583_1;    relay_conn far_4_4583_1_a(.in(far_4_4583_0[0]), .out(far_4_4583_1[0]));    relay_conn far_4_4583_1_b(.in(far_4_4583_0[1]), .out(far_4_4583_1[1]));
    assign layer_4[503] = far_4_4583_1[0] & far_4_4583_1[1]; 
    assign layer_4[504] = ~layer_3[97] | (layer_3[97] & layer_3[77]); 
    wire [1:0] far_4_4585_0;    relay_conn far_4_4585_0_a(.in(layer_3[815]), .out(far_4_4585_0[0]));    relay_conn far_4_4585_0_b(.in(layer_3[708]), .out(far_4_4585_0[1]));
    wire [1:0] far_4_4585_1;    relay_conn far_4_4585_1_a(.in(far_4_4585_0[0]), .out(far_4_4585_1[0]));    relay_conn far_4_4585_1_b(.in(far_4_4585_0[1]), .out(far_4_4585_1[1]));
    wire [1:0] far_4_4585_2;    relay_conn far_4_4585_2_a(.in(far_4_4585_1[0]), .out(far_4_4585_2[0]));    relay_conn far_4_4585_2_b(.in(far_4_4585_1[1]), .out(far_4_4585_2[1]));
    assign layer_4[505] = far_4_4585_2[0] | far_4_4585_2[1]; 
    wire [1:0] far_4_4586_0;    relay_conn far_4_4586_0_a(.in(layer_3[345]), .out(far_4_4586_0[0]));    relay_conn far_4_4586_0_b(.in(layer_3[272]), .out(far_4_4586_0[1]));
    wire [1:0] far_4_4586_1;    relay_conn far_4_4586_1_a(.in(far_4_4586_0[0]), .out(far_4_4586_1[0]));    relay_conn far_4_4586_1_b(.in(far_4_4586_0[1]), .out(far_4_4586_1[1]));
    assign layer_4[506] = far_4_4586_1[0] | far_4_4586_1[1]; 
    wire [1:0] far_4_4587_0;    relay_conn far_4_4587_0_a(.in(layer_3[129]), .out(far_4_4587_0[0]));    relay_conn far_4_4587_0_b(.in(layer_3[222]), .out(far_4_4587_0[1]));
    wire [1:0] far_4_4587_1;    relay_conn far_4_4587_1_a(.in(far_4_4587_0[0]), .out(far_4_4587_1[0]));    relay_conn far_4_4587_1_b(.in(far_4_4587_0[1]), .out(far_4_4587_1[1]));
    assign layer_4[507] = far_4_4587_1[0] & far_4_4587_1[1]; 
    wire [1:0] far_4_4588_0;    relay_conn far_4_4588_0_a(.in(layer_3[503]), .out(far_4_4588_0[0]));    relay_conn far_4_4588_0_b(.in(layer_3[577]), .out(far_4_4588_0[1]));
    wire [1:0] far_4_4588_1;    relay_conn far_4_4588_1_a(.in(far_4_4588_0[0]), .out(far_4_4588_1[0]));    relay_conn far_4_4588_1_b(.in(far_4_4588_0[1]), .out(far_4_4588_1[1]));
    assign layer_4[508] = ~far_4_4588_1[0] | (far_4_4588_1[0] & far_4_4588_1[1]); 
    wire [1:0] far_4_4589_0;    relay_conn far_4_4589_0_a(.in(layer_3[342]), .out(far_4_4589_0[0]));    relay_conn far_4_4589_0_b(.in(layer_3[451]), .out(far_4_4589_0[1]));
    wire [1:0] far_4_4589_1;    relay_conn far_4_4589_1_a(.in(far_4_4589_0[0]), .out(far_4_4589_1[0]));    relay_conn far_4_4589_1_b(.in(far_4_4589_0[1]), .out(far_4_4589_1[1]));
    wire [1:0] far_4_4589_2;    relay_conn far_4_4589_2_a(.in(far_4_4589_1[0]), .out(far_4_4589_2[0]));    relay_conn far_4_4589_2_b(.in(far_4_4589_1[1]), .out(far_4_4589_2[1]));
    assign layer_4[509] = far_4_4589_2[0] & ~far_4_4589_2[1]; 
    assign layer_4[510] = layer_3[813] | layer_3[800]; 
    assign layer_4[511] = layer_3[972] | layer_3[1003]; 
    wire [1:0] far_4_4592_0;    relay_conn far_4_4592_0_a(.in(layer_3[778]), .out(far_4_4592_0[0]));    relay_conn far_4_4592_0_b(.in(layer_3[815]), .out(far_4_4592_0[1]));
    assign layer_4[512] = far_4_4592_0[0]; 
    wire [1:0] far_4_4593_0;    relay_conn far_4_4593_0_a(.in(layer_3[402]), .out(far_4_4593_0[0]));    relay_conn far_4_4593_0_b(.in(layer_3[369]), .out(far_4_4593_0[1]));
    assign layer_4[513] = ~far_4_4593_0[0] | (far_4_4593_0[0] & far_4_4593_0[1]); 
    wire [1:0] far_4_4594_0;    relay_conn far_4_4594_0_a(.in(layer_3[608]), .out(far_4_4594_0[0]));    relay_conn far_4_4594_0_b(.in(layer_3[726]), .out(far_4_4594_0[1]));
    wire [1:0] far_4_4594_1;    relay_conn far_4_4594_1_a(.in(far_4_4594_0[0]), .out(far_4_4594_1[0]));    relay_conn far_4_4594_1_b(.in(far_4_4594_0[1]), .out(far_4_4594_1[1]));
    wire [1:0] far_4_4594_2;    relay_conn far_4_4594_2_a(.in(far_4_4594_1[0]), .out(far_4_4594_2[0]));    relay_conn far_4_4594_2_b(.in(far_4_4594_1[1]), .out(far_4_4594_2[1]));
    assign layer_4[514] = far_4_4594_2[0] & far_4_4594_2[1]; 
    wire [1:0] far_4_4595_0;    relay_conn far_4_4595_0_a(.in(layer_3[937]), .out(far_4_4595_0[0]));    relay_conn far_4_4595_0_b(.in(layer_3[866]), .out(far_4_4595_0[1]));
    wire [1:0] far_4_4595_1;    relay_conn far_4_4595_1_a(.in(far_4_4595_0[0]), .out(far_4_4595_1[0]));    relay_conn far_4_4595_1_b(.in(far_4_4595_0[1]), .out(far_4_4595_1[1]));
    assign layer_4[515] = far_4_4595_1[0] & far_4_4595_1[1]; 
    assign layer_4[516] = ~layer_3[671] | (layer_3[664] & layer_3[671]); 
    wire [1:0] far_4_4597_0;    relay_conn far_4_4597_0_a(.in(layer_3[905]), .out(far_4_4597_0[0]));    relay_conn far_4_4597_0_b(.in(layer_3[823]), .out(far_4_4597_0[1]));
    wire [1:0] far_4_4597_1;    relay_conn far_4_4597_1_a(.in(far_4_4597_0[0]), .out(far_4_4597_1[0]));    relay_conn far_4_4597_1_b(.in(far_4_4597_0[1]), .out(far_4_4597_1[1]));
    assign layer_4[517] = far_4_4597_1[0] | far_4_4597_1[1]; 
    wire [1:0] far_4_4598_0;    relay_conn far_4_4598_0_a(.in(layer_3[35]), .out(far_4_4598_0[0]));    relay_conn far_4_4598_0_b(.in(layer_3[112]), .out(far_4_4598_0[1]));
    wire [1:0] far_4_4598_1;    relay_conn far_4_4598_1_a(.in(far_4_4598_0[0]), .out(far_4_4598_1[0]));    relay_conn far_4_4598_1_b(.in(far_4_4598_0[1]), .out(far_4_4598_1[1]));
    assign layer_4[518] = ~far_4_4598_1[0] | (far_4_4598_1[0] & far_4_4598_1[1]); 
    assign layer_4[519] = ~layer_3[581]; 
    wire [1:0] far_4_4600_0;    relay_conn far_4_4600_0_a(.in(layer_3[567]), .out(far_4_4600_0[0]));    relay_conn far_4_4600_0_b(.in(layer_3[670]), .out(far_4_4600_0[1]));
    wire [1:0] far_4_4600_1;    relay_conn far_4_4600_1_a(.in(far_4_4600_0[0]), .out(far_4_4600_1[0]));    relay_conn far_4_4600_1_b(.in(far_4_4600_0[1]), .out(far_4_4600_1[1]));
    wire [1:0] far_4_4600_2;    relay_conn far_4_4600_2_a(.in(far_4_4600_1[0]), .out(far_4_4600_2[0]));    relay_conn far_4_4600_2_b(.in(far_4_4600_1[1]), .out(far_4_4600_2[1]));
    assign layer_4[520] = far_4_4600_2[0]; 
    wire [1:0] far_4_4601_0;    relay_conn far_4_4601_0_a(.in(layer_3[147]), .out(far_4_4601_0[0]));    relay_conn far_4_4601_0_b(.in(layer_3[37]), .out(far_4_4601_0[1]));
    wire [1:0] far_4_4601_1;    relay_conn far_4_4601_1_a(.in(far_4_4601_0[0]), .out(far_4_4601_1[0]));    relay_conn far_4_4601_1_b(.in(far_4_4601_0[1]), .out(far_4_4601_1[1]));
    wire [1:0] far_4_4601_2;    relay_conn far_4_4601_2_a(.in(far_4_4601_1[0]), .out(far_4_4601_2[0]));    relay_conn far_4_4601_2_b(.in(far_4_4601_1[1]), .out(far_4_4601_2[1]));
    assign layer_4[521] = far_4_4601_2[0] | far_4_4601_2[1]; 
    wire [1:0] far_4_4602_0;    relay_conn far_4_4602_0_a(.in(layer_3[455]), .out(far_4_4602_0[0]));    relay_conn far_4_4602_0_b(.in(layer_3[345]), .out(far_4_4602_0[1]));
    wire [1:0] far_4_4602_1;    relay_conn far_4_4602_1_a(.in(far_4_4602_0[0]), .out(far_4_4602_1[0]));    relay_conn far_4_4602_1_b(.in(far_4_4602_0[1]), .out(far_4_4602_1[1]));
    wire [1:0] far_4_4602_2;    relay_conn far_4_4602_2_a(.in(far_4_4602_1[0]), .out(far_4_4602_2[0]));    relay_conn far_4_4602_2_b(.in(far_4_4602_1[1]), .out(far_4_4602_2[1]));
    assign layer_4[522] = ~(far_4_4602_2[0] & far_4_4602_2[1]); 
    wire [1:0] far_4_4603_0;    relay_conn far_4_4603_0_a(.in(layer_3[202]), .out(far_4_4603_0[0]));    relay_conn far_4_4603_0_b(.in(layer_3[316]), .out(far_4_4603_0[1]));
    wire [1:0] far_4_4603_1;    relay_conn far_4_4603_1_a(.in(far_4_4603_0[0]), .out(far_4_4603_1[0]));    relay_conn far_4_4603_1_b(.in(far_4_4603_0[1]), .out(far_4_4603_1[1]));
    wire [1:0] far_4_4603_2;    relay_conn far_4_4603_2_a(.in(far_4_4603_1[0]), .out(far_4_4603_2[0]));    relay_conn far_4_4603_2_b(.in(far_4_4603_1[1]), .out(far_4_4603_2[1]));
    assign layer_4[523] = ~far_4_4603_2[1] | (far_4_4603_2[0] & far_4_4603_2[1]); 
    wire [1:0] far_4_4604_0;    relay_conn far_4_4604_0_a(.in(layer_3[627]), .out(far_4_4604_0[0]));    relay_conn far_4_4604_0_b(.in(layer_3[572]), .out(far_4_4604_0[1]));
    assign layer_4[524] = far_4_4604_0[0] | far_4_4604_0[1]; 
    wire [1:0] far_4_4605_0;    relay_conn far_4_4605_0_a(.in(layer_3[408]), .out(far_4_4605_0[0]));    relay_conn far_4_4605_0_b(.in(layer_3[374]), .out(far_4_4605_0[1]));
    assign layer_4[525] = far_4_4605_0[0]; 
    wire [1:0] far_4_4606_0;    relay_conn far_4_4606_0_a(.in(layer_3[953]), .out(far_4_4606_0[0]));    relay_conn far_4_4606_0_b(.in(layer_3[846]), .out(far_4_4606_0[1]));
    wire [1:0] far_4_4606_1;    relay_conn far_4_4606_1_a(.in(far_4_4606_0[0]), .out(far_4_4606_1[0]));    relay_conn far_4_4606_1_b(.in(far_4_4606_0[1]), .out(far_4_4606_1[1]));
    wire [1:0] far_4_4606_2;    relay_conn far_4_4606_2_a(.in(far_4_4606_1[0]), .out(far_4_4606_2[0]));    relay_conn far_4_4606_2_b(.in(far_4_4606_1[1]), .out(far_4_4606_2[1]));
    assign layer_4[526] = far_4_4606_2[0] ^ far_4_4606_2[1]; 
    wire [1:0] far_4_4607_0;    relay_conn far_4_4607_0_a(.in(layer_3[830]), .out(far_4_4607_0[0]));    relay_conn far_4_4607_0_b(.in(layer_3[775]), .out(far_4_4607_0[1]));
    assign layer_4[527] = far_4_4607_0[0]; 
    assign layer_4[528] = layer_3[348] & ~layer_3[354]; 
    wire [1:0] far_4_4609_0;    relay_conn far_4_4609_0_a(.in(layer_3[274]), .out(far_4_4609_0[0]));    relay_conn far_4_4609_0_b(.in(layer_3[323]), .out(far_4_4609_0[1]));
    assign layer_4[529] = ~(far_4_4609_0[0] ^ far_4_4609_0[1]); 
    wire [1:0] far_4_4610_0;    relay_conn far_4_4610_0_a(.in(layer_3[868]), .out(far_4_4610_0[0]));    relay_conn far_4_4610_0_b(.in(layer_3[782]), .out(far_4_4610_0[1]));
    wire [1:0] far_4_4610_1;    relay_conn far_4_4610_1_a(.in(far_4_4610_0[0]), .out(far_4_4610_1[0]));    relay_conn far_4_4610_1_b(.in(far_4_4610_0[1]), .out(far_4_4610_1[1]));
    assign layer_4[530] = far_4_4610_1[1]; 
    wire [1:0] far_4_4611_0;    relay_conn far_4_4611_0_a(.in(layer_3[255]), .out(far_4_4611_0[0]));    relay_conn far_4_4611_0_b(.in(layer_3[212]), .out(far_4_4611_0[1]));
    assign layer_4[531] = ~far_4_4611_0[1] | (far_4_4611_0[0] & far_4_4611_0[1]); 
    wire [1:0] far_4_4612_0;    relay_conn far_4_4612_0_a(.in(layer_3[297]), .out(far_4_4612_0[0]));    relay_conn far_4_4612_0_b(.in(layer_3[179]), .out(far_4_4612_0[1]));
    wire [1:0] far_4_4612_1;    relay_conn far_4_4612_1_a(.in(far_4_4612_0[0]), .out(far_4_4612_1[0]));    relay_conn far_4_4612_1_b(.in(far_4_4612_0[1]), .out(far_4_4612_1[1]));
    wire [1:0] far_4_4612_2;    relay_conn far_4_4612_2_a(.in(far_4_4612_1[0]), .out(far_4_4612_2[0]));    relay_conn far_4_4612_2_b(.in(far_4_4612_1[1]), .out(far_4_4612_2[1]));
    assign layer_4[532] = ~far_4_4612_2[0]; 
    wire [1:0] far_4_4613_0;    relay_conn far_4_4613_0_a(.in(layer_3[420]), .out(far_4_4613_0[0]));    relay_conn far_4_4613_0_b(.in(layer_3[525]), .out(far_4_4613_0[1]));
    wire [1:0] far_4_4613_1;    relay_conn far_4_4613_1_a(.in(far_4_4613_0[0]), .out(far_4_4613_1[0]));    relay_conn far_4_4613_1_b(.in(far_4_4613_0[1]), .out(far_4_4613_1[1]));
    wire [1:0] far_4_4613_2;    relay_conn far_4_4613_2_a(.in(far_4_4613_1[0]), .out(far_4_4613_2[0]));    relay_conn far_4_4613_2_b(.in(far_4_4613_1[1]), .out(far_4_4613_2[1]));
    assign layer_4[533] = ~far_4_4613_2[0] | (far_4_4613_2[0] & far_4_4613_2[1]); 
    wire [1:0] far_4_4614_0;    relay_conn far_4_4614_0_a(.in(layer_3[169]), .out(far_4_4614_0[0]));    relay_conn far_4_4614_0_b(.in(layer_3[113]), .out(far_4_4614_0[1]));
    assign layer_4[534] = ~far_4_4614_0[1]; 
    wire [1:0] far_4_4615_0;    relay_conn far_4_4615_0_a(.in(layer_3[498]), .out(far_4_4615_0[0]));    relay_conn far_4_4615_0_b(.in(layer_3[391]), .out(far_4_4615_0[1]));
    wire [1:0] far_4_4615_1;    relay_conn far_4_4615_1_a(.in(far_4_4615_0[0]), .out(far_4_4615_1[0]));    relay_conn far_4_4615_1_b(.in(far_4_4615_0[1]), .out(far_4_4615_1[1]));
    wire [1:0] far_4_4615_2;    relay_conn far_4_4615_2_a(.in(far_4_4615_1[0]), .out(far_4_4615_2[0]));    relay_conn far_4_4615_2_b(.in(far_4_4615_1[1]), .out(far_4_4615_2[1]));
    assign layer_4[535] = far_4_4615_2[1] & ~far_4_4615_2[0]; 
    assign layer_4[536] = layer_3[931] | layer_3[919]; 
    wire [1:0] far_4_4617_0;    relay_conn far_4_4617_0_a(.in(layer_3[179]), .out(far_4_4617_0[0]));    relay_conn far_4_4617_0_b(.in(layer_3[147]), .out(far_4_4617_0[1]));
    assign layer_4[537] = far_4_4617_0[1] & ~far_4_4617_0[0]; 
    wire [1:0] far_4_4618_0;    relay_conn far_4_4618_0_a(.in(layer_3[478]), .out(far_4_4618_0[0]));    relay_conn far_4_4618_0_b(.in(layer_3[433]), .out(far_4_4618_0[1]));
    assign layer_4[538] = far_4_4618_0[0] | far_4_4618_0[1]; 
    assign layer_4[539] = ~layer_3[605]; 
    wire [1:0] far_4_4620_0;    relay_conn far_4_4620_0_a(.in(layer_3[317]), .out(far_4_4620_0[0]));    relay_conn far_4_4620_0_b(.in(layer_3[443]), .out(far_4_4620_0[1]));
    wire [1:0] far_4_4620_1;    relay_conn far_4_4620_1_a(.in(far_4_4620_0[0]), .out(far_4_4620_1[0]));    relay_conn far_4_4620_1_b(.in(far_4_4620_0[1]), .out(far_4_4620_1[1]));
    wire [1:0] far_4_4620_2;    relay_conn far_4_4620_2_a(.in(far_4_4620_1[0]), .out(far_4_4620_2[0]));    relay_conn far_4_4620_2_b(.in(far_4_4620_1[1]), .out(far_4_4620_2[1]));
    assign layer_4[540] = far_4_4620_2[0] & ~far_4_4620_2[1]; 
    wire [1:0] far_4_4621_0;    relay_conn far_4_4621_0_a(.in(layer_3[846]), .out(far_4_4621_0[0]));    relay_conn far_4_4621_0_b(.in(layer_3[738]), .out(far_4_4621_0[1]));
    wire [1:0] far_4_4621_1;    relay_conn far_4_4621_1_a(.in(far_4_4621_0[0]), .out(far_4_4621_1[0]));    relay_conn far_4_4621_1_b(.in(far_4_4621_0[1]), .out(far_4_4621_1[1]));
    wire [1:0] far_4_4621_2;    relay_conn far_4_4621_2_a(.in(far_4_4621_1[0]), .out(far_4_4621_2[0]));    relay_conn far_4_4621_2_b(.in(far_4_4621_1[1]), .out(far_4_4621_2[1]));
    assign layer_4[541] = ~(far_4_4621_2[0] | far_4_4621_2[1]); 
    wire [1:0] far_4_4622_0;    relay_conn far_4_4622_0_a(.in(layer_3[323]), .out(far_4_4622_0[0]));    relay_conn far_4_4622_0_b(.in(layer_3[416]), .out(far_4_4622_0[1]));
    wire [1:0] far_4_4622_1;    relay_conn far_4_4622_1_a(.in(far_4_4622_0[0]), .out(far_4_4622_1[0]));    relay_conn far_4_4622_1_b(.in(far_4_4622_0[1]), .out(far_4_4622_1[1]));
    assign layer_4[542] = ~far_4_4622_1[0] | (far_4_4622_1[0] & far_4_4622_1[1]); 
    assign layer_4[543] = ~layer_3[143]; 
    wire [1:0] far_4_4624_0;    relay_conn far_4_4624_0_a(.in(layer_3[337]), .out(far_4_4624_0[0]));    relay_conn far_4_4624_0_b(.in(layer_3[408]), .out(far_4_4624_0[1]));
    wire [1:0] far_4_4624_1;    relay_conn far_4_4624_1_a(.in(far_4_4624_0[0]), .out(far_4_4624_1[0]));    relay_conn far_4_4624_1_b(.in(far_4_4624_0[1]), .out(far_4_4624_1[1]));
    assign layer_4[544] = ~far_4_4624_1[0] | (far_4_4624_1[0] & far_4_4624_1[1]); 
    wire [1:0] far_4_4625_0;    relay_conn far_4_4625_0_a(.in(layer_3[165]), .out(far_4_4625_0[0]));    relay_conn far_4_4625_0_b(.in(layer_3[105]), .out(far_4_4625_0[1]));
    assign layer_4[545] = ~(far_4_4625_0[0] | far_4_4625_0[1]); 
    wire [1:0] far_4_4626_0;    relay_conn far_4_4626_0_a(.in(layer_3[908]), .out(far_4_4626_0[0]));    relay_conn far_4_4626_0_b(.in(layer_3[781]), .out(far_4_4626_0[1]));
    wire [1:0] far_4_4626_1;    relay_conn far_4_4626_1_a(.in(far_4_4626_0[0]), .out(far_4_4626_1[0]));    relay_conn far_4_4626_1_b(.in(far_4_4626_0[1]), .out(far_4_4626_1[1]));
    wire [1:0] far_4_4626_2;    relay_conn far_4_4626_2_a(.in(far_4_4626_1[0]), .out(far_4_4626_2[0]));    relay_conn far_4_4626_2_b(.in(far_4_4626_1[1]), .out(far_4_4626_2[1]));
    assign layer_4[546] = ~far_4_4626_2[1] | (far_4_4626_2[0] & far_4_4626_2[1]); 
    wire [1:0] far_4_4627_0;    relay_conn far_4_4627_0_a(.in(layer_3[305]), .out(far_4_4627_0[0]));    relay_conn far_4_4627_0_b(.in(layer_3[243]), .out(far_4_4627_0[1]));
    assign layer_4[547] = far_4_4627_0[1] & ~far_4_4627_0[0]; 
    wire [1:0] far_4_4628_0;    relay_conn far_4_4628_0_a(.in(layer_3[143]), .out(far_4_4628_0[0]));    relay_conn far_4_4628_0_b(.in(layer_3[266]), .out(far_4_4628_0[1]));
    wire [1:0] far_4_4628_1;    relay_conn far_4_4628_1_a(.in(far_4_4628_0[0]), .out(far_4_4628_1[0]));    relay_conn far_4_4628_1_b(.in(far_4_4628_0[1]), .out(far_4_4628_1[1]));
    wire [1:0] far_4_4628_2;    relay_conn far_4_4628_2_a(.in(far_4_4628_1[0]), .out(far_4_4628_2[0]));    relay_conn far_4_4628_2_b(.in(far_4_4628_1[1]), .out(far_4_4628_2[1]));
    assign layer_4[548] = ~far_4_4628_2[1]; 
    wire [1:0] far_4_4629_0;    relay_conn far_4_4629_0_a(.in(layer_3[674]), .out(far_4_4629_0[0]));    relay_conn far_4_4629_0_b(.in(layer_3[589]), .out(far_4_4629_0[1]));
    wire [1:0] far_4_4629_1;    relay_conn far_4_4629_1_a(.in(far_4_4629_0[0]), .out(far_4_4629_1[0]));    relay_conn far_4_4629_1_b(.in(far_4_4629_0[1]), .out(far_4_4629_1[1]));
    assign layer_4[549] = far_4_4629_1[1] & ~far_4_4629_1[0]; 
    wire [1:0] far_4_4630_0;    relay_conn far_4_4630_0_a(.in(layer_3[398]), .out(far_4_4630_0[0]));    relay_conn far_4_4630_0_b(.in(layer_3[498]), .out(far_4_4630_0[1]));
    wire [1:0] far_4_4630_1;    relay_conn far_4_4630_1_a(.in(far_4_4630_0[0]), .out(far_4_4630_1[0]));    relay_conn far_4_4630_1_b(.in(far_4_4630_0[1]), .out(far_4_4630_1[1]));
    wire [1:0] far_4_4630_2;    relay_conn far_4_4630_2_a(.in(far_4_4630_1[0]), .out(far_4_4630_2[0]));    relay_conn far_4_4630_2_b(.in(far_4_4630_1[1]), .out(far_4_4630_2[1]));
    assign layer_4[550] = far_4_4630_2[1] & ~far_4_4630_2[0]; 
    assign layer_4[551] = ~(layer_3[537] ^ layer_3[568]); 
    wire [1:0] far_4_4632_0;    relay_conn far_4_4632_0_a(.in(layer_3[909]), .out(far_4_4632_0[0]));    relay_conn far_4_4632_0_b(.in(layer_3[860]), .out(far_4_4632_0[1]));
    assign layer_4[552] = ~(far_4_4632_0[0] & far_4_4632_0[1]); 
    wire [1:0] far_4_4633_0;    relay_conn far_4_4633_0_a(.in(layer_3[470]), .out(far_4_4633_0[0]));    relay_conn far_4_4633_0_b(.in(layer_3[376]), .out(far_4_4633_0[1]));
    wire [1:0] far_4_4633_1;    relay_conn far_4_4633_1_a(.in(far_4_4633_0[0]), .out(far_4_4633_1[0]));    relay_conn far_4_4633_1_b(.in(far_4_4633_0[1]), .out(far_4_4633_1[1]));
    assign layer_4[553] = far_4_4633_1[1] & ~far_4_4633_1[0]; 
    wire [1:0] far_4_4634_0;    relay_conn far_4_4634_0_a(.in(layer_3[953]), .out(far_4_4634_0[0]));    relay_conn far_4_4634_0_b(.in(layer_3[843]), .out(far_4_4634_0[1]));
    wire [1:0] far_4_4634_1;    relay_conn far_4_4634_1_a(.in(far_4_4634_0[0]), .out(far_4_4634_1[0]));    relay_conn far_4_4634_1_b(.in(far_4_4634_0[1]), .out(far_4_4634_1[1]));
    wire [1:0] far_4_4634_2;    relay_conn far_4_4634_2_a(.in(far_4_4634_1[0]), .out(far_4_4634_2[0]));    relay_conn far_4_4634_2_b(.in(far_4_4634_1[1]), .out(far_4_4634_2[1]));
    assign layer_4[554] = far_4_4634_2[0] | far_4_4634_2[1]; 
    assign layer_4[555] = ~(layer_3[35] & layer_3[46]); 
    wire [1:0] far_4_4636_0;    relay_conn far_4_4636_0_a(.in(layer_3[121]), .out(far_4_4636_0[0]));    relay_conn far_4_4636_0_b(.in(layer_3[31]), .out(far_4_4636_0[1]));
    wire [1:0] far_4_4636_1;    relay_conn far_4_4636_1_a(.in(far_4_4636_0[0]), .out(far_4_4636_1[0]));    relay_conn far_4_4636_1_b(.in(far_4_4636_0[1]), .out(far_4_4636_1[1]));
    assign layer_4[556] = ~far_4_4636_1[1] | (far_4_4636_1[0] & far_4_4636_1[1]); 
    assign layer_4[557] = layer_3[276] & ~layer_3[289]; 
    assign layer_4[558] = layer_3[129] & ~layer_3[100]; 
    wire [1:0] far_4_4639_0;    relay_conn far_4_4639_0_a(.in(layer_3[556]), .out(far_4_4639_0[0]));    relay_conn far_4_4639_0_b(.in(layer_3[428]), .out(far_4_4639_0[1]));
    wire [1:0] far_4_4639_1;    relay_conn far_4_4639_1_a(.in(far_4_4639_0[0]), .out(far_4_4639_1[0]));    relay_conn far_4_4639_1_b(.in(far_4_4639_0[1]), .out(far_4_4639_1[1]));
    wire [1:0] far_4_4639_2;    relay_conn far_4_4639_2_a(.in(far_4_4639_1[0]), .out(far_4_4639_2[0]));    relay_conn far_4_4639_2_b(.in(far_4_4639_1[1]), .out(far_4_4639_2[1]));
    wire [1:0] far_4_4639_3;    relay_conn far_4_4639_3_a(.in(far_4_4639_2[0]), .out(far_4_4639_3[0]));    relay_conn far_4_4639_3_b(.in(far_4_4639_2[1]), .out(far_4_4639_3[1]));
    assign layer_4[559] = ~far_4_4639_3[1]; 
    wire [1:0] far_4_4640_0;    relay_conn far_4_4640_0_a(.in(layer_3[568]), .out(far_4_4640_0[0]));    relay_conn far_4_4640_0_b(.in(layer_3[525]), .out(far_4_4640_0[1]));
    assign layer_4[560] = ~far_4_4640_0[1]; 
    wire [1:0] far_4_4641_0;    relay_conn far_4_4641_0_a(.in(layer_3[525]), .out(far_4_4641_0[0]));    relay_conn far_4_4641_0_b(.in(layer_3[459]), .out(far_4_4641_0[1]));
    wire [1:0] far_4_4641_1;    relay_conn far_4_4641_1_a(.in(far_4_4641_0[0]), .out(far_4_4641_1[0]));    relay_conn far_4_4641_1_b(.in(far_4_4641_0[1]), .out(far_4_4641_1[1]));
    assign layer_4[561] = far_4_4641_1[1]; 
    wire [1:0] far_4_4642_0;    relay_conn far_4_4642_0_a(.in(layer_3[951]), .out(far_4_4642_0[0]));    relay_conn far_4_4642_0_b(.in(layer_3[847]), .out(far_4_4642_0[1]));
    wire [1:0] far_4_4642_1;    relay_conn far_4_4642_1_a(.in(far_4_4642_0[0]), .out(far_4_4642_1[0]));    relay_conn far_4_4642_1_b(.in(far_4_4642_0[1]), .out(far_4_4642_1[1]));
    wire [1:0] far_4_4642_2;    relay_conn far_4_4642_2_a(.in(far_4_4642_1[0]), .out(far_4_4642_2[0]));    relay_conn far_4_4642_2_b(.in(far_4_4642_1[1]), .out(far_4_4642_2[1]));
    assign layer_4[562] = ~(far_4_4642_2[0] | far_4_4642_2[1]); 
    wire [1:0] far_4_4643_0;    relay_conn far_4_4643_0_a(.in(layer_3[30]), .out(far_4_4643_0[0]));    relay_conn far_4_4643_0_b(.in(layer_3[104]), .out(far_4_4643_0[1]));
    wire [1:0] far_4_4643_1;    relay_conn far_4_4643_1_a(.in(far_4_4643_0[0]), .out(far_4_4643_1[0]));    relay_conn far_4_4643_1_b(.in(far_4_4643_0[1]), .out(far_4_4643_1[1]));
    assign layer_4[563] = ~far_4_4643_1[1]; 
    wire [1:0] far_4_4644_0;    relay_conn far_4_4644_0_a(.in(layer_3[498]), .out(far_4_4644_0[0]));    relay_conn far_4_4644_0_b(.in(layer_3[400]), .out(far_4_4644_0[1]));
    wire [1:0] far_4_4644_1;    relay_conn far_4_4644_1_a(.in(far_4_4644_0[0]), .out(far_4_4644_1[0]));    relay_conn far_4_4644_1_b(.in(far_4_4644_0[1]), .out(far_4_4644_1[1]));
    wire [1:0] far_4_4644_2;    relay_conn far_4_4644_2_a(.in(far_4_4644_1[0]), .out(far_4_4644_2[0]));    relay_conn far_4_4644_2_b(.in(far_4_4644_1[1]), .out(far_4_4644_2[1]));
    assign layer_4[564] = ~(far_4_4644_2[0] ^ far_4_4644_2[1]); 
    wire [1:0] far_4_4645_0;    relay_conn far_4_4645_0_a(.in(layer_3[70]), .out(far_4_4645_0[0]));    relay_conn far_4_4645_0_b(.in(layer_3[154]), .out(far_4_4645_0[1]));
    wire [1:0] far_4_4645_1;    relay_conn far_4_4645_1_a(.in(far_4_4645_0[0]), .out(far_4_4645_1[0]));    relay_conn far_4_4645_1_b(.in(far_4_4645_0[1]), .out(far_4_4645_1[1]));
    assign layer_4[565] = ~far_4_4645_1[0] | (far_4_4645_1[0] & far_4_4645_1[1]); 
    assign layer_4[566] = ~layer_3[779] | (layer_3[779] & layer_3[801]); 
    wire [1:0] far_4_4647_0;    relay_conn far_4_4647_0_a(.in(layer_3[718]), .out(far_4_4647_0[0]));    relay_conn far_4_4647_0_b(.in(layer_3[629]), .out(far_4_4647_0[1]));
    wire [1:0] far_4_4647_1;    relay_conn far_4_4647_1_a(.in(far_4_4647_0[0]), .out(far_4_4647_1[0]));    relay_conn far_4_4647_1_b(.in(far_4_4647_0[1]), .out(far_4_4647_1[1]));
    assign layer_4[567] = ~far_4_4647_1[0]; 
    wire [1:0] far_4_4648_0;    relay_conn far_4_4648_0_a(.in(layer_3[865]), .out(far_4_4648_0[0]));    relay_conn far_4_4648_0_b(.in(layer_3[950]), .out(far_4_4648_0[1]));
    wire [1:0] far_4_4648_1;    relay_conn far_4_4648_1_a(.in(far_4_4648_0[0]), .out(far_4_4648_1[0]));    relay_conn far_4_4648_1_b(.in(far_4_4648_0[1]), .out(far_4_4648_1[1]));
    assign layer_4[568] = far_4_4648_1[1] & ~far_4_4648_1[0]; 
    assign layer_4[569] = layer_3[708] | layer_3[738]; 
    assign layer_4[570] = ~(layer_3[953] | layer_3[941]); 
    assign layer_4[571] = ~(layer_3[402] & layer_3[428]); 
    wire [1:0] far_4_4652_0;    relay_conn far_4_4652_0_a(.in(layer_3[28]), .out(far_4_4652_0[0]));    relay_conn far_4_4652_0_b(.in(layer_3[72]), .out(far_4_4652_0[1]));
    assign layer_4[572] = ~far_4_4652_0[1] | (far_4_4652_0[0] & far_4_4652_0[1]); 
    assign layer_4[573] = ~layer_3[726] | (layer_3[726] & layer_3[725]); 
    wire [1:0] far_4_4654_0;    relay_conn far_4_4654_0_a(.in(layer_3[157]), .out(far_4_4654_0[0]));    relay_conn far_4_4654_0_b(.in(layer_3[210]), .out(far_4_4654_0[1]));
    assign layer_4[574] = far_4_4654_0[0]; 
    assign layer_4[575] = layer_3[248] & ~layer_3[274]; 
    wire [1:0] far_4_4656_0;    relay_conn far_4_4656_0_a(.in(layer_3[320]), .out(far_4_4656_0[0]));    relay_conn far_4_4656_0_b(.in(layer_3[194]), .out(far_4_4656_0[1]));
    wire [1:0] far_4_4656_1;    relay_conn far_4_4656_1_a(.in(far_4_4656_0[0]), .out(far_4_4656_1[0]));    relay_conn far_4_4656_1_b(.in(far_4_4656_0[1]), .out(far_4_4656_1[1]));
    wire [1:0] far_4_4656_2;    relay_conn far_4_4656_2_a(.in(far_4_4656_1[0]), .out(far_4_4656_2[0]));    relay_conn far_4_4656_2_b(.in(far_4_4656_1[1]), .out(far_4_4656_2[1]));
    assign layer_4[576] = ~far_4_4656_2[1]; 
    assign layer_4[577] = ~layer_3[673]; 
    wire [1:0] far_4_4658_0;    relay_conn far_4_4658_0_a(.in(layer_3[772]), .out(far_4_4658_0[0]));    relay_conn far_4_4658_0_b(.in(layer_3[839]), .out(far_4_4658_0[1]));
    wire [1:0] far_4_4658_1;    relay_conn far_4_4658_1_a(.in(far_4_4658_0[0]), .out(far_4_4658_1[0]));    relay_conn far_4_4658_1_b(.in(far_4_4658_0[1]), .out(far_4_4658_1[1]));
    assign layer_4[578] = far_4_4658_1[0] & ~far_4_4658_1[1]; 
    assign layer_4[579] = ~layer_3[632]; 
    assign layer_4[580] = ~layer_3[681]; 
    wire [1:0] far_4_4661_0;    relay_conn far_4_4661_0_a(.in(layer_3[255]), .out(far_4_4661_0[0]));    relay_conn far_4_4661_0_b(.in(layer_3[363]), .out(far_4_4661_0[1]));
    wire [1:0] far_4_4661_1;    relay_conn far_4_4661_1_a(.in(far_4_4661_0[0]), .out(far_4_4661_1[0]));    relay_conn far_4_4661_1_b(.in(far_4_4661_0[1]), .out(far_4_4661_1[1]));
    wire [1:0] far_4_4661_2;    relay_conn far_4_4661_2_a(.in(far_4_4661_1[0]), .out(far_4_4661_2[0]));    relay_conn far_4_4661_2_b(.in(far_4_4661_1[1]), .out(far_4_4661_2[1]));
    assign layer_4[581] = far_4_4661_2[0] & ~far_4_4661_2[1]; 
    wire [1:0] far_4_4662_0;    relay_conn far_4_4662_0_a(.in(layer_3[674]), .out(far_4_4662_0[0]));    relay_conn far_4_4662_0_b(.in(layer_3[609]), .out(far_4_4662_0[1]));
    wire [1:0] far_4_4662_1;    relay_conn far_4_4662_1_a(.in(far_4_4662_0[0]), .out(far_4_4662_1[0]));    relay_conn far_4_4662_1_b(.in(far_4_4662_0[1]), .out(far_4_4662_1[1]));
    assign layer_4[582] = ~(far_4_4662_1[0] & far_4_4662_1[1]); 
    wire [1:0] far_4_4663_0;    relay_conn far_4_4663_0_a(.in(layer_3[113]), .out(far_4_4663_0[0]));    relay_conn far_4_4663_0_b(.in(layer_3[32]), .out(far_4_4663_0[1]));
    wire [1:0] far_4_4663_1;    relay_conn far_4_4663_1_a(.in(far_4_4663_0[0]), .out(far_4_4663_1[0]));    relay_conn far_4_4663_1_b(.in(far_4_4663_0[1]), .out(far_4_4663_1[1]));
    assign layer_4[583] = far_4_4663_1[0] & far_4_4663_1[1]; 
    wire [1:0] far_4_4664_0;    relay_conn far_4_4664_0_a(.in(layer_3[801]), .out(far_4_4664_0[0]));    relay_conn far_4_4664_0_b(.in(layer_3[835]), .out(far_4_4664_0[1]));
    assign layer_4[584] = ~(far_4_4664_0[0] | far_4_4664_0[1]); 
    wire [1:0] far_4_4665_0;    relay_conn far_4_4665_0_a(.in(layer_3[101]), .out(far_4_4665_0[0]));    relay_conn far_4_4665_0_b(.in(layer_3[19]), .out(far_4_4665_0[1]));
    wire [1:0] far_4_4665_1;    relay_conn far_4_4665_1_a(.in(far_4_4665_0[0]), .out(far_4_4665_1[0]));    relay_conn far_4_4665_1_b(.in(far_4_4665_0[1]), .out(far_4_4665_1[1]));
    assign layer_4[585] = far_4_4665_1[1] & ~far_4_4665_1[0]; 
    assign layer_4[586] = layer_3[398]; 
    wire [1:0] far_4_4667_0;    relay_conn far_4_4667_0_a(.in(layer_3[443]), .out(far_4_4667_0[0]));    relay_conn far_4_4667_0_b(.in(layer_3[356]), .out(far_4_4667_0[1]));
    wire [1:0] far_4_4667_1;    relay_conn far_4_4667_1_a(.in(far_4_4667_0[0]), .out(far_4_4667_1[0]));    relay_conn far_4_4667_1_b(.in(far_4_4667_0[1]), .out(far_4_4667_1[1]));
    assign layer_4[587] = ~far_4_4667_1[1] | (far_4_4667_1[0] & far_4_4667_1[1]); 
    wire [1:0] far_4_4668_0;    relay_conn far_4_4668_0_a(.in(layer_3[75]), .out(far_4_4668_0[0]));    relay_conn far_4_4668_0_b(.in(layer_3[155]), .out(far_4_4668_0[1]));
    wire [1:0] far_4_4668_1;    relay_conn far_4_4668_1_a(.in(far_4_4668_0[0]), .out(far_4_4668_1[0]));    relay_conn far_4_4668_1_b(.in(far_4_4668_0[1]), .out(far_4_4668_1[1]));
    assign layer_4[588] = far_4_4668_1[0]; 
    wire [1:0] far_4_4669_0;    relay_conn far_4_4669_0_a(.in(layer_3[44]), .out(far_4_4669_0[0]));    relay_conn far_4_4669_0_b(.in(layer_3[140]), .out(far_4_4669_0[1]));
    wire [1:0] far_4_4669_1;    relay_conn far_4_4669_1_a(.in(far_4_4669_0[0]), .out(far_4_4669_1[0]));    relay_conn far_4_4669_1_b(.in(far_4_4669_0[1]), .out(far_4_4669_1[1]));
    wire [1:0] far_4_4669_2;    relay_conn far_4_4669_2_a(.in(far_4_4669_1[0]), .out(far_4_4669_2[0]));    relay_conn far_4_4669_2_b(.in(far_4_4669_1[1]), .out(far_4_4669_2[1]));
    assign layer_4[589] = ~(far_4_4669_2[0] | far_4_4669_2[1]); 
    wire [1:0] far_4_4670_0;    relay_conn far_4_4670_0_a(.in(layer_3[106]), .out(far_4_4670_0[0]));    relay_conn far_4_4670_0_b(.in(layer_3[35]), .out(far_4_4670_0[1]));
    wire [1:0] far_4_4670_1;    relay_conn far_4_4670_1_a(.in(far_4_4670_0[0]), .out(far_4_4670_1[0]));    relay_conn far_4_4670_1_b(.in(far_4_4670_0[1]), .out(far_4_4670_1[1]));
    assign layer_4[590] = ~(far_4_4670_1[0] & far_4_4670_1[1]); 
    assign layer_4[591] = layer_3[547] ^ layer_3[567]; 
    wire [1:0] far_4_4672_0;    relay_conn far_4_4672_0_a(.in(layer_3[744]), .out(far_4_4672_0[0]));    relay_conn far_4_4672_0_b(.in(layer_3[859]), .out(far_4_4672_0[1]));
    wire [1:0] far_4_4672_1;    relay_conn far_4_4672_1_a(.in(far_4_4672_0[0]), .out(far_4_4672_1[0]));    relay_conn far_4_4672_1_b(.in(far_4_4672_0[1]), .out(far_4_4672_1[1]));
    wire [1:0] far_4_4672_2;    relay_conn far_4_4672_2_a(.in(far_4_4672_1[0]), .out(far_4_4672_2[0]));    relay_conn far_4_4672_2_b(.in(far_4_4672_1[1]), .out(far_4_4672_2[1]));
    assign layer_4[592] = far_4_4672_2[0] & far_4_4672_2[1]; 
    assign layer_4[593] = ~layer_3[323]; 
    wire [1:0] far_4_4674_0;    relay_conn far_4_4674_0_a(.in(layer_3[556]), .out(far_4_4674_0[0]));    relay_conn far_4_4674_0_b(.in(layer_3[490]), .out(far_4_4674_0[1]));
    wire [1:0] far_4_4674_1;    relay_conn far_4_4674_1_a(.in(far_4_4674_0[0]), .out(far_4_4674_1[0]));    relay_conn far_4_4674_1_b(.in(far_4_4674_0[1]), .out(far_4_4674_1[1]));
    assign layer_4[594] = far_4_4674_1[0] & ~far_4_4674_1[1]; 
    wire [1:0] far_4_4675_0;    relay_conn far_4_4675_0_a(.in(layer_3[323]), .out(far_4_4675_0[0]));    relay_conn far_4_4675_0_b(.in(layer_3[264]), .out(far_4_4675_0[1]));
    assign layer_4[595] = ~(far_4_4675_0[0] & far_4_4675_0[1]); 
    wire [1:0] far_4_4676_0;    relay_conn far_4_4676_0_a(.in(layer_3[408]), .out(far_4_4676_0[0]));    relay_conn far_4_4676_0_b(.in(layer_3[318]), .out(far_4_4676_0[1]));
    wire [1:0] far_4_4676_1;    relay_conn far_4_4676_1_a(.in(far_4_4676_0[0]), .out(far_4_4676_1[0]));    relay_conn far_4_4676_1_b(.in(far_4_4676_0[1]), .out(far_4_4676_1[1]));
    assign layer_4[596] = ~(far_4_4676_1[0] | far_4_4676_1[1]); 
    wire [1:0] far_4_4677_0;    relay_conn far_4_4677_0_a(.in(layer_3[816]), .out(far_4_4677_0[0]));    relay_conn far_4_4677_0_b(.in(layer_3[927]), .out(far_4_4677_0[1]));
    wire [1:0] far_4_4677_1;    relay_conn far_4_4677_1_a(.in(far_4_4677_0[0]), .out(far_4_4677_1[0]));    relay_conn far_4_4677_1_b(.in(far_4_4677_0[1]), .out(far_4_4677_1[1]));
    wire [1:0] far_4_4677_2;    relay_conn far_4_4677_2_a(.in(far_4_4677_1[0]), .out(far_4_4677_2[0]));    relay_conn far_4_4677_2_b(.in(far_4_4677_1[1]), .out(far_4_4677_2[1]));
    assign layer_4[597] = ~far_4_4677_2[0] | (far_4_4677_2[0] & far_4_4677_2[1]); 
    wire [1:0] far_4_4678_0;    relay_conn far_4_4678_0_a(.in(layer_3[58]), .out(far_4_4678_0[0]));    relay_conn far_4_4678_0_b(.in(layer_3[94]), .out(far_4_4678_0[1]));
    assign layer_4[598] = far_4_4678_0[1] & ~far_4_4678_0[0]; 
    wire [1:0] far_4_4679_0;    relay_conn far_4_4679_0_a(.in(layer_3[692]), .out(far_4_4679_0[0]));    relay_conn far_4_4679_0_b(.in(layer_3[780]), .out(far_4_4679_0[1]));
    wire [1:0] far_4_4679_1;    relay_conn far_4_4679_1_a(.in(far_4_4679_0[0]), .out(far_4_4679_1[0]));    relay_conn far_4_4679_1_b(.in(far_4_4679_0[1]), .out(far_4_4679_1[1]));
    assign layer_4[599] = ~(far_4_4679_1[0] | far_4_4679_1[1]); 
    assign layer_4[600] = layer_3[681]; 
    wire [1:0] far_4_4681_0;    relay_conn far_4_4681_0_a(.in(layer_3[147]), .out(far_4_4681_0[0]));    relay_conn far_4_4681_0_b(.in(layer_3[36]), .out(far_4_4681_0[1]));
    wire [1:0] far_4_4681_1;    relay_conn far_4_4681_1_a(.in(far_4_4681_0[0]), .out(far_4_4681_1[0]));    relay_conn far_4_4681_1_b(.in(far_4_4681_0[1]), .out(far_4_4681_1[1]));
    wire [1:0] far_4_4681_2;    relay_conn far_4_4681_2_a(.in(far_4_4681_1[0]), .out(far_4_4681_2[0]));    relay_conn far_4_4681_2_b(.in(far_4_4681_1[1]), .out(far_4_4681_2[1]));
    assign layer_4[601] = far_4_4681_2[1] & ~far_4_4681_2[0]; 
    wire [1:0] far_4_4682_0;    relay_conn far_4_4682_0_a(.in(layer_3[394]), .out(far_4_4682_0[0]));    relay_conn far_4_4682_0_b(.in(layer_3[475]), .out(far_4_4682_0[1]));
    wire [1:0] far_4_4682_1;    relay_conn far_4_4682_1_a(.in(far_4_4682_0[0]), .out(far_4_4682_1[0]));    relay_conn far_4_4682_1_b(.in(far_4_4682_0[1]), .out(far_4_4682_1[1]));
    assign layer_4[602] = ~(far_4_4682_1[0] | far_4_4682_1[1]); 
    wire [1:0] far_4_4683_0;    relay_conn far_4_4683_0_a(.in(layer_3[716]), .out(far_4_4683_0[0]));    relay_conn far_4_4683_0_b(.in(layer_3[795]), .out(far_4_4683_0[1]));
    wire [1:0] far_4_4683_1;    relay_conn far_4_4683_1_a(.in(far_4_4683_0[0]), .out(far_4_4683_1[0]));    relay_conn far_4_4683_1_b(.in(far_4_4683_0[1]), .out(far_4_4683_1[1]));
    assign layer_4[603] = ~far_4_4683_1[1]; 
    wire [1:0] far_4_4684_0;    relay_conn far_4_4684_0_a(.in(layer_3[756]), .out(far_4_4684_0[0]));    relay_conn far_4_4684_0_b(.in(layer_3[855]), .out(far_4_4684_0[1]));
    wire [1:0] far_4_4684_1;    relay_conn far_4_4684_1_a(.in(far_4_4684_0[0]), .out(far_4_4684_1[0]));    relay_conn far_4_4684_1_b(.in(far_4_4684_0[1]), .out(far_4_4684_1[1]));
    wire [1:0] far_4_4684_2;    relay_conn far_4_4684_2_a(.in(far_4_4684_1[0]), .out(far_4_4684_2[0]));    relay_conn far_4_4684_2_b(.in(far_4_4684_1[1]), .out(far_4_4684_2[1]));
    assign layer_4[604] = ~far_4_4684_2[0]; 
    wire [1:0] far_4_4685_0;    relay_conn far_4_4685_0_a(.in(layer_3[113]), .out(far_4_4685_0[0]));    relay_conn far_4_4685_0_b(.in(layer_3[0]), .out(far_4_4685_0[1]));
    wire [1:0] far_4_4685_1;    relay_conn far_4_4685_1_a(.in(far_4_4685_0[0]), .out(far_4_4685_1[0]));    relay_conn far_4_4685_1_b(.in(far_4_4685_0[1]), .out(far_4_4685_1[1]));
    wire [1:0] far_4_4685_2;    relay_conn far_4_4685_2_a(.in(far_4_4685_1[0]), .out(far_4_4685_2[0]));    relay_conn far_4_4685_2_b(.in(far_4_4685_1[1]), .out(far_4_4685_2[1]));
    assign layer_4[605] = ~far_4_4685_2[0] | (far_4_4685_2[0] & far_4_4685_2[1]); 
    wire [1:0] far_4_4686_0;    relay_conn far_4_4686_0_a(.in(layer_3[532]), .out(far_4_4686_0[0]));    relay_conn far_4_4686_0_b(.in(layer_3[598]), .out(far_4_4686_0[1]));
    wire [1:0] far_4_4686_1;    relay_conn far_4_4686_1_a(.in(far_4_4686_0[0]), .out(far_4_4686_1[0]));    relay_conn far_4_4686_1_b(.in(far_4_4686_0[1]), .out(far_4_4686_1[1]));
    assign layer_4[606] = ~far_4_4686_1[1]; 
    assign layer_4[607] = layer_3[670]; 
    wire [1:0] far_4_4688_0;    relay_conn far_4_4688_0_a(.in(layer_3[868]), .out(far_4_4688_0[0]));    relay_conn far_4_4688_0_b(.in(layer_3[979]), .out(far_4_4688_0[1]));
    wire [1:0] far_4_4688_1;    relay_conn far_4_4688_1_a(.in(far_4_4688_0[0]), .out(far_4_4688_1[0]));    relay_conn far_4_4688_1_b(.in(far_4_4688_0[1]), .out(far_4_4688_1[1]));
    wire [1:0] far_4_4688_2;    relay_conn far_4_4688_2_a(.in(far_4_4688_1[0]), .out(far_4_4688_2[0]));    relay_conn far_4_4688_2_b(.in(far_4_4688_1[1]), .out(far_4_4688_2[1]));
    assign layer_4[608] = ~far_4_4688_2[1]; 
    assign layer_4[609] = layer_3[59]; 
    wire [1:0] far_4_4690_0;    relay_conn far_4_4690_0_a(.in(layer_3[846]), .out(far_4_4690_0[0]));    relay_conn far_4_4690_0_b(.in(layer_3[953]), .out(far_4_4690_0[1]));
    wire [1:0] far_4_4690_1;    relay_conn far_4_4690_1_a(.in(far_4_4690_0[0]), .out(far_4_4690_1[0]));    relay_conn far_4_4690_1_b(.in(far_4_4690_0[1]), .out(far_4_4690_1[1]));
    wire [1:0] far_4_4690_2;    relay_conn far_4_4690_2_a(.in(far_4_4690_1[0]), .out(far_4_4690_2[0]));    relay_conn far_4_4690_2_b(.in(far_4_4690_1[1]), .out(far_4_4690_2[1]));
    assign layer_4[610] = ~(far_4_4690_2[0] ^ far_4_4690_2[1]); 
    assign layer_4[611] = layer_3[837]; 
    wire [1:0] far_4_4692_0;    relay_conn far_4_4692_0_a(.in(layer_3[712]), .out(far_4_4692_0[0]));    relay_conn far_4_4692_0_b(.in(layer_3[826]), .out(far_4_4692_0[1]));
    wire [1:0] far_4_4692_1;    relay_conn far_4_4692_1_a(.in(far_4_4692_0[0]), .out(far_4_4692_1[0]));    relay_conn far_4_4692_1_b(.in(far_4_4692_0[1]), .out(far_4_4692_1[1]));
    wire [1:0] far_4_4692_2;    relay_conn far_4_4692_2_a(.in(far_4_4692_1[0]), .out(far_4_4692_2[0]));    relay_conn far_4_4692_2_b(.in(far_4_4692_1[1]), .out(far_4_4692_2[1]));
    assign layer_4[612] = far_4_4692_2[1] & ~far_4_4692_2[0]; 
    wire [1:0] far_4_4693_0;    relay_conn far_4_4693_0_a(.in(layer_3[113]), .out(far_4_4693_0[0]));    relay_conn far_4_4693_0_b(.in(layer_3[15]), .out(far_4_4693_0[1]));
    wire [1:0] far_4_4693_1;    relay_conn far_4_4693_1_a(.in(far_4_4693_0[0]), .out(far_4_4693_1[0]));    relay_conn far_4_4693_1_b(.in(far_4_4693_0[1]), .out(far_4_4693_1[1]));
    wire [1:0] far_4_4693_2;    relay_conn far_4_4693_2_a(.in(far_4_4693_1[0]), .out(far_4_4693_2[0]));    relay_conn far_4_4693_2_b(.in(far_4_4693_1[1]), .out(far_4_4693_2[1]));
    assign layer_4[613] = ~far_4_4693_2[1]; 
    wire [1:0] far_4_4694_0;    relay_conn far_4_4694_0_a(.in(layer_3[773]), .out(far_4_4694_0[0]));    relay_conn far_4_4694_0_b(.in(layer_3[831]), .out(far_4_4694_0[1]));
    assign layer_4[614] = far_4_4694_0[1] & ~far_4_4694_0[0]; 
    wire [1:0] far_4_4695_0;    relay_conn far_4_4695_0_a(.in(layer_3[589]), .out(far_4_4695_0[0]));    relay_conn far_4_4695_0_b(.in(layer_3[555]), .out(far_4_4695_0[1]));
    assign layer_4[615] = ~(far_4_4695_0[0] & far_4_4695_0[1]); 
    wire [1:0] far_4_4696_0;    relay_conn far_4_4696_0_a(.in(layer_3[492]), .out(far_4_4696_0[0]));    relay_conn far_4_4696_0_b(.in(layer_3[619]), .out(far_4_4696_0[1]));
    wire [1:0] far_4_4696_1;    relay_conn far_4_4696_1_a(.in(far_4_4696_0[0]), .out(far_4_4696_1[0]));    relay_conn far_4_4696_1_b(.in(far_4_4696_0[1]), .out(far_4_4696_1[1]));
    wire [1:0] far_4_4696_2;    relay_conn far_4_4696_2_a(.in(far_4_4696_1[0]), .out(far_4_4696_2[0]));    relay_conn far_4_4696_2_b(.in(far_4_4696_1[1]), .out(far_4_4696_2[1]));
    assign layer_4[616] = far_4_4696_2[0]; 
    wire [1:0] far_4_4697_0;    relay_conn far_4_4697_0_a(.in(layer_3[796]), .out(far_4_4697_0[0]));    relay_conn far_4_4697_0_b(.in(layer_3[674]), .out(far_4_4697_0[1]));
    wire [1:0] far_4_4697_1;    relay_conn far_4_4697_1_a(.in(far_4_4697_0[0]), .out(far_4_4697_1[0]));    relay_conn far_4_4697_1_b(.in(far_4_4697_0[1]), .out(far_4_4697_1[1]));
    wire [1:0] far_4_4697_2;    relay_conn far_4_4697_2_a(.in(far_4_4697_1[0]), .out(far_4_4697_2[0]));    relay_conn far_4_4697_2_b(.in(far_4_4697_1[1]), .out(far_4_4697_2[1]));
    assign layer_4[617] = far_4_4697_2[0] & ~far_4_4697_2[1]; 
    wire [1:0] far_4_4698_0;    relay_conn far_4_4698_0_a(.in(layer_3[18]), .out(far_4_4698_0[0]));    relay_conn far_4_4698_0_b(.in(layer_3[136]), .out(far_4_4698_0[1]));
    wire [1:0] far_4_4698_1;    relay_conn far_4_4698_1_a(.in(far_4_4698_0[0]), .out(far_4_4698_1[0]));    relay_conn far_4_4698_1_b(.in(far_4_4698_0[1]), .out(far_4_4698_1[1]));
    wire [1:0] far_4_4698_2;    relay_conn far_4_4698_2_a(.in(far_4_4698_1[0]), .out(far_4_4698_2[0]));    relay_conn far_4_4698_2_b(.in(far_4_4698_1[1]), .out(far_4_4698_2[1]));
    assign layer_4[618] = far_4_4698_2[1] & ~far_4_4698_2[0]; 
    assign layer_4[619] = ~(layer_3[210] | layer_3[217]); 
    wire [1:0] far_4_4700_0;    relay_conn far_4_4700_0_a(.in(layer_3[593]), .out(far_4_4700_0[0]));    relay_conn far_4_4700_0_b(.in(layer_3[477]), .out(far_4_4700_0[1]));
    wire [1:0] far_4_4700_1;    relay_conn far_4_4700_1_a(.in(far_4_4700_0[0]), .out(far_4_4700_1[0]));    relay_conn far_4_4700_1_b(.in(far_4_4700_0[1]), .out(far_4_4700_1[1]));
    wire [1:0] far_4_4700_2;    relay_conn far_4_4700_2_a(.in(far_4_4700_1[0]), .out(far_4_4700_2[0]));    relay_conn far_4_4700_2_b(.in(far_4_4700_1[1]), .out(far_4_4700_2[1]));
    assign layer_4[620] = far_4_4700_2[1]; 
    wire [1:0] far_4_4701_0;    relay_conn far_4_4701_0_a(.in(layer_3[221]), .out(far_4_4701_0[0]));    relay_conn far_4_4701_0_b(.in(layer_3[303]), .out(far_4_4701_0[1]));
    wire [1:0] far_4_4701_1;    relay_conn far_4_4701_1_a(.in(far_4_4701_0[0]), .out(far_4_4701_1[0]));    relay_conn far_4_4701_1_b(.in(far_4_4701_0[1]), .out(far_4_4701_1[1]));
    assign layer_4[621] = far_4_4701_1[0] ^ far_4_4701_1[1]; 
    wire [1:0] far_4_4702_0;    relay_conn far_4_4702_0_a(.in(layer_3[667]), .out(far_4_4702_0[0]));    relay_conn far_4_4702_0_b(.in(layer_3[712]), .out(far_4_4702_0[1]));
    assign layer_4[622] = ~far_4_4702_0[1]; 
    wire [1:0] far_4_4703_0;    relay_conn far_4_4703_0_a(.in(layer_3[893]), .out(far_4_4703_0[0]));    relay_conn far_4_4703_0_b(.in(layer_3[935]), .out(far_4_4703_0[1]));
    assign layer_4[623] = far_4_4703_0[0] & far_4_4703_0[1]; 
    wire [1:0] far_4_4704_0;    relay_conn far_4_4704_0_a(.in(layer_3[634]), .out(far_4_4704_0[0]));    relay_conn far_4_4704_0_b(.in(layer_3[512]), .out(far_4_4704_0[1]));
    wire [1:0] far_4_4704_1;    relay_conn far_4_4704_1_a(.in(far_4_4704_0[0]), .out(far_4_4704_1[0]));    relay_conn far_4_4704_1_b(.in(far_4_4704_0[1]), .out(far_4_4704_1[1]));
    wire [1:0] far_4_4704_2;    relay_conn far_4_4704_2_a(.in(far_4_4704_1[0]), .out(far_4_4704_2[0]));    relay_conn far_4_4704_2_b(.in(far_4_4704_1[1]), .out(far_4_4704_2[1]));
    assign layer_4[624] = ~far_4_4704_2[1]; 
    wire [1:0] far_4_4705_0;    relay_conn far_4_4705_0_a(.in(layer_3[125]), .out(far_4_4705_0[0]));    relay_conn far_4_4705_0_b(.in(layer_3[196]), .out(far_4_4705_0[1]));
    wire [1:0] far_4_4705_1;    relay_conn far_4_4705_1_a(.in(far_4_4705_0[0]), .out(far_4_4705_1[0]));    relay_conn far_4_4705_1_b(.in(far_4_4705_0[1]), .out(far_4_4705_1[1]));
    assign layer_4[625] = ~far_4_4705_1[1] | (far_4_4705_1[0] & far_4_4705_1[1]); 
    wire [1:0] far_4_4706_0;    relay_conn far_4_4706_0_a(.in(layer_3[922]), .out(far_4_4706_0[0]));    relay_conn far_4_4706_0_b(.in(layer_3[859]), .out(far_4_4706_0[1]));
    assign layer_4[626] = ~(far_4_4706_0[0] ^ far_4_4706_0[1]); 
    wire [1:0] far_4_4707_0;    relay_conn far_4_4707_0_a(.in(layer_3[486]), .out(far_4_4707_0[0]));    relay_conn far_4_4707_0_b(.in(layer_3[426]), .out(far_4_4707_0[1]));
    assign layer_4[627] = far_4_4707_0[1]; 
    wire [1:0] far_4_4708_0;    relay_conn far_4_4708_0_a(.in(layer_3[535]), .out(far_4_4708_0[0]));    relay_conn far_4_4708_0_b(.in(layer_3[433]), .out(far_4_4708_0[1]));
    wire [1:0] far_4_4708_1;    relay_conn far_4_4708_1_a(.in(far_4_4708_0[0]), .out(far_4_4708_1[0]));    relay_conn far_4_4708_1_b(.in(far_4_4708_0[1]), .out(far_4_4708_1[1]));
    wire [1:0] far_4_4708_2;    relay_conn far_4_4708_2_a(.in(far_4_4708_1[0]), .out(far_4_4708_2[0]));    relay_conn far_4_4708_2_b(.in(far_4_4708_1[1]), .out(far_4_4708_2[1]));
    assign layer_4[628] = far_4_4708_2[0] & far_4_4708_2[1]; 
    assign layer_4[629] = ~layer_3[887] | (layer_3[887] & layer_3[908]); 
    wire [1:0] far_4_4710_0;    relay_conn far_4_4710_0_a(.in(layer_3[882]), .out(far_4_4710_0[0]));    relay_conn far_4_4710_0_b(.in(layer_3[977]), .out(far_4_4710_0[1]));
    wire [1:0] far_4_4710_1;    relay_conn far_4_4710_1_a(.in(far_4_4710_0[0]), .out(far_4_4710_1[0]));    relay_conn far_4_4710_1_b(.in(far_4_4710_0[1]), .out(far_4_4710_1[1]));
    assign layer_4[630] = far_4_4710_1[0] | far_4_4710_1[1]; 
    assign layer_4[631] = layer_3[504] & layer_3[497]; 
    wire [1:0] far_4_4712_0;    relay_conn far_4_4712_0_a(.in(layer_3[511]), .out(far_4_4712_0[0]));    relay_conn far_4_4712_0_b(.in(layer_3[623]), .out(far_4_4712_0[1]));
    wire [1:0] far_4_4712_1;    relay_conn far_4_4712_1_a(.in(far_4_4712_0[0]), .out(far_4_4712_1[0]));    relay_conn far_4_4712_1_b(.in(far_4_4712_0[1]), .out(far_4_4712_1[1]));
    wire [1:0] far_4_4712_2;    relay_conn far_4_4712_2_a(.in(far_4_4712_1[0]), .out(far_4_4712_2[0]));    relay_conn far_4_4712_2_b(.in(far_4_4712_1[1]), .out(far_4_4712_2[1]));
    assign layer_4[632] = far_4_4712_2[1] & ~far_4_4712_2[0]; 
    wire [1:0] far_4_4713_0;    relay_conn far_4_4713_0_a(.in(layer_3[855]), .out(far_4_4713_0[0]));    relay_conn far_4_4713_0_b(.in(layer_3[774]), .out(far_4_4713_0[1]));
    wire [1:0] far_4_4713_1;    relay_conn far_4_4713_1_a(.in(far_4_4713_0[0]), .out(far_4_4713_1[0]));    relay_conn far_4_4713_1_b(.in(far_4_4713_0[1]), .out(far_4_4713_1[1]));
    assign layer_4[633] = far_4_4713_1[1] & ~far_4_4713_1[0]; 
    wire [1:0] far_4_4714_0;    relay_conn far_4_4714_0_a(.in(layer_3[72]), .out(far_4_4714_0[0]));    relay_conn far_4_4714_0_b(.in(layer_3[194]), .out(far_4_4714_0[1]));
    wire [1:0] far_4_4714_1;    relay_conn far_4_4714_1_a(.in(far_4_4714_0[0]), .out(far_4_4714_1[0]));    relay_conn far_4_4714_1_b(.in(far_4_4714_0[1]), .out(far_4_4714_1[1]));
    wire [1:0] far_4_4714_2;    relay_conn far_4_4714_2_a(.in(far_4_4714_1[0]), .out(far_4_4714_2[0]));    relay_conn far_4_4714_2_b(.in(far_4_4714_1[1]), .out(far_4_4714_2[1]));
    assign layer_4[634] = far_4_4714_2[0]; 
    wire [1:0] far_4_4715_0;    relay_conn far_4_4715_0_a(.in(layer_3[943]), .out(far_4_4715_0[0]));    relay_conn far_4_4715_0_b(.in(layer_3[837]), .out(far_4_4715_0[1]));
    wire [1:0] far_4_4715_1;    relay_conn far_4_4715_1_a(.in(far_4_4715_0[0]), .out(far_4_4715_1[0]));    relay_conn far_4_4715_1_b(.in(far_4_4715_0[1]), .out(far_4_4715_1[1]));
    wire [1:0] far_4_4715_2;    relay_conn far_4_4715_2_a(.in(far_4_4715_1[0]), .out(far_4_4715_2[0]));    relay_conn far_4_4715_2_b(.in(far_4_4715_1[1]), .out(far_4_4715_2[1]));
    assign layer_4[635] = ~far_4_4715_2[0] | (far_4_4715_2[0] & far_4_4715_2[1]); 
    wire [1:0] far_4_4716_0;    relay_conn far_4_4716_0_a(.in(layer_3[576]), .out(far_4_4716_0[0]));    relay_conn far_4_4716_0_b(.in(layer_3[676]), .out(far_4_4716_0[1]));
    wire [1:0] far_4_4716_1;    relay_conn far_4_4716_1_a(.in(far_4_4716_0[0]), .out(far_4_4716_1[0]));    relay_conn far_4_4716_1_b(.in(far_4_4716_0[1]), .out(far_4_4716_1[1]));
    wire [1:0] far_4_4716_2;    relay_conn far_4_4716_2_a(.in(far_4_4716_1[0]), .out(far_4_4716_2[0]));    relay_conn far_4_4716_2_b(.in(far_4_4716_1[1]), .out(far_4_4716_2[1]));
    assign layer_4[636] = ~far_4_4716_2[0] | (far_4_4716_2[0] & far_4_4716_2[1]); 
    wire [1:0] far_4_4717_0;    relay_conn far_4_4717_0_a(.in(layer_3[12]), .out(far_4_4717_0[0]));    relay_conn far_4_4717_0_b(.in(layer_3[49]), .out(far_4_4717_0[1]));
    assign layer_4[637] = far_4_4717_0[1]; 
    wire [1:0] far_4_4718_0;    relay_conn far_4_4718_0_a(.in(layer_3[649]), .out(far_4_4718_0[0]));    relay_conn far_4_4718_0_b(.in(layer_3[612]), .out(far_4_4718_0[1]));
    assign layer_4[638] = ~far_4_4718_0[0] | (far_4_4718_0[0] & far_4_4718_0[1]); 
    wire [1:0] far_4_4719_0;    relay_conn far_4_4719_0_a(.in(layer_3[622]), .out(far_4_4719_0[0]));    relay_conn far_4_4719_0_b(.in(layer_3[682]), .out(far_4_4719_0[1]));
    assign layer_4[639] = ~far_4_4719_0[0] | (far_4_4719_0[0] & far_4_4719_0[1]); 
    wire [1:0] far_4_4720_0;    relay_conn far_4_4720_0_a(.in(layer_3[363]), .out(far_4_4720_0[0]));    relay_conn far_4_4720_0_b(.in(layer_3[261]), .out(far_4_4720_0[1]));
    wire [1:0] far_4_4720_1;    relay_conn far_4_4720_1_a(.in(far_4_4720_0[0]), .out(far_4_4720_1[0]));    relay_conn far_4_4720_1_b(.in(far_4_4720_0[1]), .out(far_4_4720_1[1]));
    wire [1:0] far_4_4720_2;    relay_conn far_4_4720_2_a(.in(far_4_4720_1[0]), .out(far_4_4720_2[0]));    relay_conn far_4_4720_2_b(.in(far_4_4720_1[1]), .out(far_4_4720_2[1]));
    assign layer_4[640] = ~(far_4_4720_2[0] | far_4_4720_2[1]); 
    wire [1:0] far_4_4721_0;    relay_conn far_4_4721_0_a(.in(layer_3[478]), .out(far_4_4721_0[0]));    relay_conn far_4_4721_0_b(.in(layer_3[395]), .out(far_4_4721_0[1]));
    wire [1:0] far_4_4721_1;    relay_conn far_4_4721_1_a(.in(far_4_4721_0[0]), .out(far_4_4721_1[0]));    relay_conn far_4_4721_1_b(.in(far_4_4721_0[1]), .out(far_4_4721_1[1]));
    assign layer_4[641] = far_4_4721_1[0] | far_4_4721_1[1]; 
    wire [1:0] far_4_4722_0;    relay_conn far_4_4722_0_a(.in(layer_3[780]), .out(far_4_4722_0[0]));    relay_conn far_4_4722_0_b(.in(layer_3[726]), .out(far_4_4722_0[1]));
    assign layer_4[642] = ~far_4_4722_0[1]; 
    assign layer_4[643] = layer_3[695] | layer_3[664]; 
    wire [1:0] far_4_4724_0;    relay_conn far_4_4724_0_a(.in(layer_3[535]), .out(far_4_4724_0[0]));    relay_conn far_4_4724_0_b(.in(layer_3[586]), .out(far_4_4724_0[1]));
    assign layer_4[644] = far_4_4724_0[0] & ~far_4_4724_0[1]; 
    wire [1:0] far_4_4725_0;    relay_conn far_4_4725_0_a(.in(layer_3[797]), .out(far_4_4725_0[0]));    relay_conn far_4_4725_0_b(.in(layer_3[754]), .out(far_4_4725_0[1]));
    assign layer_4[645] = far_4_4725_0[0] & far_4_4725_0[1]; 
    assign layer_4[646] = ~layer_3[664] | (layer_3[664] & layer_3[633]); 
    assign layer_4[647] = layer_3[140] | layer_3[143]; 
    wire [1:0] far_4_4728_0;    relay_conn far_4_4728_0_a(.in(layer_3[329]), .out(far_4_4728_0[0]));    relay_conn far_4_4728_0_b(.in(layer_3[434]), .out(far_4_4728_0[1]));
    wire [1:0] far_4_4728_1;    relay_conn far_4_4728_1_a(.in(far_4_4728_0[0]), .out(far_4_4728_1[0]));    relay_conn far_4_4728_1_b(.in(far_4_4728_0[1]), .out(far_4_4728_1[1]));
    wire [1:0] far_4_4728_2;    relay_conn far_4_4728_2_a(.in(far_4_4728_1[0]), .out(far_4_4728_2[0]));    relay_conn far_4_4728_2_b(.in(far_4_4728_1[1]), .out(far_4_4728_2[1]));
    assign layer_4[648] = far_4_4728_2[1]; 
    wire [1:0] far_4_4729_0;    relay_conn far_4_4729_0_a(.in(layer_3[507]), .out(far_4_4729_0[0]));    relay_conn far_4_4729_0_b(.in(layer_3[598]), .out(far_4_4729_0[1]));
    wire [1:0] far_4_4729_1;    relay_conn far_4_4729_1_a(.in(far_4_4729_0[0]), .out(far_4_4729_1[0]));    relay_conn far_4_4729_1_b(.in(far_4_4729_0[1]), .out(far_4_4729_1[1]));
    assign layer_4[649] = ~(far_4_4729_1[0] | far_4_4729_1[1]); 
    wire [1:0] far_4_4730_0;    relay_conn far_4_4730_0_a(.in(layer_3[973]), .out(far_4_4730_0[0]));    relay_conn far_4_4730_0_b(.in(layer_3[903]), .out(far_4_4730_0[1]));
    wire [1:0] far_4_4730_1;    relay_conn far_4_4730_1_a(.in(far_4_4730_0[0]), .out(far_4_4730_1[0]));    relay_conn far_4_4730_1_b(.in(far_4_4730_0[1]), .out(far_4_4730_1[1]));
    assign layer_4[650] = ~far_4_4730_1[0]; 
    wire [1:0] far_4_4731_0;    relay_conn far_4_4731_0_a(.in(layer_3[402]), .out(far_4_4731_0[0]));    relay_conn far_4_4731_0_b(.in(layer_3[310]), .out(far_4_4731_0[1]));
    wire [1:0] far_4_4731_1;    relay_conn far_4_4731_1_a(.in(far_4_4731_0[0]), .out(far_4_4731_1[0]));    relay_conn far_4_4731_1_b(.in(far_4_4731_0[1]), .out(far_4_4731_1[1]));
    assign layer_4[651] = ~(far_4_4731_1[0] | far_4_4731_1[1]); 
    wire [1:0] far_4_4732_0;    relay_conn far_4_4732_0_a(.in(layer_3[179]), .out(far_4_4732_0[0]));    relay_conn far_4_4732_0_b(.in(layer_3[100]), .out(far_4_4732_0[1]));
    wire [1:0] far_4_4732_1;    relay_conn far_4_4732_1_a(.in(far_4_4732_0[0]), .out(far_4_4732_1[0]));    relay_conn far_4_4732_1_b(.in(far_4_4732_0[1]), .out(far_4_4732_1[1]));
    assign layer_4[652] = ~far_4_4732_1[1]; 
    wire [1:0] far_4_4733_0;    relay_conn far_4_4733_0_a(.in(layer_3[448]), .out(far_4_4733_0[0]));    relay_conn far_4_4733_0_b(.in(layer_3[546]), .out(far_4_4733_0[1]));
    wire [1:0] far_4_4733_1;    relay_conn far_4_4733_1_a(.in(far_4_4733_0[0]), .out(far_4_4733_1[0]));    relay_conn far_4_4733_1_b(.in(far_4_4733_0[1]), .out(far_4_4733_1[1]));
    wire [1:0] far_4_4733_2;    relay_conn far_4_4733_2_a(.in(far_4_4733_1[0]), .out(far_4_4733_2[0]));    relay_conn far_4_4733_2_b(.in(far_4_4733_1[1]), .out(far_4_4733_2[1]));
    assign layer_4[653] = ~(far_4_4733_2[0] | far_4_4733_2[1]); 
    wire [1:0] far_4_4734_0;    relay_conn far_4_4734_0_a(.in(layer_3[855]), .out(far_4_4734_0[0]));    relay_conn far_4_4734_0_b(.in(layer_3[909]), .out(far_4_4734_0[1]));
    assign layer_4[654] = far_4_4734_0[1] & ~far_4_4734_0[0]; 
    wire [1:0] far_4_4735_0;    relay_conn far_4_4735_0_a(.in(layer_3[811]), .out(far_4_4735_0[0]));    relay_conn far_4_4735_0_b(.in(layer_3[769]), .out(far_4_4735_0[1]));
    assign layer_4[655] = far_4_4735_0[0] & far_4_4735_0[1]; 
    wire [1:0] far_4_4736_0;    relay_conn far_4_4736_0_a(.in(layer_3[368]), .out(far_4_4736_0[0]));    relay_conn far_4_4736_0_b(.in(layer_3[303]), .out(far_4_4736_0[1]));
    wire [1:0] far_4_4736_1;    relay_conn far_4_4736_1_a(.in(far_4_4736_0[0]), .out(far_4_4736_1[0]));    relay_conn far_4_4736_1_b(.in(far_4_4736_0[1]), .out(far_4_4736_1[1]));
    assign layer_4[656] = ~(far_4_4736_1[0] & far_4_4736_1[1]); 
    wire [1:0] far_4_4737_0;    relay_conn far_4_4737_0_a(.in(layer_3[664]), .out(far_4_4737_0[0]));    relay_conn far_4_4737_0_b(.in(layer_3[599]), .out(far_4_4737_0[1]));
    wire [1:0] far_4_4737_1;    relay_conn far_4_4737_1_a(.in(far_4_4737_0[0]), .out(far_4_4737_1[0]));    relay_conn far_4_4737_1_b(.in(far_4_4737_0[1]), .out(far_4_4737_1[1]));
    assign layer_4[657] = ~far_4_4737_1[1] | (far_4_4737_1[0] & far_4_4737_1[1]); 
    assign layer_4[658] = layer_3[645] & ~layer_3[661]; 
    wire [1:0] far_4_4739_0;    relay_conn far_4_4739_0_a(.in(layer_3[310]), .out(far_4_4739_0[0]));    relay_conn far_4_4739_0_b(.in(layer_3[398]), .out(far_4_4739_0[1]));
    wire [1:0] far_4_4739_1;    relay_conn far_4_4739_1_a(.in(far_4_4739_0[0]), .out(far_4_4739_1[0]));    relay_conn far_4_4739_1_b(.in(far_4_4739_0[1]), .out(far_4_4739_1[1]));
    assign layer_4[659] = ~far_4_4739_1[0] | (far_4_4739_1[0] & far_4_4739_1[1]); 
    assign layer_4[660] = ~(layer_3[285] | layer_3[269]); 
    wire [1:0] far_4_4741_0;    relay_conn far_4_4741_0_a(.in(layer_3[116]), .out(far_4_4741_0[0]));    relay_conn far_4_4741_0_b(.in(layer_3[46]), .out(far_4_4741_0[1]));
    wire [1:0] far_4_4741_1;    relay_conn far_4_4741_1_a(.in(far_4_4741_0[0]), .out(far_4_4741_1[0]));    relay_conn far_4_4741_1_b(.in(far_4_4741_0[1]), .out(far_4_4741_1[1]));
    assign layer_4[661] = ~far_4_4741_1[1] | (far_4_4741_1[0] & far_4_4741_1[1]); 
    assign layer_4[662] = ~layer_3[195] | (layer_3[195] & layer_3[188]); 
    wire [1:0] far_4_4743_0;    relay_conn far_4_4743_0_a(.in(layer_3[302]), .out(far_4_4743_0[0]));    relay_conn far_4_4743_0_b(.in(layer_3[387]), .out(far_4_4743_0[1]));
    wire [1:0] far_4_4743_1;    relay_conn far_4_4743_1_a(.in(far_4_4743_0[0]), .out(far_4_4743_1[0]));    relay_conn far_4_4743_1_b(.in(far_4_4743_0[1]), .out(far_4_4743_1[1]));
    assign layer_4[663] = ~far_4_4743_1[0] | (far_4_4743_1[0] & far_4_4743_1[1]); 
    wire [1:0] far_4_4744_0;    relay_conn far_4_4744_0_a(.in(layer_3[58]), .out(far_4_4744_0[0]));    relay_conn far_4_4744_0_b(.in(layer_3[169]), .out(far_4_4744_0[1]));
    wire [1:0] far_4_4744_1;    relay_conn far_4_4744_1_a(.in(far_4_4744_0[0]), .out(far_4_4744_1[0]));    relay_conn far_4_4744_1_b(.in(far_4_4744_0[1]), .out(far_4_4744_1[1]));
    wire [1:0] far_4_4744_2;    relay_conn far_4_4744_2_a(.in(far_4_4744_1[0]), .out(far_4_4744_2[0]));    relay_conn far_4_4744_2_b(.in(far_4_4744_1[1]), .out(far_4_4744_2[1]));
    assign layer_4[664] = far_4_4744_2[0] ^ far_4_4744_2[1]; 
    wire [1:0] far_4_4745_0;    relay_conn far_4_4745_0_a(.in(layer_3[664]), .out(far_4_4745_0[0]));    relay_conn far_4_4745_0_b(.in(layer_3[721]), .out(far_4_4745_0[1]));
    assign layer_4[665] = far_4_4745_0[1]; 
    wire [1:0] far_4_4746_0;    relay_conn far_4_4746_0_a(.in(layer_3[697]), .out(far_4_4746_0[0]));    relay_conn far_4_4746_0_b(.in(layer_3[569]), .out(far_4_4746_0[1]));
    wire [1:0] far_4_4746_1;    relay_conn far_4_4746_1_a(.in(far_4_4746_0[0]), .out(far_4_4746_1[0]));    relay_conn far_4_4746_1_b(.in(far_4_4746_0[1]), .out(far_4_4746_1[1]));
    wire [1:0] far_4_4746_2;    relay_conn far_4_4746_2_a(.in(far_4_4746_1[0]), .out(far_4_4746_2[0]));    relay_conn far_4_4746_2_b(.in(far_4_4746_1[1]), .out(far_4_4746_2[1]));
    wire [1:0] far_4_4746_3;    relay_conn far_4_4746_3_a(.in(far_4_4746_2[0]), .out(far_4_4746_3[0]));    relay_conn far_4_4746_3_b(.in(far_4_4746_2[1]), .out(far_4_4746_3[1]));
    assign layer_4[666] = ~(far_4_4746_3[0] & far_4_4746_3[1]); 
    assign layer_4[667] = ~layer_3[492] | (layer_3[497] & layer_3[492]); 
    assign layer_4[668] = ~(layer_3[926] & layer_3[934]); 
    wire [1:0] far_4_4749_0;    relay_conn far_4_4749_0_a(.in(layer_3[466]), .out(far_4_4749_0[0]));    relay_conn far_4_4749_0_b(.in(layer_3[507]), .out(far_4_4749_0[1]));
    assign layer_4[669] = far_4_4749_0[0] | far_4_4749_0[1]; 
    assign layer_4[670] = layer_3[964]; 
    wire [1:0] far_4_4751_0;    relay_conn far_4_4751_0_a(.in(layer_3[718]), .out(far_4_4751_0[0]));    relay_conn far_4_4751_0_b(.in(layer_3[771]), .out(far_4_4751_0[1]));
    assign layer_4[671] = far_4_4751_0[0] & ~far_4_4751_0[1]; 
    assign layer_4[672] = layer_3[865]; 
    wire [1:0] far_4_4753_0;    relay_conn far_4_4753_0_a(.in(layer_3[674]), .out(far_4_4753_0[0]));    relay_conn far_4_4753_0_b(.in(layer_3[570]), .out(far_4_4753_0[1]));
    wire [1:0] far_4_4753_1;    relay_conn far_4_4753_1_a(.in(far_4_4753_0[0]), .out(far_4_4753_1[0]));    relay_conn far_4_4753_1_b(.in(far_4_4753_0[1]), .out(far_4_4753_1[1]));
    wire [1:0] far_4_4753_2;    relay_conn far_4_4753_2_a(.in(far_4_4753_1[0]), .out(far_4_4753_2[0]));    relay_conn far_4_4753_2_b(.in(far_4_4753_1[1]), .out(far_4_4753_2[1]));
    assign layer_4[673] = far_4_4753_2[0] | far_4_4753_2[1]; 
    wire [1:0] far_4_4754_0;    relay_conn far_4_4754_0_a(.in(layer_3[150]), .out(far_4_4754_0[0]));    relay_conn far_4_4754_0_b(.in(layer_3[48]), .out(far_4_4754_0[1]));
    wire [1:0] far_4_4754_1;    relay_conn far_4_4754_1_a(.in(far_4_4754_0[0]), .out(far_4_4754_1[0]));    relay_conn far_4_4754_1_b(.in(far_4_4754_0[1]), .out(far_4_4754_1[1]));
    wire [1:0] far_4_4754_2;    relay_conn far_4_4754_2_a(.in(far_4_4754_1[0]), .out(far_4_4754_2[0]));    relay_conn far_4_4754_2_b(.in(far_4_4754_1[1]), .out(far_4_4754_2[1]));
    assign layer_4[674] = ~(far_4_4754_2[0] & far_4_4754_2[1]); 
    wire [1:0] far_4_4755_0;    relay_conn far_4_4755_0_a(.in(layer_3[252]), .out(far_4_4755_0[0]));    relay_conn far_4_4755_0_b(.in(layer_3[192]), .out(far_4_4755_0[1]));
    assign layer_4[675] = ~far_4_4755_0[1]; 
    wire [1:0] far_4_4756_0;    relay_conn far_4_4756_0_a(.in(layer_3[281]), .out(far_4_4756_0[0]));    relay_conn far_4_4756_0_b(.in(layer_3[178]), .out(far_4_4756_0[1]));
    wire [1:0] far_4_4756_1;    relay_conn far_4_4756_1_a(.in(far_4_4756_0[0]), .out(far_4_4756_1[0]));    relay_conn far_4_4756_1_b(.in(far_4_4756_0[1]), .out(far_4_4756_1[1]));
    wire [1:0] far_4_4756_2;    relay_conn far_4_4756_2_a(.in(far_4_4756_1[0]), .out(far_4_4756_2[0]));    relay_conn far_4_4756_2_b(.in(far_4_4756_1[1]), .out(far_4_4756_2[1]));
    assign layer_4[676] = ~(far_4_4756_2[0] | far_4_4756_2[1]); 
    assign layer_4[677] = ~layer_3[666] | (layer_3[680] & layer_3[666]); 
    wire [1:0] far_4_4758_0;    relay_conn far_4_4758_0_a(.in(layer_3[563]), .out(far_4_4758_0[0]));    relay_conn far_4_4758_0_b(.in(layer_3[471]), .out(far_4_4758_0[1]));
    wire [1:0] far_4_4758_1;    relay_conn far_4_4758_1_a(.in(far_4_4758_0[0]), .out(far_4_4758_1[0]));    relay_conn far_4_4758_1_b(.in(far_4_4758_0[1]), .out(far_4_4758_1[1]));
    assign layer_4[678] = ~(far_4_4758_1[0] | far_4_4758_1[1]); 
    wire [1:0] far_4_4759_0;    relay_conn far_4_4759_0_a(.in(layer_3[322]), .out(far_4_4759_0[0]));    relay_conn far_4_4759_0_b(.in(layer_3[433]), .out(far_4_4759_0[1]));
    wire [1:0] far_4_4759_1;    relay_conn far_4_4759_1_a(.in(far_4_4759_0[0]), .out(far_4_4759_1[0]));    relay_conn far_4_4759_1_b(.in(far_4_4759_0[1]), .out(far_4_4759_1[1]));
    wire [1:0] far_4_4759_2;    relay_conn far_4_4759_2_a(.in(far_4_4759_1[0]), .out(far_4_4759_2[0]));    relay_conn far_4_4759_2_b(.in(far_4_4759_1[1]), .out(far_4_4759_2[1]));
    assign layer_4[679] = ~far_4_4759_2[1] | (far_4_4759_2[0] & far_4_4759_2[1]); 
    assign layer_4[680] = ~layer_3[972]; 
    assign layer_4[681] = layer_3[629] ^ layer_3[619]; 
    wire [1:0] far_4_4762_0;    relay_conn far_4_4762_0_a(.in(layer_3[625]), .out(far_4_4762_0[0]));    relay_conn far_4_4762_0_b(.in(layer_3[497]), .out(far_4_4762_0[1]));
    wire [1:0] far_4_4762_1;    relay_conn far_4_4762_1_a(.in(far_4_4762_0[0]), .out(far_4_4762_1[0]));    relay_conn far_4_4762_1_b(.in(far_4_4762_0[1]), .out(far_4_4762_1[1]));
    wire [1:0] far_4_4762_2;    relay_conn far_4_4762_2_a(.in(far_4_4762_1[0]), .out(far_4_4762_2[0]));    relay_conn far_4_4762_2_b(.in(far_4_4762_1[1]), .out(far_4_4762_2[1]));
    wire [1:0] far_4_4762_3;    relay_conn far_4_4762_3_a(.in(far_4_4762_2[0]), .out(far_4_4762_3[0]));    relay_conn far_4_4762_3_b(.in(far_4_4762_2[1]), .out(far_4_4762_3[1]));
    assign layer_4[682] = ~far_4_4762_3[1] | (far_4_4762_3[0] & far_4_4762_3[1]); 
    wire [1:0] far_4_4763_0;    relay_conn far_4_4763_0_a(.in(layer_3[466]), .out(far_4_4763_0[0]));    relay_conn far_4_4763_0_b(.in(layer_3[415]), .out(far_4_4763_0[1]));
    assign layer_4[683] = ~far_4_4763_0[0]; 
    wire [1:0] far_4_4764_0;    relay_conn far_4_4764_0_a(.in(layer_3[903]), .out(far_4_4764_0[0]));    relay_conn far_4_4764_0_b(.in(layer_3[943]), .out(far_4_4764_0[1]));
    assign layer_4[684] = far_4_4764_0[0]; 
    assign layer_4[685] = layer_3[769] & ~layer_3[741]; 
    wire [1:0] far_4_4766_0;    relay_conn far_4_4766_0_a(.in(layer_3[874]), .out(far_4_4766_0[0]));    relay_conn far_4_4766_0_b(.in(layer_3[931]), .out(far_4_4766_0[1]));
    assign layer_4[686] = ~(far_4_4766_0[0] | far_4_4766_0[1]); 
    wire [1:0] far_4_4767_0;    relay_conn far_4_4767_0_a(.in(layer_3[514]), .out(far_4_4767_0[0]));    relay_conn far_4_4767_0_b(.in(layer_3[576]), .out(far_4_4767_0[1]));
    assign layer_4[687] = ~far_4_4767_0[0]; 
    wire [1:0] far_4_4768_0;    relay_conn far_4_4768_0_a(.in(layer_3[142]), .out(far_4_4768_0[0]));    relay_conn far_4_4768_0_b(.in(layer_3[179]), .out(far_4_4768_0[1]));
    assign layer_4[688] = far_4_4768_0[0]; 
    wire [1:0] far_4_4769_0;    relay_conn far_4_4769_0_a(.in(layer_3[303]), .out(far_4_4769_0[0]));    relay_conn far_4_4769_0_b(.in(layer_3[189]), .out(far_4_4769_0[1]));
    wire [1:0] far_4_4769_1;    relay_conn far_4_4769_1_a(.in(far_4_4769_0[0]), .out(far_4_4769_1[0]));    relay_conn far_4_4769_1_b(.in(far_4_4769_0[1]), .out(far_4_4769_1[1]));
    wire [1:0] far_4_4769_2;    relay_conn far_4_4769_2_a(.in(far_4_4769_1[0]), .out(far_4_4769_2[0]));    relay_conn far_4_4769_2_b(.in(far_4_4769_1[1]), .out(far_4_4769_2[1]));
    assign layer_4[689] = far_4_4769_2[1]; 
    wire [1:0] far_4_4770_0;    relay_conn far_4_4770_0_a(.in(layer_3[414]), .out(far_4_4770_0[0]));    relay_conn far_4_4770_0_b(.in(layer_3[470]), .out(far_4_4770_0[1]));
    assign layer_4[690] = ~far_4_4770_0[0]; 
    wire [1:0] far_4_4771_0;    relay_conn far_4_4771_0_a(.in(layer_3[102]), .out(far_4_4771_0[0]));    relay_conn far_4_4771_0_b(.in(layer_3[178]), .out(far_4_4771_0[1]));
    wire [1:0] far_4_4771_1;    relay_conn far_4_4771_1_a(.in(far_4_4771_0[0]), .out(far_4_4771_1[0]));    relay_conn far_4_4771_1_b(.in(far_4_4771_0[1]), .out(far_4_4771_1[1]));
    assign layer_4[691] = ~(far_4_4771_1[0] & far_4_4771_1[1]); 
    wire [1:0] far_4_4772_0;    relay_conn far_4_4772_0_a(.in(layer_3[527]), .out(far_4_4772_0[0]));    relay_conn far_4_4772_0_b(.in(layer_3[456]), .out(far_4_4772_0[1]));
    wire [1:0] far_4_4772_1;    relay_conn far_4_4772_1_a(.in(far_4_4772_0[0]), .out(far_4_4772_1[0]));    relay_conn far_4_4772_1_b(.in(far_4_4772_0[1]), .out(far_4_4772_1[1]));
    assign layer_4[692] = ~far_4_4772_1[1] | (far_4_4772_1[0] & far_4_4772_1[1]); 
    wire [1:0] far_4_4773_0;    relay_conn far_4_4773_0_a(.in(layer_3[424]), .out(far_4_4773_0[0]));    relay_conn far_4_4773_0_b(.in(layer_3[478]), .out(far_4_4773_0[1]));
    assign layer_4[693] = ~(far_4_4773_0[0] & far_4_4773_0[1]); 
    wire [1:0] far_4_4774_0;    relay_conn far_4_4774_0_a(.in(layer_3[813]), .out(far_4_4774_0[0]));    relay_conn far_4_4774_0_b(.in(layer_3[880]), .out(far_4_4774_0[1]));
    wire [1:0] far_4_4774_1;    relay_conn far_4_4774_1_a(.in(far_4_4774_0[0]), .out(far_4_4774_1[0]));    relay_conn far_4_4774_1_b(.in(far_4_4774_0[1]), .out(far_4_4774_1[1]));
    assign layer_4[694] = ~(far_4_4774_1[0] & far_4_4774_1[1]); 
    wire [1:0] far_4_4775_0;    relay_conn far_4_4775_0_a(.in(layer_3[274]), .out(far_4_4775_0[0]));    relay_conn far_4_4775_0_b(.in(layer_3[386]), .out(far_4_4775_0[1]));
    wire [1:0] far_4_4775_1;    relay_conn far_4_4775_1_a(.in(far_4_4775_0[0]), .out(far_4_4775_1[0]));    relay_conn far_4_4775_1_b(.in(far_4_4775_0[1]), .out(far_4_4775_1[1]));
    wire [1:0] far_4_4775_2;    relay_conn far_4_4775_2_a(.in(far_4_4775_1[0]), .out(far_4_4775_2[0]));    relay_conn far_4_4775_2_b(.in(far_4_4775_1[1]), .out(far_4_4775_2[1]));
    assign layer_4[695] = far_4_4775_2[0] & far_4_4775_2[1]; 
    wire [1:0] far_4_4776_0;    relay_conn far_4_4776_0_a(.in(layer_3[61]), .out(far_4_4776_0[0]));    relay_conn far_4_4776_0_b(.in(layer_3[102]), .out(far_4_4776_0[1]));
    assign layer_4[696] = ~far_4_4776_0[1]; 
    wire [1:0] far_4_4777_0;    relay_conn far_4_4777_0_a(.in(layer_3[629]), .out(far_4_4777_0[0]));    relay_conn far_4_4777_0_b(.in(layer_3[707]), .out(far_4_4777_0[1]));
    wire [1:0] far_4_4777_1;    relay_conn far_4_4777_1_a(.in(far_4_4777_0[0]), .out(far_4_4777_1[0]));    relay_conn far_4_4777_1_b(.in(far_4_4777_0[1]), .out(far_4_4777_1[1]));
    assign layer_4[697] = far_4_4777_1[1] & ~far_4_4777_1[0]; 
    wire [1:0] far_4_4778_0;    relay_conn far_4_4778_0_a(.in(layer_3[299]), .out(far_4_4778_0[0]));    relay_conn far_4_4778_0_b(.in(layer_3[179]), .out(far_4_4778_0[1]));
    wire [1:0] far_4_4778_1;    relay_conn far_4_4778_1_a(.in(far_4_4778_0[0]), .out(far_4_4778_1[0]));    relay_conn far_4_4778_1_b(.in(far_4_4778_0[1]), .out(far_4_4778_1[1]));
    wire [1:0] far_4_4778_2;    relay_conn far_4_4778_2_a(.in(far_4_4778_1[0]), .out(far_4_4778_2[0]));    relay_conn far_4_4778_2_b(.in(far_4_4778_1[1]), .out(far_4_4778_2[1]));
    assign layer_4[698] = ~far_4_4778_2[0] | (far_4_4778_2[0] & far_4_4778_2[1]); 
    wire [1:0] far_4_4779_0;    relay_conn far_4_4779_0_a(.in(layer_3[853]), .out(far_4_4779_0[0]));    relay_conn far_4_4779_0_b(.in(layer_3[900]), .out(far_4_4779_0[1]));
    assign layer_4[699] = far_4_4779_0[0] & far_4_4779_0[1]; 
    assign layer_4[700] = ~(layer_3[457] | layer_3[439]); 
    wire [1:0] far_4_4781_0;    relay_conn far_4_4781_0_a(.in(layer_3[368]), .out(far_4_4781_0[0]));    relay_conn far_4_4781_0_b(.in(layer_3[424]), .out(far_4_4781_0[1]));
    assign layer_4[701] = ~(far_4_4781_0[0] ^ far_4_4781_0[1]); 
    wire [1:0] far_4_4782_0;    relay_conn far_4_4782_0_a(.in(layer_3[179]), .out(far_4_4782_0[0]));    relay_conn far_4_4782_0_b(.in(layer_3[212]), .out(far_4_4782_0[1]));
    assign layer_4[702] = far_4_4782_0[0] & far_4_4782_0[1]; 
    assign layer_4[703] = ~layer_3[189]; 
    wire [1:0] far_4_4784_0;    relay_conn far_4_4784_0_a(.in(layer_3[251]), .out(far_4_4784_0[0]));    relay_conn far_4_4784_0_b(.in(layer_3[140]), .out(far_4_4784_0[1]));
    wire [1:0] far_4_4784_1;    relay_conn far_4_4784_1_a(.in(far_4_4784_0[0]), .out(far_4_4784_1[0]));    relay_conn far_4_4784_1_b(.in(far_4_4784_0[1]), .out(far_4_4784_1[1]));
    wire [1:0] far_4_4784_2;    relay_conn far_4_4784_2_a(.in(far_4_4784_1[0]), .out(far_4_4784_2[0]));    relay_conn far_4_4784_2_b(.in(far_4_4784_1[1]), .out(far_4_4784_2[1]));
    assign layer_4[704] = ~far_4_4784_2[0] | (far_4_4784_2[0] & far_4_4784_2[1]); 
    wire [1:0] far_4_4785_0;    relay_conn far_4_4785_0_a(.in(layer_3[235]), .out(far_4_4785_0[0]));    relay_conn far_4_4785_0_b(.in(layer_3[169]), .out(far_4_4785_0[1]));
    wire [1:0] far_4_4785_1;    relay_conn far_4_4785_1_a(.in(far_4_4785_0[0]), .out(far_4_4785_1[0]));    relay_conn far_4_4785_1_b(.in(far_4_4785_0[1]), .out(far_4_4785_1[1]));
    assign layer_4[705] = ~(far_4_4785_1[0] | far_4_4785_1[1]); 
    wire [1:0] far_4_4786_0;    relay_conn far_4_4786_0_a(.in(layer_3[531]), .out(far_4_4786_0[0]));    relay_conn far_4_4786_0_b(.in(layer_3[416]), .out(far_4_4786_0[1]));
    wire [1:0] far_4_4786_1;    relay_conn far_4_4786_1_a(.in(far_4_4786_0[0]), .out(far_4_4786_1[0]));    relay_conn far_4_4786_1_b(.in(far_4_4786_0[1]), .out(far_4_4786_1[1]));
    wire [1:0] far_4_4786_2;    relay_conn far_4_4786_2_a(.in(far_4_4786_1[0]), .out(far_4_4786_2[0]));    relay_conn far_4_4786_2_b(.in(far_4_4786_1[1]), .out(far_4_4786_2[1]));
    assign layer_4[706] = far_4_4786_2[0]; 
    wire [1:0] far_4_4787_0;    relay_conn far_4_4787_0_a(.in(layer_3[771]), .out(far_4_4787_0[0]));    relay_conn far_4_4787_0_b(.in(layer_3[649]), .out(far_4_4787_0[1]));
    wire [1:0] far_4_4787_1;    relay_conn far_4_4787_1_a(.in(far_4_4787_0[0]), .out(far_4_4787_1[0]));    relay_conn far_4_4787_1_b(.in(far_4_4787_0[1]), .out(far_4_4787_1[1]));
    wire [1:0] far_4_4787_2;    relay_conn far_4_4787_2_a(.in(far_4_4787_1[0]), .out(far_4_4787_2[0]));    relay_conn far_4_4787_2_b(.in(far_4_4787_1[1]), .out(far_4_4787_2[1]));
    assign layer_4[707] = ~far_4_4787_2[0] | (far_4_4787_2[0] & far_4_4787_2[1]); 
    assign layer_4[708] = ~(layer_3[164] ^ layer_3[140]); 
    wire [1:0] far_4_4789_0;    relay_conn far_4_4789_0_a(.in(layer_3[660]), .out(far_4_4789_0[0]));    relay_conn far_4_4789_0_b(.in(layer_3[556]), .out(far_4_4789_0[1]));
    wire [1:0] far_4_4789_1;    relay_conn far_4_4789_1_a(.in(far_4_4789_0[0]), .out(far_4_4789_1[0]));    relay_conn far_4_4789_1_b(.in(far_4_4789_0[1]), .out(far_4_4789_1[1]));
    wire [1:0] far_4_4789_2;    relay_conn far_4_4789_2_a(.in(far_4_4789_1[0]), .out(far_4_4789_2[0]));    relay_conn far_4_4789_2_b(.in(far_4_4789_1[1]), .out(far_4_4789_2[1]));
    assign layer_4[709] = ~(far_4_4789_2[0] & far_4_4789_2[1]); 
    wire [1:0] far_4_4790_0;    relay_conn far_4_4790_0_a(.in(layer_3[196]), .out(far_4_4790_0[0]));    relay_conn far_4_4790_0_b(.in(layer_3[100]), .out(far_4_4790_0[1]));
    wire [1:0] far_4_4790_1;    relay_conn far_4_4790_1_a(.in(far_4_4790_0[0]), .out(far_4_4790_1[0]));    relay_conn far_4_4790_1_b(.in(far_4_4790_0[1]), .out(far_4_4790_1[1]));
    wire [1:0] far_4_4790_2;    relay_conn far_4_4790_2_a(.in(far_4_4790_1[0]), .out(far_4_4790_2[0]));    relay_conn far_4_4790_2_b(.in(far_4_4790_1[1]), .out(far_4_4790_2[1]));
    assign layer_4[710] = ~far_4_4790_2[0] | (far_4_4790_2[0] & far_4_4790_2[1]); 
    wire [1:0] far_4_4791_0;    relay_conn far_4_4791_0_a(.in(layer_3[50]), .out(far_4_4791_0[0]));    relay_conn far_4_4791_0_b(.in(layer_3[158]), .out(far_4_4791_0[1]));
    wire [1:0] far_4_4791_1;    relay_conn far_4_4791_1_a(.in(far_4_4791_0[0]), .out(far_4_4791_1[0]));    relay_conn far_4_4791_1_b(.in(far_4_4791_0[1]), .out(far_4_4791_1[1]));
    wire [1:0] far_4_4791_2;    relay_conn far_4_4791_2_a(.in(far_4_4791_1[0]), .out(far_4_4791_2[0]));    relay_conn far_4_4791_2_b(.in(far_4_4791_1[1]), .out(far_4_4791_2[1]));
    assign layer_4[711] = far_4_4791_2[1]; 
    wire [1:0] far_4_4792_0;    relay_conn far_4_4792_0_a(.in(layer_3[742]), .out(far_4_4792_0[0]));    relay_conn far_4_4792_0_b(.in(layer_3[654]), .out(far_4_4792_0[1]));
    wire [1:0] far_4_4792_1;    relay_conn far_4_4792_1_a(.in(far_4_4792_0[0]), .out(far_4_4792_1[0]));    relay_conn far_4_4792_1_b(.in(far_4_4792_0[1]), .out(far_4_4792_1[1]));
    assign layer_4[712] = far_4_4792_1[1]; 
    wire [1:0] far_4_4793_0;    relay_conn far_4_4793_0_a(.in(layer_3[973]), .out(far_4_4793_0[0]));    relay_conn far_4_4793_0_b(.in(layer_3[1018]), .out(far_4_4793_0[1]));
    assign layer_4[713] = far_4_4793_0[0] | far_4_4793_0[1]; 
    wire [1:0] far_4_4794_0;    relay_conn far_4_4794_0_a(.in(layer_3[675]), .out(far_4_4794_0[0]));    relay_conn far_4_4794_0_b(.in(layer_3[620]), .out(far_4_4794_0[1]));
    assign layer_4[714] = ~far_4_4794_0[0] | (far_4_4794_0[0] & far_4_4794_0[1]); 
    wire [1:0] far_4_4795_0;    relay_conn far_4_4795_0_a(.in(layer_3[258]), .out(far_4_4795_0[0]));    relay_conn far_4_4795_0_b(.in(layer_3[364]), .out(far_4_4795_0[1]));
    wire [1:0] far_4_4795_1;    relay_conn far_4_4795_1_a(.in(far_4_4795_0[0]), .out(far_4_4795_1[0]));    relay_conn far_4_4795_1_b(.in(far_4_4795_0[1]), .out(far_4_4795_1[1]));
    wire [1:0] far_4_4795_2;    relay_conn far_4_4795_2_a(.in(far_4_4795_1[0]), .out(far_4_4795_2[0]));    relay_conn far_4_4795_2_b(.in(far_4_4795_1[1]), .out(far_4_4795_2[1]));
    assign layer_4[715] = ~(far_4_4795_2[0] ^ far_4_4795_2[1]); 
    wire [1:0] far_4_4796_0;    relay_conn far_4_4796_0_a(.in(layer_3[142]), .out(far_4_4796_0[0]));    relay_conn far_4_4796_0_b(.in(layer_3[232]), .out(far_4_4796_0[1]));
    wire [1:0] far_4_4796_1;    relay_conn far_4_4796_1_a(.in(far_4_4796_0[0]), .out(far_4_4796_1[0]));    relay_conn far_4_4796_1_b(.in(far_4_4796_0[1]), .out(far_4_4796_1[1]));
    assign layer_4[716] = ~far_4_4796_1[0]; 
    wire [1:0] far_4_4797_0;    relay_conn far_4_4797_0_a(.in(layer_3[25]), .out(far_4_4797_0[0]));    relay_conn far_4_4797_0_b(.in(layer_3[127]), .out(far_4_4797_0[1]));
    wire [1:0] far_4_4797_1;    relay_conn far_4_4797_1_a(.in(far_4_4797_0[0]), .out(far_4_4797_1[0]));    relay_conn far_4_4797_1_b(.in(far_4_4797_0[1]), .out(far_4_4797_1[1]));
    wire [1:0] far_4_4797_2;    relay_conn far_4_4797_2_a(.in(far_4_4797_1[0]), .out(far_4_4797_2[0]));    relay_conn far_4_4797_2_b(.in(far_4_4797_1[1]), .out(far_4_4797_2[1]));
    assign layer_4[717] = far_4_4797_2[0] & far_4_4797_2[1]; 
    assign layer_4[718] = ~layer_3[700] | (layer_3[727] & layer_3[700]); 
    wire [1:0] far_4_4799_0;    relay_conn far_4_4799_0_a(.in(layer_3[582]), .out(far_4_4799_0[0]));    relay_conn far_4_4799_0_b(.in(layer_3[645]), .out(far_4_4799_0[1]));
    assign layer_4[719] = ~(far_4_4799_0[0] & far_4_4799_0[1]); 
    wire [1:0] far_4_4800_0;    relay_conn far_4_4800_0_a(.in(layer_3[0]), .out(far_4_4800_0[0]));    relay_conn far_4_4800_0_b(.in(layer_3[75]), .out(far_4_4800_0[1]));
    wire [1:0] far_4_4800_1;    relay_conn far_4_4800_1_a(.in(far_4_4800_0[0]), .out(far_4_4800_1[0]));    relay_conn far_4_4800_1_b(.in(far_4_4800_0[1]), .out(far_4_4800_1[1]));
    assign layer_4[720] = far_4_4800_1[0] & far_4_4800_1[1]; 
    wire [1:0] far_4_4801_0;    relay_conn far_4_4801_0_a(.in(layer_3[312]), .out(far_4_4801_0[0]));    relay_conn far_4_4801_0_b(.in(layer_3[420]), .out(far_4_4801_0[1]));
    wire [1:0] far_4_4801_1;    relay_conn far_4_4801_1_a(.in(far_4_4801_0[0]), .out(far_4_4801_1[0]));    relay_conn far_4_4801_1_b(.in(far_4_4801_0[1]), .out(far_4_4801_1[1]));
    wire [1:0] far_4_4801_2;    relay_conn far_4_4801_2_a(.in(far_4_4801_1[0]), .out(far_4_4801_2[0]));    relay_conn far_4_4801_2_b(.in(far_4_4801_1[1]), .out(far_4_4801_2[1]));
    assign layer_4[721] = far_4_4801_2[0] & ~far_4_4801_2[1]; 
    assign layer_4[722] = layer_3[878] ^ layer_3[909]; 
    wire [1:0] far_4_4803_0;    relay_conn far_4_4803_0_a(.in(layer_3[834]), .out(far_4_4803_0[0]));    relay_conn far_4_4803_0_b(.in(layer_3[941]), .out(far_4_4803_0[1]));
    wire [1:0] far_4_4803_1;    relay_conn far_4_4803_1_a(.in(far_4_4803_0[0]), .out(far_4_4803_1[0]));    relay_conn far_4_4803_1_b(.in(far_4_4803_0[1]), .out(far_4_4803_1[1]));
    wire [1:0] far_4_4803_2;    relay_conn far_4_4803_2_a(.in(far_4_4803_1[0]), .out(far_4_4803_2[0]));    relay_conn far_4_4803_2_b(.in(far_4_4803_1[1]), .out(far_4_4803_2[1]));
    assign layer_4[723] = ~(far_4_4803_2[0] & far_4_4803_2[1]); 
    wire [1:0] far_4_4804_0;    relay_conn far_4_4804_0_a(.in(layer_3[112]), .out(far_4_4804_0[0]));    relay_conn far_4_4804_0_b(.in(layer_3[195]), .out(far_4_4804_0[1]));
    wire [1:0] far_4_4804_1;    relay_conn far_4_4804_1_a(.in(far_4_4804_0[0]), .out(far_4_4804_1[0]));    relay_conn far_4_4804_1_b(.in(far_4_4804_0[1]), .out(far_4_4804_1[1]));
    assign layer_4[724] = ~far_4_4804_1[0] | (far_4_4804_1[0] & far_4_4804_1[1]); 
    wire [1:0] far_4_4805_0;    relay_conn far_4_4805_0_a(.in(layer_3[486]), .out(far_4_4805_0[0]));    relay_conn far_4_4805_0_b(.in(layer_3[401]), .out(far_4_4805_0[1]));
    wire [1:0] far_4_4805_1;    relay_conn far_4_4805_1_a(.in(far_4_4805_0[0]), .out(far_4_4805_1[0]));    relay_conn far_4_4805_1_b(.in(far_4_4805_0[1]), .out(far_4_4805_1[1]));
    assign layer_4[725] = ~(far_4_4805_1[0] | far_4_4805_1[1]); 
    wire [1:0] far_4_4806_0;    relay_conn far_4_4806_0_a(.in(layer_3[568]), .out(far_4_4806_0[0]));    relay_conn far_4_4806_0_b(.in(layer_3[648]), .out(far_4_4806_0[1]));
    wire [1:0] far_4_4806_1;    relay_conn far_4_4806_1_a(.in(far_4_4806_0[0]), .out(far_4_4806_1[0]));    relay_conn far_4_4806_1_b(.in(far_4_4806_0[1]), .out(far_4_4806_1[1]));
    assign layer_4[726] = far_4_4806_1[1] & ~far_4_4806_1[0]; 
    assign layer_4[727] = ~(layer_3[782] ^ layer_3[778]); 
    wire [1:0] far_4_4808_0;    relay_conn far_4_4808_0_a(.in(layer_3[176]), .out(far_4_4808_0[0]));    relay_conn far_4_4808_0_b(.in(layer_3[135]), .out(far_4_4808_0[1]));
    assign layer_4[728] = ~far_4_4808_0[1] | (far_4_4808_0[0] & far_4_4808_0[1]); 
    wire [1:0] far_4_4809_0;    relay_conn far_4_4809_0_a(.in(layer_3[944]), .out(far_4_4809_0[0]));    relay_conn far_4_4809_0_b(.in(layer_3[823]), .out(far_4_4809_0[1]));
    wire [1:0] far_4_4809_1;    relay_conn far_4_4809_1_a(.in(far_4_4809_0[0]), .out(far_4_4809_1[0]));    relay_conn far_4_4809_1_b(.in(far_4_4809_0[1]), .out(far_4_4809_1[1]));
    wire [1:0] far_4_4809_2;    relay_conn far_4_4809_2_a(.in(far_4_4809_1[0]), .out(far_4_4809_2[0]));    relay_conn far_4_4809_2_b(.in(far_4_4809_1[1]), .out(far_4_4809_2[1]));
    assign layer_4[729] = far_4_4809_2[1]; 
    assign layer_4[730] = layer_3[981] & layer_3[982]; 
    assign layer_4[731] = layer_3[212]; 
    wire [1:0] far_4_4812_0;    relay_conn far_4_4812_0_a(.in(layer_3[65]), .out(far_4_4812_0[0]));    relay_conn far_4_4812_0_b(.in(layer_3[179]), .out(far_4_4812_0[1]));
    wire [1:0] far_4_4812_1;    relay_conn far_4_4812_1_a(.in(far_4_4812_0[0]), .out(far_4_4812_1[0]));    relay_conn far_4_4812_1_b(.in(far_4_4812_0[1]), .out(far_4_4812_1[1]));
    wire [1:0] far_4_4812_2;    relay_conn far_4_4812_2_a(.in(far_4_4812_1[0]), .out(far_4_4812_2[0]));    relay_conn far_4_4812_2_b(.in(far_4_4812_1[1]), .out(far_4_4812_2[1]));
    assign layer_4[732] = ~(far_4_4812_2[0] & far_4_4812_2[1]); 
    wire [1:0] far_4_4813_0;    relay_conn far_4_4813_0_a(.in(layer_3[985]), .out(far_4_4813_0[0]));    relay_conn far_4_4813_0_b(.in(layer_3[884]), .out(far_4_4813_0[1]));
    wire [1:0] far_4_4813_1;    relay_conn far_4_4813_1_a(.in(far_4_4813_0[0]), .out(far_4_4813_1[0]));    relay_conn far_4_4813_1_b(.in(far_4_4813_0[1]), .out(far_4_4813_1[1]));
    wire [1:0] far_4_4813_2;    relay_conn far_4_4813_2_a(.in(far_4_4813_1[0]), .out(far_4_4813_2[0]));    relay_conn far_4_4813_2_b(.in(far_4_4813_1[1]), .out(far_4_4813_2[1]));
    assign layer_4[733] = ~(far_4_4813_2[0] & far_4_4813_2[1]); 
    wire [1:0] far_4_4814_0;    relay_conn far_4_4814_0_a(.in(layer_3[128]), .out(far_4_4814_0[0]));    relay_conn far_4_4814_0_b(.in(layer_3[80]), .out(far_4_4814_0[1]));
    assign layer_4[734] = ~(far_4_4814_0[0] ^ far_4_4814_0[1]); 
    assign layer_4[735] = ~(layer_3[47] & layer_3[35]); 
    wire [1:0] far_4_4816_0;    relay_conn far_4_4816_0_a(.in(layer_3[416]), .out(far_4_4816_0[0]));    relay_conn far_4_4816_0_b(.in(layer_3[458]), .out(far_4_4816_0[1]));
    assign layer_4[736] = ~far_4_4816_0[1]; 
    wire [1:0] far_4_4817_0;    relay_conn far_4_4817_0_a(.in(layer_3[834]), .out(far_4_4817_0[0]));    relay_conn far_4_4817_0_b(.in(layer_3[893]), .out(far_4_4817_0[1]));
    assign layer_4[737] = far_4_4817_0[0]; 
    assign layer_4[738] = ~(layer_3[106] & layer_3[135]); 
    assign layer_4[739] = layer_3[879]; 
    assign layer_4[740] = ~(layer_3[807] | layer_3[818]); 
    assign layer_4[741] = layer_3[762]; 
    assign layer_4[742] = ~(layer_3[321] & layer_3[307]); 
    wire [1:0] far_4_4823_0;    relay_conn far_4_4823_0_a(.in(layer_3[943]), .out(far_4_4823_0[0]));    relay_conn far_4_4823_0_b(.in(layer_3[991]), .out(far_4_4823_0[1]));
    assign layer_4[743] = ~far_4_4823_0[0]; 
    wire [1:0] far_4_4824_0;    relay_conn far_4_4824_0_a(.in(layer_3[442]), .out(far_4_4824_0[0]));    relay_conn far_4_4824_0_b(.in(layer_3[323]), .out(far_4_4824_0[1]));
    wire [1:0] far_4_4824_1;    relay_conn far_4_4824_1_a(.in(far_4_4824_0[0]), .out(far_4_4824_1[0]));    relay_conn far_4_4824_1_b(.in(far_4_4824_0[1]), .out(far_4_4824_1[1]));
    wire [1:0] far_4_4824_2;    relay_conn far_4_4824_2_a(.in(far_4_4824_1[0]), .out(far_4_4824_2[0]));    relay_conn far_4_4824_2_b(.in(far_4_4824_1[1]), .out(far_4_4824_2[1]));
    assign layer_4[744] = far_4_4824_2[0] | far_4_4824_2[1]; 
    wire [1:0] far_4_4825_0;    relay_conn far_4_4825_0_a(.in(layer_3[477]), .out(far_4_4825_0[0]));    relay_conn far_4_4825_0_b(.in(layer_3[429]), .out(far_4_4825_0[1]));
    assign layer_4[745] = ~far_4_4825_0[0] | (far_4_4825_0[0] & far_4_4825_0[1]); 
    wire [1:0] far_4_4826_0;    relay_conn far_4_4826_0_a(.in(layer_3[248]), .out(far_4_4826_0[0]));    relay_conn far_4_4826_0_b(.in(layer_3[368]), .out(far_4_4826_0[1]));
    wire [1:0] far_4_4826_1;    relay_conn far_4_4826_1_a(.in(far_4_4826_0[0]), .out(far_4_4826_1[0]));    relay_conn far_4_4826_1_b(.in(far_4_4826_0[1]), .out(far_4_4826_1[1]));
    wire [1:0] far_4_4826_2;    relay_conn far_4_4826_2_a(.in(far_4_4826_1[0]), .out(far_4_4826_2[0]));    relay_conn far_4_4826_2_b(.in(far_4_4826_1[1]), .out(far_4_4826_2[1]));
    assign layer_4[746] = far_4_4826_2[0]; 
    wire [1:0] far_4_4827_0;    relay_conn far_4_4827_0_a(.in(layer_3[768]), .out(far_4_4827_0[0]));    relay_conn far_4_4827_0_b(.in(layer_3[801]), .out(far_4_4827_0[1]));
    assign layer_4[747] = ~(far_4_4827_0[0] & far_4_4827_0[1]); 
    wire [1:0] far_4_4828_0;    relay_conn far_4_4828_0_a(.in(layer_3[232]), .out(far_4_4828_0[0]));    relay_conn far_4_4828_0_b(.in(layer_3[352]), .out(far_4_4828_0[1]));
    wire [1:0] far_4_4828_1;    relay_conn far_4_4828_1_a(.in(far_4_4828_0[0]), .out(far_4_4828_1[0]));    relay_conn far_4_4828_1_b(.in(far_4_4828_0[1]), .out(far_4_4828_1[1]));
    wire [1:0] far_4_4828_2;    relay_conn far_4_4828_2_a(.in(far_4_4828_1[0]), .out(far_4_4828_2[0]));    relay_conn far_4_4828_2_b(.in(far_4_4828_1[1]), .out(far_4_4828_2[1]));
    assign layer_4[748] = far_4_4828_2[1]; 
    assign layer_4[749] = layer_3[51] & layer_3[72]; 
    wire [1:0] far_4_4830_0;    relay_conn far_4_4830_0_a(.in(layer_3[717]), .out(far_4_4830_0[0]));    relay_conn far_4_4830_0_b(.in(layer_3[816]), .out(far_4_4830_0[1]));
    wire [1:0] far_4_4830_1;    relay_conn far_4_4830_1_a(.in(far_4_4830_0[0]), .out(far_4_4830_1[0]));    relay_conn far_4_4830_1_b(.in(far_4_4830_0[1]), .out(far_4_4830_1[1]));
    wire [1:0] far_4_4830_2;    relay_conn far_4_4830_2_a(.in(far_4_4830_1[0]), .out(far_4_4830_2[0]));    relay_conn far_4_4830_2_b(.in(far_4_4830_1[1]), .out(far_4_4830_2[1]));
    assign layer_4[750] = far_4_4830_2[0] & ~far_4_4830_2[1]; 
    wire [1:0] far_4_4831_0;    relay_conn far_4_4831_0_a(.in(layer_3[981]), .out(far_4_4831_0[0]));    relay_conn far_4_4831_0_b(.in(layer_3[861]), .out(far_4_4831_0[1]));
    wire [1:0] far_4_4831_1;    relay_conn far_4_4831_1_a(.in(far_4_4831_0[0]), .out(far_4_4831_1[0]));    relay_conn far_4_4831_1_b(.in(far_4_4831_0[1]), .out(far_4_4831_1[1]));
    wire [1:0] far_4_4831_2;    relay_conn far_4_4831_2_a(.in(far_4_4831_1[0]), .out(far_4_4831_2[0]));    relay_conn far_4_4831_2_b(.in(far_4_4831_1[1]), .out(far_4_4831_2[1]));
    assign layer_4[751] = ~(far_4_4831_2[0] ^ far_4_4831_2[1]); 
    assign layer_4[752] = ~layer_3[512] | (layer_3[488] & layer_3[512]); 
    assign layer_4[753] = ~layer_3[152]; 
    wire [1:0] far_4_4834_0;    relay_conn far_4_4834_0_a(.in(layer_3[212]), .out(far_4_4834_0[0]));    relay_conn far_4_4834_0_b(.in(layer_3[100]), .out(far_4_4834_0[1]));
    wire [1:0] far_4_4834_1;    relay_conn far_4_4834_1_a(.in(far_4_4834_0[0]), .out(far_4_4834_1[0]));    relay_conn far_4_4834_1_b(.in(far_4_4834_0[1]), .out(far_4_4834_1[1]));
    wire [1:0] far_4_4834_2;    relay_conn far_4_4834_2_a(.in(far_4_4834_1[0]), .out(far_4_4834_2[0]));    relay_conn far_4_4834_2_b(.in(far_4_4834_1[1]), .out(far_4_4834_2[1]));
    assign layer_4[754] = ~far_4_4834_2[1]; 
    wire [1:0] far_4_4835_0;    relay_conn far_4_4835_0_a(.in(layer_3[834]), .out(far_4_4835_0[0]));    relay_conn far_4_4835_0_b(.in(layer_3[800]), .out(far_4_4835_0[1]));
    assign layer_4[755] = far_4_4835_0[0] | far_4_4835_0[1]; 
    assign layer_4[756] = ~(layer_3[682] & layer_3[678]); 
    wire [1:0] far_4_4837_0;    relay_conn far_4_4837_0_a(.in(layer_3[222]), .out(far_4_4837_0[0]));    relay_conn far_4_4837_0_b(.in(layer_3[169]), .out(far_4_4837_0[1]));
    assign layer_4[757] = far_4_4837_0[1] & ~far_4_4837_0[0]; 
    wire [1:0] far_4_4838_0;    relay_conn far_4_4838_0_a(.in(layer_3[112]), .out(far_4_4838_0[0]));    relay_conn far_4_4838_0_b(.in(layer_3[0]), .out(far_4_4838_0[1]));
    wire [1:0] far_4_4838_1;    relay_conn far_4_4838_1_a(.in(far_4_4838_0[0]), .out(far_4_4838_1[0]));    relay_conn far_4_4838_1_b(.in(far_4_4838_0[1]), .out(far_4_4838_1[1]));
    wire [1:0] far_4_4838_2;    relay_conn far_4_4838_2_a(.in(far_4_4838_1[0]), .out(far_4_4838_2[0]));    relay_conn far_4_4838_2_b(.in(far_4_4838_1[1]), .out(far_4_4838_2[1]));
    assign layer_4[758] = ~far_4_4838_2[0]; 
    assign layer_4[759] = layer_3[134]; 
    assign layer_4[760] = layer_3[542] | layer_3[569]; 
    wire [1:0] far_4_4841_0;    relay_conn far_4_4841_0_a(.in(layer_3[623]), .out(far_4_4841_0[0]));    relay_conn far_4_4841_0_b(.in(layer_3[512]), .out(far_4_4841_0[1]));
    wire [1:0] far_4_4841_1;    relay_conn far_4_4841_1_a(.in(far_4_4841_0[0]), .out(far_4_4841_1[0]));    relay_conn far_4_4841_1_b(.in(far_4_4841_0[1]), .out(far_4_4841_1[1]));
    wire [1:0] far_4_4841_2;    relay_conn far_4_4841_2_a(.in(far_4_4841_1[0]), .out(far_4_4841_2[0]));    relay_conn far_4_4841_2_b(.in(far_4_4841_1[1]), .out(far_4_4841_2[1]));
    assign layer_4[761] = far_4_4841_2[1] & ~far_4_4841_2[0]; 
    wire [1:0] far_4_4842_0;    relay_conn far_4_4842_0_a(.in(layer_3[12]), .out(far_4_4842_0[0]));    relay_conn far_4_4842_0_b(.in(layer_3[113]), .out(far_4_4842_0[1]));
    wire [1:0] far_4_4842_1;    relay_conn far_4_4842_1_a(.in(far_4_4842_0[0]), .out(far_4_4842_1[0]));    relay_conn far_4_4842_1_b(.in(far_4_4842_0[1]), .out(far_4_4842_1[1]));
    wire [1:0] far_4_4842_2;    relay_conn far_4_4842_2_a(.in(far_4_4842_1[0]), .out(far_4_4842_2[0]));    relay_conn far_4_4842_2_b(.in(far_4_4842_1[1]), .out(far_4_4842_2[1]));
    assign layer_4[762] = ~far_4_4842_2[1] | (far_4_4842_2[0] & far_4_4842_2[1]); 
    assign layer_4[763] = layer_3[198]; 
    assign layer_4[764] = ~layer_3[963] | (layer_3[963] & layer_3[988]); 
    wire [1:0] far_4_4845_0;    relay_conn far_4_4845_0_a(.in(layer_3[942]), .out(far_4_4845_0[0]));    relay_conn far_4_4845_0_b(.in(layer_3[994]), .out(far_4_4845_0[1]));
    assign layer_4[765] = far_4_4845_0[0] & ~far_4_4845_0[1]; 
    wire [1:0] far_4_4846_0;    relay_conn far_4_4846_0_a(.in(layer_3[408]), .out(far_4_4846_0[0]));    relay_conn far_4_4846_0_b(.in(layer_3[467]), .out(far_4_4846_0[1]));
    assign layer_4[766] = ~far_4_4846_0[0]; 
    wire [1:0] far_4_4847_0;    relay_conn far_4_4847_0_a(.in(layer_3[726]), .out(far_4_4847_0[0]));    relay_conn far_4_4847_0_b(.in(layer_3[823]), .out(far_4_4847_0[1]));
    wire [1:0] far_4_4847_1;    relay_conn far_4_4847_1_a(.in(far_4_4847_0[0]), .out(far_4_4847_1[0]));    relay_conn far_4_4847_1_b(.in(far_4_4847_0[1]), .out(far_4_4847_1[1]));
    wire [1:0] far_4_4847_2;    relay_conn far_4_4847_2_a(.in(far_4_4847_1[0]), .out(far_4_4847_2[0]));    relay_conn far_4_4847_2_b(.in(far_4_4847_1[1]), .out(far_4_4847_2[1]));
    assign layer_4[767] = ~(far_4_4847_2[0] & far_4_4847_2[1]); 
    assign layer_4[768] = ~layer_3[341] | (layer_3[341] & layer_3[323]); 
    wire [1:0] far_4_4849_0;    relay_conn far_4_4849_0_a(.in(layer_3[900]), .out(far_4_4849_0[0]));    relay_conn far_4_4849_0_b(.in(layer_3[953]), .out(far_4_4849_0[1]));
    assign layer_4[769] = ~(far_4_4849_0[0] & far_4_4849_0[1]); 
    wire [1:0] far_4_4850_0;    relay_conn far_4_4850_0_a(.in(layer_3[164]), .out(far_4_4850_0[0]));    relay_conn far_4_4850_0_b(.in(layer_3[56]), .out(far_4_4850_0[1]));
    wire [1:0] far_4_4850_1;    relay_conn far_4_4850_1_a(.in(far_4_4850_0[0]), .out(far_4_4850_1[0]));    relay_conn far_4_4850_1_b(.in(far_4_4850_0[1]), .out(far_4_4850_1[1]));
    wire [1:0] far_4_4850_2;    relay_conn far_4_4850_2_a(.in(far_4_4850_1[0]), .out(far_4_4850_2[0]));    relay_conn far_4_4850_2_b(.in(far_4_4850_1[1]), .out(far_4_4850_2[1]));
    assign layer_4[770] = far_4_4850_2[0] | far_4_4850_2[1]; 
    assign layer_4[771] = ~layer_3[981]; 
    wire [1:0] far_4_4852_0;    relay_conn far_4_4852_0_a(.in(layer_3[887]), .out(far_4_4852_0[0]));    relay_conn far_4_4852_0_b(.in(layer_3[990]), .out(far_4_4852_0[1]));
    wire [1:0] far_4_4852_1;    relay_conn far_4_4852_1_a(.in(far_4_4852_0[0]), .out(far_4_4852_1[0]));    relay_conn far_4_4852_1_b(.in(far_4_4852_0[1]), .out(far_4_4852_1[1]));
    wire [1:0] far_4_4852_2;    relay_conn far_4_4852_2_a(.in(far_4_4852_1[0]), .out(far_4_4852_2[0]));    relay_conn far_4_4852_2_b(.in(far_4_4852_1[1]), .out(far_4_4852_2[1]));
    assign layer_4[772] = ~(far_4_4852_2[0] | far_4_4852_2[1]); 
    assign layer_4[773] = layer_3[807]; 
    wire [1:0] far_4_4854_0;    relay_conn far_4_4854_0_a(.in(layer_3[115]), .out(far_4_4854_0[0]));    relay_conn far_4_4854_0_b(.in(layer_3[222]), .out(far_4_4854_0[1]));
    wire [1:0] far_4_4854_1;    relay_conn far_4_4854_1_a(.in(far_4_4854_0[0]), .out(far_4_4854_1[0]));    relay_conn far_4_4854_1_b(.in(far_4_4854_0[1]), .out(far_4_4854_1[1]));
    wire [1:0] far_4_4854_2;    relay_conn far_4_4854_2_a(.in(far_4_4854_1[0]), .out(far_4_4854_2[0]));    relay_conn far_4_4854_2_b(.in(far_4_4854_1[1]), .out(far_4_4854_2[1]));
    assign layer_4[774] = ~far_4_4854_2[1]; 
    wire [1:0] far_4_4855_0;    relay_conn far_4_4855_0_a(.in(layer_3[756]), .out(far_4_4855_0[0]));    relay_conn far_4_4855_0_b(.in(layer_3[838]), .out(far_4_4855_0[1]));
    wire [1:0] far_4_4855_1;    relay_conn far_4_4855_1_a(.in(far_4_4855_0[0]), .out(far_4_4855_1[0]));    relay_conn far_4_4855_1_b(.in(far_4_4855_0[1]), .out(far_4_4855_1[1]));
    assign layer_4[775] = far_4_4855_1[1] & ~far_4_4855_1[0]; 
    wire [1:0] far_4_4856_0;    relay_conn far_4_4856_0_a(.in(layer_3[829]), .out(far_4_4856_0[0]));    relay_conn far_4_4856_0_b(.in(layer_3[702]), .out(far_4_4856_0[1]));
    wire [1:0] far_4_4856_1;    relay_conn far_4_4856_1_a(.in(far_4_4856_0[0]), .out(far_4_4856_1[0]));    relay_conn far_4_4856_1_b(.in(far_4_4856_0[1]), .out(far_4_4856_1[1]));
    wire [1:0] far_4_4856_2;    relay_conn far_4_4856_2_a(.in(far_4_4856_1[0]), .out(far_4_4856_2[0]));    relay_conn far_4_4856_2_b(.in(far_4_4856_1[1]), .out(far_4_4856_2[1]));
    assign layer_4[776] = ~far_4_4856_2[1] | (far_4_4856_2[0] & far_4_4856_2[1]); 
    wire [1:0] far_4_4857_0;    relay_conn far_4_4857_0_a(.in(layer_3[287]), .out(far_4_4857_0[0]));    relay_conn far_4_4857_0_b(.in(layer_3[402]), .out(far_4_4857_0[1]));
    wire [1:0] far_4_4857_1;    relay_conn far_4_4857_1_a(.in(far_4_4857_0[0]), .out(far_4_4857_1[0]));    relay_conn far_4_4857_1_b(.in(far_4_4857_0[1]), .out(far_4_4857_1[1]));
    wire [1:0] far_4_4857_2;    relay_conn far_4_4857_2_a(.in(far_4_4857_1[0]), .out(far_4_4857_2[0]));    relay_conn far_4_4857_2_b(.in(far_4_4857_1[1]), .out(far_4_4857_2[1]));
    assign layer_4[777] = ~far_4_4857_2[1]; 
    wire [1:0] far_4_4858_0;    relay_conn far_4_4858_0_a(.in(layer_3[572]), .out(far_4_4858_0[0]));    relay_conn far_4_4858_0_b(.in(layer_3[674]), .out(far_4_4858_0[1]));
    wire [1:0] far_4_4858_1;    relay_conn far_4_4858_1_a(.in(far_4_4858_0[0]), .out(far_4_4858_1[0]));    relay_conn far_4_4858_1_b(.in(far_4_4858_0[1]), .out(far_4_4858_1[1]));
    wire [1:0] far_4_4858_2;    relay_conn far_4_4858_2_a(.in(far_4_4858_1[0]), .out(far_4_4858_2[0]));    relay_conn far_4_4858_2_b(.in(far_4_4858_1[1]), .out(far_4_4858_2[1]));
    assign layer_4[778] = far_4_4858_2[0] & ~far_4_4858_2[1]; 
    wire [1:0] far_4_4859_0;    relay_conn far_4_4859_0_a(.in(layer_3[780]), .out(far_4_4859_0[0]));    relay_conn far_4_4859_0_b(.in(layer_3[871]), .out(far_4_4859_0[1]));
    wire [1:0] far_4_4859_1;    relay_conn far_4_4859_1_a(.in(far_4_4859_0[0]), .out(far_4_4859_1[0]));    relay_conn far_4_4859_1_b(.in(far_4_4859_0[1]), .out(far_4_4859_1[1]));
    assign layer_4[779] = far_4_4859_1[0] ^ far_4_4859_1[1]; 
    assign layer_4[780] = ~layer_3[979]; 
    wire [1:0] far_4_4861_0;    relay_conn far_4_4861_0_a(.in(layer_3[935]), .out(far_4_4861_0[0]));    relay_conn far_4_4861_0_b(.in(layer_3[986]), .out(far_4_4861_0[1]));
    assign layer_4[781] = ~far_4_4861_0[1] | (far_4_4861_0[0] & far_4_4861_0[1]); 
    assign layer_4[782] = ~(layer_3[329] | layer_3[337]); 
    wire [1:0] far_4_4863_0;    relay_conn far_4_4863_0_a(.in(layer_3[0]), .out(far_4_4863_0[0]));    relay_conn far_4_4863_0_b(.in(layer_3[62]), .out(far_4_4863_0[1]));
    assign layer_4[783] = ~(far_4_4863_0[0] & far_4_4863_0[1]); 
    wire [1:0] far_4_4864_0;    relay_conn far_4_4864_0_a(.in(layer_3[332]), .out(far_4_4864_0[0]));    relay_conn far_4_4864_0_b(.in(layer_3[239]), .out(far_4_4864_0[1]));
    wire [1:0] far_4_4864_1;    relay_conn far_4_4864_1_a(.in(far_4_4864_0[0]), .out(far_4_4864_1[0]));    relay_conn far_4_4864_1_b(.in(far_4_4864_0[1]), .out(far_4_4864_1[1]));
    assign layer_4[784] = ~far_4_4864_1[0] | (far_4_4864_1[0] & far_4_4864_1[1]); 
    assign layer_4[785] = ~layer_3[604]; 
    wire [1:0] far_4_4866_0;    relay_conn far_4_4866_0_a(.in(layer_3[948]), .out(far_4_4866_0[0]));    relay_conn far_4_4866_0_b(.in(layer_3[1008]), .out(far_4_4866_0[1]));
    assign layer_4[786] = far_4_4866_0[0]; 
    wire [1:0] far_4_4867_0;    relay_conn far_4_4867_0_a(.in(layer_3[692]), .out(far_4_4867_0[0]));    relay_conn far_4_4867_0_b(.in(layer_3[815]), .out(far_4_4867_0[1]));
    wire [1:0] far_4_4867_1;    relay_conn far_4_4867_1_a(.in(far_4_4867_0[0]), .out(far_4_4867_1[0]));    relay_conn far_4_4867_1_b(.in(far_4_4867_0[1]), .out(far_4_4867_1[1]));
    wire [1:0] far_4_4867_2;    relay_conn far_4_4867_2_a(.in(far_4_4867_1[0]), .out(far_4_4867_2[0]));    relay_conn far_4_4867_2_b(.in(far_4_4867_1[1]), .out(far_4_4867_2[1]));
    assign layer_4[787] = far_4_4867_2[0] & ~far_4_4867_2[1]; 
    wire [1:0] far_4_4868_0;    relay_conn far_4_4868_0_a(.in(layer_3[334]), .out(far_4_4868_0[0]));    relay_conn far_4_4868_0_b(.in(layer_3[375]), .out(far_4_4868_0[1]));
    assign layer_4[788] = ~far_4_4868_0[1] | (far_4_4868_0[0] & far_4_4868_0[1]); 
    wire [1:0] far_4_4869_0;    relay_conn far_4_4869_0_a(.in(layer_3[837]), .out(far_4_4869_0[0]));    relay_conn far_4_4869_0_b(.in(layer_3[942]), .out(far_4_4869_0[1]));
    wire [1:0] far_4_4869_1;    relay_conn far_4_4869_1_a(.in(far_4_4869_0[0]), .out(far_4_4869_1[0]));    relay_conn far_4_4869_1_b(.in(far_4_4869_0[1]), .out(far_4_4869_1[1]));
    wire [1:0] far_4_4869_2;    relay_conn far_4_4869_2_a(.in(far_4_4869_1[0]), .out(far_4_4869_2[0]));    relay_conn far_4_4869_2_b(.in(far_4_4869_1[1]), .out(far_4_4869_2[1]));
    assign layer_4[789] = ~(far_4_4869_2[0] & far_4_4869_2[1]); 
    assign layer_4[790] = layer_3[516]; 
    wire [1:0] far_4_4871_0;    relay_conn far_4_4871_0_a(.in(layer_3[223]), .out(far_4_4871_0[0]));    relay_conn far_4_4871_0_b(.in(layer_3[302]), .out(far_4_4871_0[1]));
    wire [1:0] far_4_4871_1;    relay_conn far_4_4871_1_a(.in(far_4_4871_0[0]), .out(far_4_4871_1[0]));    relay_conn far_4_4871_1_b(.in(far_4_4871_0[1]), .out(far_4_4871_1[1]));
    assign layer_4[791] = ~(far_4_4871_1[0] & far_4_4871_1[1]); 
    assign layer_4[792] = ~layer_3[674]; 
    assign layer_4[793] = ~(layer_3[909] & layer_3[901]); 
    wire [1:0] far_4_4874_0;    relay_conn far_4_4874_0_a(.in(layer_3[769]), .out(far_4_4874_0[0]));    relay_conn far_4_4874_0_b(.in(layer_3[700]), .out(far_4_4874_0[1]));
    wire [1:0] far_4_4874_1;    relay_conn far_4_4874_1_a(.in(far_4_4874_0[0]), .out(far_4_4874_1[0]));    relay_conn far_4_4874_1_b(.in(far_4_4874_0[1]), .out(far_4_4874_1[1]));
    assign layer_4[794] = far_4_4874_1[1]; 
    assign layer_4[795] = ~layer_3[18] | (layer_3[18] & layer_3[10]); 
    assign layer_4[796] = layer_3[593]; 
    wire [1:0] far_4_4877_0;    relay_conn far_4_4877_0_a(.in(layer_3[475]), .out(far_4_4877_0[0]));    relay_conn far_4_4877_0_b(.in(layer_3[547]), .out(far_4_4877_0[1]));
    wire [1:0] far_4_4877_1;    relay_conn far_4_4877_1_a(.in(far_4_4877_0[0]), .out(far_4_4877_1[0]));    relay_conn far_4_4877_1_b(.in(far_4_4877_0[1]), .out(far_4_4877_1[1]));
    assign layer_4[797] = far_4_4877_1[1]; 
    assign layer_4[798] = layer_3[319] & layer_3[335]; 
    wire [1:0] far_4_4879_0;    relay_conn far_4_4879_0_a(.in(layer_3[68]), .out(far_4_4879_0[0]));    relay_conn far_4_4879_0_b(.in(layer_3[149]), .out(far_4_4879_0[1]));
    wire [1:0] far_4_4879_1;    relay_conn far_4_4879_1_a(.in(far_4_4879_0[0]), .out(far_4_4879_1[0]));    relay_conn far_4_4879_1_b(.in(far_4_4879_0[1]), .out(far_4_4879_1[1]));
    assign layer_4[799] = far_4_4879_1[0] & far_4_4879_1[1]; 
    assign layer_4[800] = layer_3[391] & ~layer_3[382]; 
    wire [1:0] far_4_4881_0;    relay_conn far_4_4881_0_a(.in(layer_3[112]), .out(far_4_4881_0[0]));    relay_conn far_4_4881_0_b(.in(layer_3[165]), .out(far_4_4881_0[1]));
    assign layer_4[801] = ~far_4_4881_0[1] | (far_4_4881_0[0] & far_4_4881_0[1]); 
    wire [1:0] far_4_4882_0;    relay_conn far_4_4882_0_a(.in(layer_3[900]), .out(far_4_4882_0[0]));    relay_conn far_4_4882_0_b(.in(layer_3[950]), .out(far_4_4882_0[1]));
    assign layer_4[802] = far_4_4882_0[1]; 
    wire [1:0] far_4_4883_0;    relay_conn far_4_4883_0_a(.in(layer_3[676]), .out(far_4_4883_0[0]));    relay_conn far_4_4883_0_b(.in(layer_3[584]), .out(far_4_4883_0[1]));
    wire [1:0] far_4_4883_1;    relay_conn far_4_4883_1_a(.in(far_4_4883_0[0]), .out(far_4_4883_1[0]));    relay_conn far_4_4883_1_b(.in(far_4_4883_0[1]), .out(far_4_4883_1[1]));
    assign layer_4[803] = far_4_4883_1[1] & ~far_4_4883_1[0]; 
    wire [1:0] far_4_4884_0;    relay_conn far_4_4884_0_a(.in(layer_3[420]), .out(far_4_4884_0[0]));    relay_conn far_4_4884_0_b(.in(layer_3[459]), .out(far_4_4884_0[1]));
    assign layer_4[804] = ~(far_4_4884_0[0] & far_4_4884_0[1]); 
    wire [1:0] far_4_4885_0;    relay_conn far_4_4885_0_a(.in(layer_3[376]), .out(far_4_4885_0[0]));    relay_conn far_4_4885_0_b(.in(layer_3[410]), .out(far_4_4885_0[1]));
    assign layer_4[805] = ~far_4_4885_0[1]; 
    wire [1:0] far_4_4886_0;    relay_conn far_4_4886_0_a(.in(layer_3[882]), .out(far_4_4886_0[0]));    relay_conn far_4_4886_0_b(.in(layer_3[956]), .out(far_4_4886_0[1]));
    wire [1:0] far_4_4886_1;    relay_conn far_4_4886_1_a(.in(far_4_4886_0[0]), .out(far_4_4886_1[0]));    relay_conn far_4_4886_1_b(.in(far_4_4886_0[1]), .out(far_4_4886_1[1]));
    assign layer_4[806] = far_4_4886_1[1] & ~far_4_4886_1[0]; 
    assign layer_4[807] = layer_3[58] ^ layer_3[81]; 
    wire [1:0] far_4_4888_0;    relay_conn far_4_4888_0_a(.in(layer_3[433]), .out(far_4_4888_0[0]));    relay_conn far_4_4888_0_b(.in(layer_3[314]), .out(far_4_4888_0[1]));
    wire [1:0] far_4_4888_1;    relay_conn far_4_4888_1_a(.in(far_4_4888_0[0]), .out(far_4_4888_1[0]));    relay_conn far_4_4888_1_b(.in(far_4_4888_0[1]), .out(far_4_4888_1[1]));
    wire [1:0] far_4_4888_2;    relay_conn far_4_4888_2_a(.in(far_4_4888_1[0]), .out(far_4_4888_2[0]));    relay_conn far_4_4888_2_b(.in(far_4_4888_1[1]), .out(far_4_4888_2[1]));
    assign layer_4[808] = ~far_4_4888_2[1]; 
    wire [1:0] far_4_4889_0;    relay_conn far_4_4889_0_a(.in(layer_3[775]), .out(far_4_4889_0[0]));    relay_conn far_4_4889_0_b(.in(layer_3[715]), .out(far_4_4889_0[1]));
    assign layer_4[809] = ~far_4_4889_0[1]; 
    wire [1:0] far_4_4890_0;    relay_conn far_4_4890_0_a(.in(layer_3[383]), .out(far_4_4890_0[0]));    relay_conn far_4_4890_0_b(.in(layer_3[454]), .out(far_4_4890_0[1]));
    wire [1:0] far_4_4890_1;    relay_conn far_4_4890_1_a(.in(far_4_4890_0[0]), .out(far_4_4890_1[0]));    relay_conn far_4_4890_1_b(.in(far_4_4890_0[1]), .out(far_4_4890_1[1]));
    assign layer_4[810] = ~far_4_4890_1[0] | (far_4_4890_1[0] & far_4_4890_1[1]); 
    assign layer_4[811] = layer_3[492]; 
    wire [1:0] far_4_4892_0;    relay_conn far_4_4892_0_a(.in(layer_3[834]), .out(far_4_4892_0[0]));    relay_conn far_4_4892_0_b(.in(layer_3[937]), .out(far_4_4892_0[1]));
    wire [1:0] far_4_4892_1;    relay_conn far_4_4892_1_a(.in(far_4_4892_0[0]), .out(far_4_4892_1[0]));    relay_conn far_4_4892_1_b(.in(far_4_4892_0[1]), .out(far_4_4892_1[1]));
    wire [1:0] far_4_4892_2;    relay_conn far_4_4892_2_a(.in(far_4_4892_1[0]), .out(far_4_4892_2[0]));    relay_conn far_4_4892_2_b(.in(far_4_4892_1[1]), .out(far_4_4892_2[1]));
    assign layer_4[812] = far_4_4892_2[0]; 
    wire [1:0] far_4_4893_0;    relay_conn far_4_4893_0_a(.in(layer_3[930]), .out(far_4_4893_0[0]));    relay_conn far_4_4893_0_b(.in(layer_3[885]), .out(far_4_4893_0[1]));
    assign layer_4[813] = far_4_4893_0[0] & ~far_4_4893_0[1]; 
    assign layer_4[814] = layer_3[153]; 
    wire [1:0] far_4_4895_0;    relay_conn far_4_4895_0_a(.in(layer_3[233]), .out(far_4_4895_0[0]));    relay_conn far_4_4895_0_b(.in(layer_3[115]), .out(far_4_4895_0[1]));
    wire [1:0] far_4_4895_1;    relay_conn far_4_4895_1_a(.in(far_4_4895_0[0]), .out(far_4_4895_1[0]));    relay_conn far_4_4895_1_b(.in(far_4_4895_0[1]), .out(far_4_4895_1[1]));
    wire [1:0] far_4_4895_2;    relay_conn far_4_4895_2_a(.in(far_4_4895_1[0]), .out(far_4_4895_2[0]));    relay_conn far_4_4895_2_b(.in(far_4_4895_1[1]), .out(far_4_4895_2[1]));
    assign layer_4[815] = ~far_4_4895_2[1]; 
    wire [1:0] far_4_4896_0;    relay_conn far_4_4896_0_a(.in(layer_3[456]), .out(far_4_4896_0[0]));    relay_conn far_4_4896_0_b(.in(layer_3[540]), .out(far_4_4896_0[1]));
    wire [1:0] far_4_4896_1;    relay_conn far_4_4896_1_a(.in(far_4_4896_0[0]), .out(far_4_4896_1[0]));    relay_conn far_4_4896_1_b(.in(far_4_4896_0[1]), .out(far_4_4896_1[1]));
    assign layer_4[816] = ~(far_4_4896_1[0] | far_4_4896_1[1]); 
    wire [1:0] far_4_4897_0;    relay_conn far_4_4897_0_a(.in(layer_3[347]), .out(far_4_4897_0[0]));    relay_conn far_4_4897_0_b(.in(layer_3[312]), .out(far_4_4897_0[1]));
    assign layer_4[817] = ~far_4_4897_0[1]; 
    wire [1:0] far_4_4898_0;    relay_conn far_4_4898_0_a(.in(layer_3[681]), .out(far_4_4898_0[0]));    relay_conn far_4_4898_0_b(.in(layer_3[755]), .out(far_4_4898_0[1]));
    wire [1:0] far_4_4898_1;    relay_conn far_4_4898_1_a(.in(far_4_4898_0[0]), .out(far_4_4898_1[0]));    relay_conn far_4_4898_1_b(.in(far_4_4898_0[1]), .out(far_4_4898_1[1]));
    assign layer_4[818] = far_4_4898_1[0] & far_4_4898_1[1]; 
    wire [1:0] far_4_4899_0;    relay_conn far_4_4899_0_a(.in(layer_3[100]), .out(far_4_4899_0[0]));    relay_conn far_4_4899_0_b(.in(layer_3[64]), .out(far_4_4899_0[1]));
    assign layer_4[819] = ~far_4_4899_0[0] | (far_4_4899_0[0] & far_4_4899_0[1]); 
    wire [1:0] far_4_4900_0;    relay_conn far_4_4900_0_a(.in(layer_3[753]), .out(far_4_4900_0[0]));    relay_conn far_4_4900_0_b(.in(layer_3[695]), .out(far_4_4900_0[1]));
    assign layer_4[820] = far_4_4900_0[0]; 
    assign layer_4[821] = layer_3[952] & layer_3[924]; 
    wire [1:0] far_4_4902_0;    relay_conn far_4_4902_0_a(.in(layer_3[979]), .out(far_4_4902_0[0]));    relay_conn far_4_4902_0_b(.in(layer_3[909]), .out(far_4_4902_0[1]));
    wire [1:0] far_4_4902_1;    relay_conn far_4_4902_1_a(.in(far_4_4902_0[0]), .out(far_4_4902_1[0]));    relay_conn far_4_4902_1_b(.in(far_4_4902_0[1]), .out(far_4_4902_1[1]));
    assign layer_4[822] = ~far_4_4902_1[0] | (far_4_4902_1[0] & far_4_4902_1[1]); 
    wire [1:0] far_4_4903_0;    relay_conn far_4_4903_0_a(.in(layer_3[113]), .out(far_4_4903_0[0]));    relay_conn far_4_4903_0_b(.in(layer_3[47]), .out(far_4_4903_0[1]));
    wire [1:0] far_4_4903_1;    relay_conn far_4_4903_1_a(.in(far_4_4903_0[0]), .out(far_4_4903_1[0]));    relay_conn far_4_4903_1_b(.in(far_4_4903_0[1]), .out(far_4_4903_1[1]));
    assign layer_4[823] = far_4_4903_1[0] | far_4_4903_1[1]; 
    wire [1:0] far_4_4904_0;    relay_conn far_4_4904_0_a(.in(layer_3[367]), .out(far_4_4904_0[0]));    relay_conn far_4_4904_0_b(.in(layer_3[299]), .out(far_4_4904_0[1]));
    wire [1:0] far_4_4904_1;    relay_conn far_4_4904_1_a(.in(far_4_4904_0[0]), .out(far_4_4904_1[0]));    relay_conn far_4_4904_1_b(.in(far_4_4904_0[1]), .out(far_4_4904_1[1]));
    assign layer_4[824] = ~far_4_4904_1[0]; 
    wire [1:0] far_4_4905_0;    relay_conn far_4_4905_0_a(.in(layer_3[1000]), .out(far_4_4905_0[0]));    relay_conn far_4_4905_0_b(.in(layer_3[909]), .out(far_4_4905_0[1]));
    wire [1:0] far_4_4905_1;    relay_conn far_4_4905_1_a(.in(far_4_4905_0[0]), .out(far_4_4905_1[0]));    relay_conn far_4_4905_1_b(.in(far_4_4905_0[1]), .out(far_4_4905_1[1]));
    assign layer_4[825] = far_4_4905_1[1] & ~far_4_4905_1[0]; 
    wire [1:0] far_4_4906_0;    relay_conn far_4_4906_0_a(.in(layer_3[744]), .out(far_4_4906_0[0]));    relay_conn far_4_4906_0_b(.in(layer_3[835]), .out(far_4_4906_0[1]));
    wire [1:0] far_4_4906_1;    relay_conn far_4_4906_1_a(.in(far_4_4906_0[0]), .out(far_4_4906_1[0]));    relay_conn far_4_4906_1_b(.in(far_4_4906_0[1]), .out(far_4_4906_1[1]));
    assign layer_4[826] = far_4_4906_1[0] & far_4_4906_1[1]; 
    wire [1:0] far_4_4907_0;    relay_conn far_4_4907_0_a(.in(layer_3[102]), .out(far_4_4907_0[0]));    relay_conn far_4_4907_0_b(.in(layer_3[222]), .out(far_4_4907_0[1]));
    wire [1:0] far_4_4907_1;    relay_conn far_4_4907_1_a(.in(far_4_4907_0[0]), .out(far_4_4907_1[0]));    relay_conn far_4_4907_1_b(.in(far_4_4907_0[1]), .out(far_4_4907_1[1]));
    wire [1:0] far_4_4907_2;    relay_conn far_4_4907_2_a(.in(far_4_4907_1[0]), .out(far_4_4907_2[0]));    relay_conn far_4_4907_2_b(.in(far_4_4907_1[1]), .out(far_4_4907_2[1]));
    assign layer_4[827] = far_4_4907_2[0] & ~far_4_4907_2[1]; 
    assign layer_4[828] = ~layer_3[443]; 
    assign layer_4[829] = ~layer_3[695]; 
    wire [1:0] far_4_4910_0;    relay_conn far_4_4910_0_a(.in(layer_3[318]), .out(far_4_4910_0[0]));    relay_conn far_4_4910_0_b(.in(layer_3[266]), .out(far_4_4910_0[1]));
    assign layer_4[830] = far_4_4910_0[1]; 
    wire [1:0] far_4_4911_0;    relay_conn far_4_4911_0_a(.in(layer_3[871]), .out(far_4_4911_0[0]));    relay_conn far_4_4911_0_b(.in(layer_3[807]), .out(far_4_4911_0[1]));
    wire [1:0] far_4_4911_1;    relay_conn far_4_4911_1_a(.in(far_4_4911_0[0]), .out(far_4_4911_1[0]));    relay_conn far_4_4911_1_b(.in(far_4_4911_0[1]), .out(far_4_4911_1[1]));
    assign layer_4[831] = far_4_4911_1[0] | far_4_4911_1[1]; 
    assign layer_4[832] = layer_3[395] | layer_3[400]; 
    wire [1:0] far_4_4913_0;    relay_conn far_4_4913_0_a(.in(layer_3[931]), .out(far_4_4913_0[0]));    relay_conn far_4_4913_0_b(.in(layer_3[884]), .out(far_4_4913_0[1]));
    assign layer_4[833] = ~(far_4_4913_0[0] & far_4_4913_0[1]); 
    assign layer_4[834] = ~layer_3[32] | (layer_3[32] & layer_3[56]); 
    wire [1:0] far_4_4915_0;    relay_conn far_4_4915_0_a(.in(layer_3[72]), .out(far_4_4915_0[0]));    relay_conn far_4_4915_0_b(.in(layer_3[122]), .out(far_4_4915_0[1]));
    assign layer_4[835] = far_4_4915_0[1]; 
    wire [1:0] far_4_4916_0;    relay_conn far_4_4916_0_a(.in(layer_3[261]), .out(far_4_4916_0[0]));    relay_conn far_4_4916_0_b(.in(layer_3[323]), .out(far_4_4916_0[1]));
    assign layer_4[836] = ~far_4_4916_0[0] | (far_4_4916_0[0] & far_4_4916_0[1]); 
    wire [1:0] far_4_4917_0;    relay_conn far_4_4917_0_a(.in(layer_3[908]), .out(far_4_4917_0[0]));    relay_conn far_4_4917_0_b(.in(layer_3[834]), .out(far_4_4917_0[1]));
    wire [1:0] far_4_4917_1;    relay_conn far_4_4917_1_a(.in(far_4_4917_0[0]), .out(far_4_4917_1[0]));    relay_conn far_4_4917_1_b(.in(far_4_4917_0[1]), .out(far_4_4917_1[1]));
    assign layer_4[837] = far_4_4917_1[1]; 
    wire [1:0] far_4_4918_0;    relay_conn far_4_4918_0_a(.in(layer_3[352]), .out(far_4_4918_0[0]));    relay_conn far_4_4918_0_b(.in(layer_3[390]), .out(far_4_4918_0[1]));
    assign layer_4[838] = ~far_4_4918_0[0]; 
    wire [1:0] far_4_4919_0;    relay_conn far_4_4919_0_a(.in(layer_3[1018]), .out(far_4_4919_0[0]));    relay_conn far_4_4919_0_b(.in(layer_3[915]), .out(far_4_4919_0[1]));
    wire [1:0] far_4_4919_1;    relay_conn far_4_4919_1_a(.in(far_4_4919_0[0]), .out(far_4_4919_1[0]));    relay_conn far_4_4919_1_b(.in(far_4_4919_0[1]), .out(far_4_4919_1[1]));
    wire [1:0] far_4_4919_2;    relay_conn far_4_4919_2_a(.in(far_4_4919_1[0]), .out(far_4_4919_2[0]));    relay_conn far_4_4919_2_b(.in(far_4_4919_1[1]), .out(far_4_4919_2[1]));
    assign layer_4[839] = far_4_4919_2[1] & ~far_4_4919_2[0]; 
    assign layer_4[840] = layer_3[56] & ~layer_3[35]; 
    assign layer_4[841] = ~(layer_3[420] ^ layer_3[398]); 
    wire [1:0] far_4_4922_0;    relay_conn far_4_4922_0_a(.in(layer_3[700]), .out(far_4_4922_0[0]));    relay_conn far_4_4922_0_b(.in(layer_3[782]), .out(far_4_4922_0[1]));
    wire [1:0] far_4_4922_1;    relay_conn far_4_4922_1_a(.in(far_4_4922_0[0]), .out(far_4_4922_1[0]));    relay_conn far_4_4922_1_b(.in(far_4_4922_0[1]), .out(far_4_4922_1[1]));
    assign layer_4[842] = far_4_4922_1[1] & ~far_4_4922_1[0]; 
    wire [1:0] far_4_4923_0;    relay_conn far_4_4923_0_a(.in(layer_3[648]), .out(far_4_4923_0[0]));    relay_conn far_4_4923_0_b(.in(layer_3[572]), .out(far_4_4923_0[1]));
    wire [1:0] far_4_4923_1;    relay_conn far_4_4923_1_a(.in(far_4_4923_0[0]), .out(far_4_4923_1[0]));    relay_conn far_4_4923_1_b(.in(far_4_4923_0[1]), .out(far_4_4923_1[1]));
    assign layer_4[843] = ~(far_4_4923_1[0] ^ far_4_4923_1[1]); 
    wire [1:0] far_4_4924_0;    relay_conn far_4_4924_0_a(.in(layer_3[419]), .out(far_4_4924_0[0]));    relay_conn far_4_4924_0_b(.in(layer_3[347]), .out(far_4_4924_0[1]));
    wire [1:0] far_4_4924_1;    relay_conn far_4_4924_1_a(.in(far_4_4924_0[0]), .out(far_4_4924_1[0]));    relay_conn far_4_4924_1_b(.in(far_4_4924_0[1]), .out(far_4_4924_1[1]));
    assign layer_4[844] = ~far_4_4924_1[0] | (far_4_4924_1[0] & far_4_4924_1[1]); 
    wire [1:0] far_4_4925_0;    relay_conn far_4_4925_0_a(.in(layer_3[843]), .out(far_4_4925_0[0]));    relay_conn far_4_4925_0_b(.in(layer_3[969]), .out(far_4_4925_0[1]));
    wire [1:0] far_4_4925_1;    relay_conn far_4_4925_1_a(.in(far_4_4925_0[0]), .out(far_4_4925_1[0]));    relay_conn far_4_4925_1_b(.in(far_4_4925_0[1]), .out(far_4_4925_1[1]));
    wire [1:0] far_4_4925_2;    relay_conn far_4_4925_2_a(.in(far_4_4925_1[0]), .out(far_4_4925_2[0]));    relay_conn far_4_4925_2_b(.in(far_4_4925_1[1]), .out(far_4_4925_2[1]));
    assign layer_4[845] = ~far_4_4925_2[0]; 
    wire [1:0] far_4_4926_0;    relay_conn far_4_4926_0_a(.in(layer_3[1003]), .out(far_4_4926_0[0]));    relay_conn far_4_4926_0_b(.in(layer_3[916]), .out(far_4_4926_0[1]));
    wire [1:0] far_4_4926_1;    relay_conn far_4_4926_1_a(.in(far_4_4926_0[0]), .out(far_4_4926_1[0]));    relay_conn far_4_4926_1_b(.in(far_4_4926_0[1]), .out(far_4_4926_1[1]));
    assign layer_4[846] = far_4_4926_1[1]; 
    wire [1:0] far_4_4927_0;    relay_conn far_4_4927_0_a(.in(layer_3[253]), .out(far_4_4927_0[0]));    relay_conn far_4_4927_0_b(.in(layer_3[352]), .out(far_4_4927_0[1]));
    wire [1:0] far_4_4927_1;    relay_conn far_4_4927_1_a(.in(far_4_4927_0[0]), .out(far_4_4927_1[0]));    relay_conn far_4_4927_1_b(.in(far_4_4927_0[1]), .out(far_4_4927_1[1]));
    wire [1:0] far_4_4927_2;    relay_conn far_4_4927_2_a(.in(far_4_4927_1[0]), .out(far_4_4927_2[0]));    relay_conn far_4_4927_2_b(.in(far_4_4927_1[1]), .out(far_4_4927_2[1]));
    assign layer_4[847] = ~far_4_4927_2[0] | (far_4_4927_2[0] & far_4_4927_2[1]); 
    wire [1:0] far_4_4928_0;    relay_conn far_4_4928_0_a(.in(layer_3[778]), .out(far_4_4928_0[0]));    relay_conn far_4_4928_0_b(.in(layer_3[823]), .out(far_4_4928_0[1]));
    assign layer_4[848] = far_4_4928_0[0]; 
    wire [1:0] far_4_4929_0;    relay_conn far_4_4929_0_a(.in(layer_3[321]), .out(far_4_4929_0[0]));    relay_conn far_4_4929_0_b(.in(layer_3[289]), .out(far_4_4929_0[1]));
    assign layer_4[849] = far_4_4929_0[0] | far_4_4929_0[1]; 
    wire [1:0] far_4_4930_0;    relay_conn far_4_4930_0_a(.in(layer_3[428]), .out(far_4_4930_0[0]));    relay_conn far_4_4930_0_b(.in(layer_3[359]), .out(far_4_4930_0[1]));
    wire [1:0] far_4_4930_1;    relay_conn far_4_4930_1_a(.in(far_4_4930_0[0]), .out(far_4_4930_1[0]));    relay_conn far_4_4930_1_b(.in(far_4_4930_0[1]), .out(far_4_4930_1[1]));
    assign layer_4[850] = far_4_4930_1[1] & ~far_4_4930_1[0]; 
    wire [1:0] far_4_4931_0;    relay_conn far_4_4931_0_a(.in(layer_3[656]), .out(far_4_4931_0[0]));    relay_conn far_4_4931_0_b(.in(layer_3[558]), .out(far_4_4931_0[1]));
    wire [1:0] far_4_4931_1;    relay_conn far_4_4931_1_a(.in(far_4_4931_0[0]), .out(far_4_4931_1[0]));    relay_conn far_4_4931_1_b(.in(far_4_4931_0[1]), .out(far_4_4931_1[1]));
    wire [1:0] far_4_4931_2;    relay_conn far_4_4931_2_a(.in(far_4_4931_1[0]), .out(far_4_4931_2[0]));    relay_conn far_4_4931_2_b(.in(far_4_4931_1[1]), .out(far_4_4931_2[1]));
    assign layer_4[851] = far_4_4931_2[0]; 
    wire [1:0] far_4_4932_0;    relay_conn far_4_4932_0_a(.in(layer_3[850]), .out(far_4_4932_0[0]));    relay_conn far_4_4932_0_b(.in(layer_3[744]), .out(far_4_4932_0[1]));
    wire [1:0] far_4_4932_1;    relay_conn far_4_4932_1_a(.in(far_4_4932_0[0]), .out(far_4_4932_1[0]));    relay_conn far_4_4932_1_b(.in(far_4_4932_0[1]), .out(far_4_4932_1[1]));
    wire [1:0] far_4_4932_2;    relay_conn far_4_4932_2_a(.in(far_4_4932_1[0]), .out(far_4_4932_2[0]));    relay_conn far_4_4932_2_b(.in(far_4_4932_1[1]), .out(far_4_4932_2[1]));
    assign layer_4[852] = far_4_4932_2[0] | far_4_4932_2[1]; 
    wire [1:0] far_4_4933_0;    relay_conn far_4_4933_0_a(.in(layer_3[637]), .out(far_4_4933_0[0]));    relay_conn far_4_4933_0_b(.in(layer_3[511]), .out(far_4_4933_0[1]));
    wire [1:0] far_4_4933_1;    relay_conn far_4_4933_1_a(.in(far_4_4933_0[0]), .out(far_4_4933_1[0]));    relay_conn far_4_4933_1_b(.in(far_4_4933_0[1]), .out(far_4_4933_1[1]));
    wire [1:0] far_4_4933_2;    relay_conn far_4_4933_2_a(.in(far_4_4933_1[0]), .out(far_4_4933_2[0]));    relay_conn far_4_4933_2_b(.in(far_4_4933_1[1]), .out(far_4_4933_2[1]));
    assign layer_4[853] = far_4_4933_2[0] ^ far_4_4933_2[1]; 
    wire [1:0] far_4_4934_0;    relay_conn far_4_4934_0_a(.in(layer_3[261]), .out(far_4_4934_0[0]));    relay_conn far_4_4934_0_b(.in(layer_3[386]), .out(far_4_4934_0[1]));
    wire [1:0] far_4_4934_1;    relay_conn far_4_4934_1_a(.in(far_4_4934_0[0]), .out(far_4_4934_1[0]));    relay_conn far_4_4934_1_b(.in(far_4_4934_0[1]), .out(far_4_4934_1[1]));
    wire [1:0] far_4_4934_2;    relay_conn far_4_4934_2_a(.in(far_4_4934_1[0]), .out(far_4_4934_2[0]));    relay_conn far_4_4934_2_b(.in(far_4_4934_1[1]), .out(far_4_4934_2[1]));
    assign layer_4[854] = far_4_4934_2[0]; 
    wire [1:0] far_4_4935_0;    relay_conn far_4_4935_0_a(.in(layer_3[329]), .out(far_4_4935_0[0]));    relay_conn far_4_4935_0_b(.in(layer_3[422]), .out(far_4_4935_0[1]));
    wire [1:0] far_4_4935_1;    relay_conn far_4_4935_1_a(.in(far_4_4935_0[0]), .out(far_4_4935_1[0]));    relay_conn far_4_4935_1_b(.in(far_4_4935_0[1]), .out(far_4_4935_1[1]));
    assign layer_4[855] = far_4_4935_1[0]; 
    wire [1:0] far_4_4936_0;    relay_conn far_4_4936_0_a(.in(layer_3[939]), .out(far_4_4936_0[0]));    relay_conn far_4_4936_0_b(.in(layer_3[850]), .out(far_4_4936_0[1]));
    wire [1:0] far_4_4936_1;    relay_conn far_4_4936_1_a(.in(far_4_4936_0[0]), .out(far_4_4936_1[0]));    relay_conn far_4_4936_1_b(.in(far_4_4936_0[1]), .out(far_4_4936_1[1]));
    assign layer_4[856] = ~(far_4_4936_1[0] & far_4_4936_1[1]); 
    assign layer_4[857] = layer_3[220] & layer_3[199]; 
    wire [1:0] far_4_4938_0;    relay_conn far_4_4938_0_a(.in(layer_3[896]), .out(far_4_4938_0[0]));    relay_conn far_4_4938_0_b(.in(layer_3[859]), .out(far_4_4938_0[1]));
    assign layer_4[858] = far_4_4938_0[0]; 
    wire [1:0] far_4_4939_0;    relay_conn far_4_4939_0_a(.in(layer_3[674]), .out(far_4_4939_0[0]));    relay_conn far_4_4939_0_b(.in(layer_3[615]), .out(far_4_4939_0[1]));
    assign layer_4[859] = far_4_4939_0[0] ^ far_4_4939_0[1]; 
    wire [1:0] far_4_4940_0;    relay_conn far_4_4940_0_a(.in(layer_3[263]), .out(far_4_4940_0[0]));    relay_conn far_4_4940_0_b(.in(layer_3[376]), .out(far_4_4940_0[1]));
    wire [1:0] far_4_4940_1;    relay_conn far_4_4940_1_a(.in(far_4_4940_0[0]), .out(far_4_4940_1[0]));    relay_conn far_4_4940_1_b(.in(far_4_4940_0[1]), .out(far_4_4940_1[1]));
    wire [1:0] far_4_4940_2;    relay_conn far_4_4940_2_a(.in(far_4_4940_1[0]), .out(far_4_4940_2[0]));    relay_conn far_4_4940_2_b(.in(far_4_4940_1[1]), .out(far_4_4940_2[1]));
    assign layer_4[860] = ~far_4_4940_2[0] | (far_4_4940_2[0] & far_4_4940_2[1]); 
    wire [1:0] far_4_4941_0;    relay_conn far_4_4941_0_a(.in(layer_3[848]), .out(far_4_4941_0[0]));    relay_conn far_4_4941_0_b(.in(layer_3[778]), .out(far_4_4941_0[1]));
    wire [1:0] far_4_4941_1;    relay_conn far_4_4941_1_a(.in(far_4_4941_0[0]), .out(far_4_4941_1[0]));    relay_conn far_4_4941_1_b(.in(far_4_4941_0[1]), .out(far_4_4941_1[1]));
    assign layer_4[861] = ~far_4_4941_1[1]; 
    wire [1:0] far_4_4942_0;    relay_conn far_4_4942_0_a(.in(layer_3[352]), .out(far_4_4942_0[0]));    relay_conn far_4_4942_0_b(.in(layer_3[467]), .out(far_4_4942_0[1]));
    wire [1:0] far_4_4942_1;    relay_conn far_4_4942_1_a(.in(far_4_4942_0[0]), .out(far_4_4942_1[0]));    relay_conn far_4_4942_1_b(.in(far_4_4942_0[1]), .out(far_4_4942_1[1]));
    wire [1:0] far_4_4942_2;    relay_conn far_4_4942_2_a(.in(far_4_4942_1[0]), .out(far_4_4942_2[0]));    relay_conn far_4_4942_2_b(.in(far_4_4942_1[1]), .out(far_4_4942_2[1]));
    assign layer_4[862] = ~far_4_4942_2[1]; 
    wire [1:0] far_4_4943_0;    relay_conn far_4_4943_0_a(.in(layer_3[761]), .out(far_4_4943_0[0]));    relay_conn far_4_4943_0_b(.in(layer_3[884]), .out(far_4_4943_0[1]));
    wire [1:0] far_4_4943_1;    relay_conn far_4_4943_1_a(.in(far_4_4943_0[0]), .out(far_4_4943_1[0]));    relay_conn far_4_4943_1_b(.in(far_4_4943_0[1]), .out(far_4_4943_1[1]));
    wire [1:0] far_4_4943_2;    relay_conn far_4_4943_2_a(.in(far_4_4943_1[0]), .out(far_4_4943_2[0]));    relay_conn far_4_4943_2_b(.in(far_4_4943_1[1]), .out(far_4_4943_2[1]));
    assign layer_4[863] = ~far_4_4943_2[0]; 
    wire [1:0] far_4_4944_0;    relay_conn far_4_4944_0_a(.in(layer_3[868]), .out(far_4_4944_0[0]));    relay_conn far_4_4944_0_b(.in(layer_3[953]), .out(far_4_4944_0[1]));
    wire [1:0] far_4_4944_1;    relay_conn far_4_4944_1_a(.in(far_4_4944_0[0]), .out(far_4_4944_1[0]));    relay_conn far_4_4944_1_b(.in(far_4_4944_0[1]), .out(far_4_4944_1[1]));
    assign layer_4[864] = ~far_4_4944_1[1]; 
    wire [1:0] far_4_4945_0;    relay_conn far_4_4945_0_a(.in(layer_3[561]), .out(far_4_4945_0[0]));    relay_conn far_4_4945_0_b(.in(layer_3[475]), .out(far_4_4945_0[1]));
    wire [1:0] far_4_4945_1;    relay_conn far_4_4945_1_a(.in(far_4_4945_0[0]), .out(far_4_4945_1[0]));    relay_conn far_4_4945_1_b(.in(far_4_4945_0[1]), .out(far_4_4945_1[1]));
    assign layer_4[865] = ~far_4_4945_1[0]; 
    wire [1:0] far_4_4946_0;    relay_conn far_4_4946_0_a(.in(layer_3[838]), .out(far_4_4946_0[0]));    relay_conn far_4_4946_0_b(.in(layer_3[953]), .out(far_4_4946_0[1]));
    wire [1:0] far_4_4946_1;    relay_conn far_4_4946_1_a(.in(far_4_4946_0[0]), .out(far_4_4946_1[0]));    relay_conn far_4_4946_1_b(.in(far_4_4946_0[1]), .out(far_4_4946_1[1]));
    wire [1:0] far_4_4946_2;    relay_conn far_4_4946_2_a(.in(far_4_4946_1[0]), .out(far_4_4946_2[0]));    relay_conn far_4_4946_2_b(.in(far_4_4946_1[1]), .out(far_4_4946_2[1]));
    assign layer_4[866] = ~far_4_4946_2[0]; 
    wire [1:0] far_4_4947_0;    relay_conn far_4_4947_0_a(.in(layer_3[837]), .out(far_4_4947_0[0]));    relay_conn far_4_4947_0_b(.in(layer_3[958]), .out(far_4_4947_0[1]));
    wire [1:0] far_4_4947_1;    relay_conn far_4_4947_1_a(.in(far_4_4947_0[0]), .out(far_4_4947_1[0]));    relay_conn far_4_4947_1_b(.in(far_4_4947_0[1]), .out(far_4_4947_1[1]));
    wire [1:0] far_4_4947_2;    relay_conn far_4_4947_2_a(.in(far_4_4947_1[0]), .out(far_4_4947_2[0]));    relay_conn far_4_4947_2_b(.in(far_4_4947_1[1]), .out(far_4_4947_2[1]));
    assign layer_4[867] = ~far_4_4947_2[0]; 
    wire [1:0] far_4_4948_0;    relay_conn far_4_4948_0_a(.in(layer_3[270]), .out(far_4_4948_0[0]));    relay_conn far_4_4948_0_b(.in(layer_3[328]), .out(far_4_4948_0[1]));
    assign layer_4[868] = ~far_4_4948_0[1]; 
    assign layer_4[869] = layer_3[930]; 
    wire [1:0] far_4_4950_0;    relay_conn far_4_4950_0_a(.in(layer_3[312]), .out(far_4_4950_0[0]));    relay_conn far_4_4950_0_b(.in(layer_3[364]), .out(far_4_4950_0[1]));
    assign layer_4[870] = ~far_4_4950_0[1]; 
    wire [1:0] far_4_4951_0;    relay_conn far_4_4951_0_a(.in(layer_3[569]), .out(far_4_4951_0[0]));    relay_conn far_4_4951_0_b(.in(layer_3[694]), .out(far_4_4951_0[1]));
    wire [1:0] far_4_4951_1;    relay_conn far_4_4951_1_a(.in(far_4_4951_0[0]), .out(far_4_4951_1[0]));    relay_conn far_4_4951_1_b(.in(far_4_4951_0[1]), .out(far_4_4951_1[1]));
    wire [1:0] far_4_4951_2;    relay_conn far_4_4951_2_a(.in(far_4_4951_1[0]), .out(far_4_4951_2[0]));    relay_conn far_4_4951_2_b(.in(far_4_4951_1[1]), .out(far_4_4951_2[1]));
    assign layer_4[871] = ~far_4_4951_2[0]; 
    wire [1:0] far_4_4952_0;    relay_conn far_4_4952_0_a(.in(layer_3[818]), .out(far_4_4952_0[0]));    relay_conn far_4_4952_0_b(.in(layer_3[770]), .out(far_4_4952_0[1]));
    assign layer_4[872] = far_4_4952_0[0]; 
    wire [1:0] far_4_4953_0;    relay_conn far_4_4953_0_a(.in(layer_3[155]), .out(far_4_4953_0[0]));    relay_conn far_4_4953_0_b(.in(layer_3[242]), .out(far_4_4953_0[1]));
    wire [1:0] far_4_4953_1;    relay_conn far_4_4953_1_a(.in(far_4_4953_0[0]), .out(far_4_4953_1[0]));    relay_conn far_4_4953_1_b(.in(far_4_4953_0[1]), .out(far_4_4953_1[1]));
    assign layer_4[873] = ~far_4_4953_1[0]; 
    wire [1:0] far_4_4954_0;    relay_conn far_4_4954_0_a(.in(layer_3[692]), .out(far_4_4954_0[0]));    relay_conn far_4_4954_0_b(.in(layer_3[569]), .out(far_4_4954_0[1]));
    wire [1:0] far_4_4954_1;    relay_conn far_4_4954_1_a(.in(far_4_4954_0[0]), .out(far_4_4954_1[0]));    relay_conn far_4_4954_1_b(.in(far_4_4954_0[1]), .out(far_4_4954_1[1]));
    wire [1:0] far_4_4954_2;    relay_conn far_4_4954_2_a(.in(far_4_4954_1[0]), .out(far_4_4954_2[0]));    relay_conn far_4_4954_2_b(.in(far_4_4954_1[1]), .out(far_4_4954_2[1]));
    assign layer_4[874] = far_4_4954_2[1] & ~far_4_4954_2[0]; 
    assign layer_4[875] = layer_3[709] & ~layer_3[680]; 
    wire [1:0] far_4_4956_0;    relay_conn far_4_4956_0_a(.in(layer_3[365]), .out(far_4_4956_0[0]));    relay_conn far_4_4956_0_b(.in(layer_3[275]), .out(far_4_4956_0[1]));
    wire [1:0] far_4_4956_1;    relay_conn far_4_4956_1_a(.in(far_4_4956_0[0]), .out(far_4_4956_1[0]));    relay_conn far_4_4956_1_b(.in(far_4_4956_0[1]), .out(far_4_4956_1[1]));
    assign layer_4[876] = far_4_4956_1[0]; 
    assign layer_4[877] = ~layer_3[674] | (layer_3[649] & layer_3[674]); 
    wire [1:0] far_4_4958_0;    relay_conn far_4_4958_0_a(.in(layer_3[212]), .out(far_4_4958_0[0]));    relay_conn far_4_4958_0_b(.in(layer_3[274]), .out(far_4_4958_0[1]));
    assign layer_4[878] = ~(far_4_4958_0[0] & far_4_4958_0[1]); 
    wire [1:0] far_4_4959_0;    relay_conn far_4_4959_0_a(.in(layer_3[410]), .out(far_4_4959_0[0]));    relay_conn far_4_4959_0_b(.in(layer_3[451]), .out(far_4_4959_0[1]));
    assign layer_4[879] = far_4_4959_0[1] & ~far_4_4959_0[0]; 
    wire [1:0] far_4_4960_0;    relay_conn far_4_4960_0_a(.in(layer_3[35]), .out(far_4_4960_0[0]));    relay_conn far_4_4960_0_b(.in(layer_3[127]), .out(far_4_4960_0[1]));
    wire [1:0] far_4_4960_1;    relay_conn far_4_4960_1_a(.in(far_4_4960_0[0]), .out(far_4_4960_1[0]));    relay_conn far_4_4960_1_b(.in(far_4_4960_0[1]), .out(far_4_4960_1[1]));
    assign layer_4[880] = ~(far_4_4960_1[0] & far_4_4960_1[1]); 
    wire [1:0] far_4_4961_0;    relay_conn far_4_4961_0_a(.in(layer_3[939]), .out(far_4_4961_0[0]));    relay_conn far_4_4961_0_b(.in(layer_3[874]), .out(far_4_4961_0[1]));
    wire [1:0] far_4_4961_1;    relay_conn far_4_4961_1_a(.in(far_4_4961_0[0]), .out(far_4_4961_1[0]));    relay_conn far_4_4961_1_b(.in(far_4_4961_0[1]), .out(far_4_4961_1[1]));
    assign layer_4[881] = far_4_4961_1[1]; 
    assign layer_4[882] = layer_3[673] & layer_3[644]; 
    wire [1:0] far_4_4963_0;    relay_conn far_4_4963_0_a(.in(layer_3[37]), .out(far_4_4963_0[0]));    relay_conn far_4_4963_0_b(.in(layer_3[149]), .out(far_4_4963_0[1]));
    wire [1:0] far_4_4963_1;    relay_conn far_4_4963_1_a(.in(far_4_4963_0[0]), .out(far_4_4963_1[0]));    relay_conn far_4_4963_1_b(.in(far_4_4963_0[1]), .out(far_4_4963_1[1]));
    wire [1:0] far_4_4963_2;    relay_conn far_4_4963_2_a(.in(far_4_4963_1[0]), .out(far_4_4963_2[0]));    relay_conn far_4_4963_2_b(.in(far_4_4963_1[1]), .out(far_4_4963_2[1]));
    assign layer_4[883] = ~(far_4_4963_2[0] ^ far_4_4963_2[1]); 
    wire [1:0] far_4_4964_0;    relay_conn far_4_4964_0_a(.in(layer_3[664]), .out(far_4_4964_0[0]));    relay_conn far_4_4964_0_b(.in(layer_3[568]), .out(far_4_4964_0[1]));
    wire [1:0] far_4_4964_1;    relay_conn far_4_4964_1_a(.in(far_4_4964_0[0]), .out(far_4_4964_1[0]));    relay_conn far_4_4964_1_b(.in(far_4_4964_0[1]), .out(far_4_4964_1[1]));
    wire [1:0] far_4_4964_2;    relay_conn far_4_4964_2_a(.in(far_4_4964_1[0]), .out(far_4_4964_2[0]));    relay_conn far_4_4964_2_b(.in(far_4_4964_1[1]), .out(far_4_4964_2[1]));
    assign layer_4[884] = ~far_4_4964_2[1]; 
    wire [1:0] far_4_4965_0;    relay_conn far_4_4965_0_a(.in(layer_3[524]), .out(far_4_4965_0[0]));    relay_conn far_4_4965_0_b(.in(layer_3[612]), .out(far_4_4965_0[1]));
    wire [1:0] far_4_4965_1;    relay_conn far_4_4965_1_a(.in(far_4_4965_0[0]), .out(far_4_4965_1[0]));    relay_conn far_4_4965_1_b(.in(far_4_4965_0[1]), .out(far_4_4965_1[1]));
    assign layer_4[885] = far_4_4965_1[1]; 
    wire [1:0] far_4_4966_0;    relay_conn far_4_4966_0_a(.in(layer_3[766]), .out(far_4_4966_0[0]));    relay_conn far_4_4966_0_b(.in(layer_3[829]), .out(far_4_4966_0[1]));
    assign layer_4[886] = ~far_4_4966_0[0]; 
    wire [1:0] far_4_4967_0;    relay_conn far_4_4967_0_a(.in(layer_3[236]), .out(far_4_4967_0[0]));    relay_conn far_4_4967_0_b(.in(layer_3[268]), .out(far_4_4967_0[1]));
    assign layer_4[887] = far_4_4967_0[0] & far_4_4967_0[1]; 
    wire [1:0] far_4_4968_0;    relay_conn far_4_4968_0_a(.in(layer_3[942]), .out(far_4_4968_0[0]));    relay_conn far_4_4968_0_b(.in(layer_3[846]), .out(far_4_4968_0[1]));
    wire [1:0] far_4_4968_1;    relay_conn far_4_4968_1_a(.in(far_4_4968_0[0]), .out(far_4_4968_1[0]));    relay_conn far_4_4968_1_b(.in(far_4_4968_0[1]), .out(far_4_4968_1[1]));
    wire [1:0] far_4_4968_2;    relay_conn far_4_4968_2_a(.in(far_4_4968_1[0]), .out(far_4_4968_2[0]));    relay_conn far_4_4968_2_b(.in(far_4_4968_1[1]), .out(far_4_4968_2[1]));
    assign layer_4[888] = far_4_4968_2[0] & far_4_4968_2[1]; 
    wire [1:0] far_4_4969_0;    relay_conn far_4_4969_0_a(.in(layer_3[630]), .out(far_4_4969_0[0]));    relay_conn far_4_4969_0_b(.in(layer_3[577]), .out(far_4_4969_0[1]));
    assign layer_4[889] = ~(far_4_4969_0[0] & far_4_4969_0[1]); 
    assign layer_4[890] = ~layer_3[805]; 
    wire [1:0] far_4_4971_0;    relay_conn far_4_4971_0_a(.in(layer_3[428]), .out(far_4_4971_0[0]));    relay_conn far_4_4971_0_b(.in(layer_3[504]), .out(far_4_4971_0[1]));
    wire [1:0] far_4_4971_1;    relay_conn far_4_4971_1_a(.in(far_4_4971_0[0]), .out(far_4_4971_1[0]));    relay_conn far_4_4971_1_b(.in(far_4_4971_0[1]), .out(far_4_4971_1[1]));
    assign layer_4[891] = far_4_4971_1[0] | far_4_4971_1[1]; 
    wire [1:0] far_4_4972_0;    relay_conn far_4_4972_0_a(.in(layer_3[780]), .out(far_4_4972_0[0]));    relay_conn far_4_4972_0_b(.in(layer_3[855]), .out(far_4_4972_0[1]));
    wire [1:0] far_4_4972_1;    relay_conn far_4_4972_1_a(.in(far_4_4972_0[0]), .out(far_4_4972_1[0]));    relay_conn far_4_4972_1_b(.in(far_4_4972_0[1]), .out(far_4_4972_1[1]));
    assign layer_4[892] = far_4_4972_1[1] & ~far_4_4972_1[0]; 
    assign layer_4[893] = layer_3[906]; 
    wire [1:0] far_4_4974_0;    relay_conn far_4_4974_0_a(.in(layer_3[169]), .out(far_4_4974_0[0]));    relay_conn far_4_4974_0_b(.in(layer_3[118]), .out(far_4_4974_0[1]));
    assign layer_4[894] = far_4_4974_0[0] & ~far_4_4974_0[1]; 
    assign layer_4[895] = layer_3[876]; 
    wire [1:0] far_4_4976_0;    relay_conn far_4_4976_0_a(.in(layer_3[478]), .out(far_4_4976_0[0]));    relay_conn far_4_4976_0_b(.in(layer_3[443]), .out(far_4_4976_0[1]));
    assign layer_4[896] = far_4_4976_0[1] & ~far_4_4976_0[0]; 
    wire [1:0] far_4_4977_0;    relay_conn far_4_4977_0_a(.in(layer_3[632]), .out(far_4_4977_0[0]));    relay_conn far_4_4977_0_b(.in(layer_3[727]), .out(far_4_4977_0[1]));
    wire [1:0] far_4_4977_1;    relay_conn far_4_4977_1_a(.in(far_4_4977_0[0]), .out(far_4_4977_1[0]));    relay_conn far_4_4977_1_b(.in(far_4_4977_0[1]), .out(far_4_4977_1[1]));
    assign layer_4[897] = ~far_4_4977_1[0] | (far_4_4977_1[0] & far_4_4977_1[1]); 
    wire [1:0] far_4_4978_0;    relay_conn far_4_4978_0_a(.in(layer_3[100]), .out(far_4_4978_0[0]));    relay_conn far_4_4978_0_b(.in(layer_3[35]), .out(far_4_4978_0[1]));
    wire [1:0] far_4_4978_1;    relay_conn far_4_4978_1_a(.in(far_4_4978_0[0]), .out(far_4_4978_1[0]));    relay_conn far_4_4978_1_b(.in(far_4_4978_0[1]), .out(far_4_4978_1[1]));
    assign layer_4[898] = far_4_4978_1[0] & ~far_4_4978_1[1]; 
    assign layer_4[899] = ~(layer_3[15] | layer_3[39]); 
    wire [1:0] far_4_4980_0;    relay_conn far_4_4980_0_a(.in(layer_3[517]), .out(far_4_4980_0[0]));    relay_conn far_4_4980_0_b(.in(layer_3[475]), .out(far_4_4980_0[1]));
    assign layer_4[900] = ~far_4_4980_0[0] | (far_4_4980_0[0] & far_4_4980_0[1]); 
    assign layer_4[901] = layer_3[778] & ~layer_3[761]; 
    assign layer_4[902] = ~layer_3[289]; 
    assign layer_4[903] = layer_3[553] & ~layer_3[556]; 
    wire [1:0] far_4_4984_0;    relay_conn far_4_4984_0_a(.in(layer_3[190]), .out(far_4_4984_0[0]));    relay_conn far_4_4984_0_b(.in(layer_3[297]), .out(far_4_4984_0[1]));
    wire [1:0] far_4_4984_1;    relay_conn far_4_4984_1_a(.in(far_4_4984_0[0]), .out(far_4_4984_1[0]));    relay_conn far_4_4984_1_b(.in(far_4_4984_0[1]), .out(far_4_4984_1[1]));
    wire [1:0] far_4_4984_2;    relay_conn far_4_4984_2_a(.in(far_4_4984_1[0]), .out(far_4_4984_2[0]));    relay_conn far_4_4984_2_b(.in(far_4_4984_1[1]), .out(far_4_4984_2[1]));
    assign layer_4[904] = ~(far_4_4984_2[0] & far_4_4984_2[1]); 
    assign layer_4[905] = layer_3[672]; 
    assign layer_4[906] = layer_3[275] & ~layer_3[284]; 
    assign layer_4[907] = layer_3[436] & ~layer_3[455]; 
    wire [1:0] far_4_4988_0;    relay_conn far_4_4988_0_a(.in(layer_3[243]), .out(far_4_4988_0[0]));    relay_conn far_4_4988_0_b(.in(layer_3[126]), .out(far_4_4988_0[1]));
    wire [1:0] far_4_4988_1;    relay_conn far_4_4988_1_a(.in(far_4_4988_0[0]), .out(far_4_4988_1[0]));    relay_conn far_4_4988_1_b(.in(far_4_4988_0[1]), .out(far_4_4988_1[1]));
    wire [1:0] far_4_4988_2;    relay_conn far_4_4988_2_a(.in(far_4_4988_1[0]), .out(far_4_4988_2[0]));    relay_conn far_4_4988_2_b(.in(far_4_4988_1[1]), .out(far_4_4988_2[1]));
    assign layer_4[908] = far_4_4988_2[1] & ~far_4_4988_2[0]; 
    wire [1:0] far_4_4989_0;    relay_conn far_4_4989_0_a(.in(layer_3[361]), .out(far_4_4989_0[0]));    relay_conn far_4_4989_0_b(.in(layer_3[253]), .out(far_4_4989_0[1]));
    wire [1:0] far_4_4989_1;    relay_conn far_4_4989_1_a(.in(far_4_4989_0[0]), .out(far_4_4989_1[0]));    relay_conn far_4_4989_1_b(.in(far_4_4989_0[1]), .out(far_4_4989_1[1]));
    wire [1:0] far_4_4989_2;    relay_conn far_4_4989_2_a(.in(far_4_4989_1[0]), .out(far_4_4989_2[0]));    relay_conn far_4_4989_2_b(.in(far_4_4989_1[1]), .out(far_4_4989_2[1]));
    assign layer_4[909] = ~(far_4_4989_2[0] ^ far_4_4989_2[1]); 
    wire [1:0] far_4_4990_0;    relay_conn far_4_4990_0_a(.in(layer_3[462]), .out(far_4_4990_0[0]));    relay_conn far_4_4990_0_b(.in(layer_3[398]), .out(far_4_4990_0[1]));
    wire [1:0] far_4_4990_1;    relay_conn far_4_4990_1_a(.in(far_4_4990_0[0]), .out(far_4_4990_1[0]));    relay_conn far_4_4990_1_b(.in(far_4_4990_0[1]), .out(far_4_4990_1[1]));
    assign layer_4[910] = ~far_4_4990_1[0] | (far_4_4990_1[0] & far_4_4990_1[1]); 
    wire [1:0] far_4_4991_0;    relay_conn far_4_4991_0_a(.in(layer_3[255]), .out(far_4_4991_0[0]));    relay_conn far_4_4991_0_b(.in(layer_3[140]), .out(far_4_4991_0[1]));
    wire [1:0] far_4_4991_1;    relay_conn far_4_4991_1_a(.in(far_4_4991_0[0]), .out(far_4_4991_1[0]));    relay_conn far_4_4991_1_b(.in(far_4_4991_0[1]), .out(far_4_4991_1[1]));
    wire [1:0] far_4_4991_2;    relay_conn far_4_4991_2_a(.in(far_4_4991_1[0]), .out(far_4_4991_2[0]));    relay_conn far_4_4991_2_b(.in(far_4_4991_1[1]), .out(far_4_4991_2[1]));
    assign layer_4[911] = far_4_4991_2[0] | far_4_4991_2[1]; 
    wire [1:0] far_4_4992_0;    relay_conn far_4_4992_0_a(.in(layer_3[829]), .out(far_4_4992_0[0]));    relay_conn far_4_4992_0_b(.in(layer_3[764]), .out(far_4_4992_0[1]));
    wire [1:0] far_4_4992_1;    relay_conn far_4_4992_1_a(.in(far_4_4992_0[0]), .out(far_4_4992_1[0]));    relay_conn far_4_4992_1_b(.in(far_4_4992_0[1]), .out(far_4_4992_1[1]));
    assign layer_4[912] = far_4_4992_1[1] & ~far_4_4992_1[0]; 
    wire [1:0] far_4_4993_0;    relay_conn far_4_4993_0_a(.in(layer_3[567]), .out(far_4_4993_0[0]));    relay_conn far_4_4993_0_b(.in(layer_3[443]), .out(far_4_4993_0[1]));
    wire [1:0] far_4_4993_1;    relay_conn far_4_4993_1_a(.in(far_4_4993_0[0]), .out(far_4_4993_1[0]));    relay_conn far_4_4993_1_b(.in(far_4_4993_0[1]), .out(far_4_4993_1[1]));
    wire [1:0] far_4_4993_2;    relay_conn far_4_4993_2_a(.in(far_4_4993_1[0]), .out(far_4_4993_2[0]));    relay_conn far_4_4993_2_b(.in(far_4_4993_1[1]), .out(far_4_4993_2[1]));
    assign layer_4[913] = ~far_4_4993_2[0] | (far_4_4993_2[0] & far_4_4993_2[1]); 
    wire [1:0] far_4_4994_0;    relay_conn far_4_4994_0_a(.in(layer_3[477]), .out(far_4_4994_0[0]));    relay_conn far_4_4994_0_b(.in(layer_3[593]), .out(far_4_4994_0[1]));
    wire [1:0] far_4_4994_1;    relay_conn far_4_4994_1_a(.in(far_4_4994_0[0]), .out(far_4_4994_1[0]));    relay_conn far_4_4994_1_b(.in(far_4_4994_0[1]), .out(far_4_4994_1[1]));
    wire [1:0] far_4_4994_2;    relay_conn far_4_4994_2_a(.in(far_4_4994_1[0]), .out(far_4_4994_2[0]));    relay_conn far_4_4994_2_b(.in(far_4_4994_1[1]), .out(far_4_4994_2[1]));
    assign layer_4[914] = far_4_4994_2[0]; 
    wire [1:0] far_4_4995_0;    relay_conn far_4_4995_0_a(.in(layer_3[636]), .out(far_4_4995_0[0]));    relay_conn far_4_4995_0_b(.in(layer_3[676]), .out(far_4_4995_0[1]));
    assign layer_4[915] = far_4_4995_0[1] & ~far_4_4995_0[0]; 
    wire [1:0] far_4_4996_0;    relay_conn far_4_4996_0_a(.in(layer_3[1009]), .out(far_4_4996_0[0]));    relay_conn far_4_4996_0_b(.in(layer_3[916]), .out(far_4_4996_0[1]));
    wire [1:0] far_4_4996_1;    relay_conn far_4_4996_1_a(.in(far_4_4996_0[0]), .out(far_4_4996_1[0]));    relay_conn far_4_4996_1_b(.in(far_4_4996_0[1]), .out(far_4_4996_1[1]));
    assign layer_4[916] = far_4_4996_1[0] | far_4_4996_1[1]; 
    wire [1:0] far_4_4997_0;    relay_conn far_4_4997_0_a(.in(layer_3[883]), .out(far_4_4997_0[0]));    relay_conn far_4_4997_0_b(.in(layer_3[788]), .out(far_4_4997_0[1]));
    wire [1:0] far_4_4997_1;    relay_conn far_4_4997_1_a(.in(far_4_4997_0[0]), .out(far_4_4997_1[0]));    relay_conn far_4_4997_1_b(.in(far_4_4997_0[1]), .out(far_4_4997_1[1]));
    assign layer_4[917] = far_4_4997_1[0] & ~far_4_4997_1[1]; 
    wire [1:0] far_4_4998_0;    relay_conn far_4_4998_0_a(.in(layer_3[281]), .out(far_4_4998_0[0]));    relay_conn far_4_4998_0_b(.in(layer_3[317]), .out(far_4_4998_0[1]));
    assign layer_4[918] = ~far_4_4998_0[0] | (far_4_4998_0[0] & far_4_4998_0[1]); 
    wire [1:0] far_4_4999_0;    relay_conn far_4_4999_0_a(.in(layer_3[414]), .out(far_4_4999_0[0]));    relay_conn far_4_4999_0_b(.in(layer_3[367]), .out(far_4_4999_0[1]));
    assign layer_4[919] = ~(far_4_4999_0[0] ^ far_4_4999_0[1]); 
    wire [1:0] far_4_5000_0;    relay_conn far_4_5000_0_a(.in(layer_3[950]), .out(far_4_5000_0[0]));    relay_conn far_4_5000_0_b(.in(layer_3[1010]), .out(far_4_5000_0[1]));
    assign layer_4[920] = far_4_5000_0[0]; 
    wire [1:0] far_4_5001_0;    relay_conn far_4_5001_0_a(.in(layer_3[384]), .out(far_4_5001_0[0]));    relay_conn far_4_5001_0_b(.in(layer_3[350]), .out(far_4_5001_0[1]));
    assign layer_4[921] = far_4_5001_0[1]; 
    wire [1:0] far_4_5002_0;    relay_conn far_4_5002_0_a(.in(layer_3[562]), .out(far_4_5002_0[0]));    relay_conn far_4_5002_0_b(.in(layer_3[457]), .out(far_4_5002_0[1]));
    wire [1:0] far_4_5002_1;    relay_conn far_4_5002_1_a(.in(far_4_5002_0[0]), .out(far_4_5002_1[0]));    relay_conn far_4_5002_1_b(.in(far_4_5002_0[1]), .out(far_4_5002_1[1]));
    wire [1:0] far_4_5002_2;    relay_conn far_4_5002_2_a(.in(far_4_5002_1[0]), .out(far_4_5002_2[0]));    relay_conn far_4_5002_2_b(.in(far_4_5002_1[1]), .out(far_4_5002_2[1]));
    assign layer_4[922] = far_4_5002_2[0]; 
    wire [1:0] far_4_5003_0;    relay_conn far_4_5003_0_a(.in(layer_3[596]), .out(far_4_5003_0[0]));    relay_conn far_4_5003_0_b(.in(layer_3[630]), .out(far_4_5003_0[1]));
    assign layer_4[923] = far_4_5003_0[1]; 
    wire [1:0] far_4_5004_0;    relay_conn far_4_5004_0_a(.in(layer_3[497]), .out(far_4_5004_0[0]));    relay_conn far_4_5004_0_b(.in(layer_3[434]), .out(far_4_5004_0[1]));
    assign layer_4[924] = ~far_4_5004_0[0]; 
    wire [1:0] far_4_5005_0;    relay_conn far_4_5005_0_a(.in(layer_3[104]), .out(far_4_5005_0[0]));    relay_conn far_4_5005_0_b(.in(layer_3[35]), .out(far_4_5005_0[1]));
    wire [1:0] far_4_5005_1;    relay_conn far_4_5005_1_a(.in(far_4_5005_0[0]), .out(far_4_5005_1[0]));    relay_conn far_4_5005_1_b(.in(far_4_5005_0[1]), .out(far_4_5005_1[1]));
    assign layer_4[925] = far_4_5005_1[0] | far_4_5005_1[1]; 
    wire [1:0] far_4_5006_0;    relay_conn far_4_5006_0_a(.in(layer_3[563]), .out(far_4_5006_0[0]));    relay_conn far_4_5006_0_b(.in(layer_3[518]), .out(far_4_5006_0[1]));
    assign layer_4[926] = far_4_5006_0[1]; 
    assign layer_4[927] = ~layer_3[323] | (layer_3[323] & layer_3[352]); 
    wire [1:0] far_4_5008_0;    relay_conn far_4_5008_0_a(.in(layer_3[337]), .out(far_4_5008_0[0]));    relay_conn far_4_5008_0_b(.in(layer_3[440]), .out(far_4_5008_0[1]));
    wire [1:0] far_4_5008_1;    relay_conn far_4_5008_1_a(.in(far_4_5008_0[0]), .out(far_4_5008_1[0]));    relay_conn far_4_5008_1_b(.in(far_4_5008_0[1]), .out(far_4_5008_1[1]));
    wire [1:0] far_4_5008_2;    relay_conn far_4_5008_2_a(.in(far_4_5008_1[0]), .out(far_4_5008_2[0]));    relay_conn far_4_5008_2_b(.in(far_4_5008_1[1]), .out(far_4_5008_2[1]));
    assign layer_4[928] = ~far_4_5008_2[0]; 
    assign layer_4[929] = ~(layer_3[19] | layer_3[2]); 
    wire [1:0] far_4_5010_0;    relay_conn far_4_5010_0_a(.in(layer_3[749]), .out(far_4_5010_0[0]));    relay_conn far_4_5010_0_b(.in(layer_3[682]), .out(far_4_5010_0[1]));
    wire [1:0] far_4_5010_1;    relay_conn far_4_5010_1_a(.in(far_4_5010_0[0]), .out(far_4_5010_1[0]));    relay_conn far_4_5010_1_b(.in(far_4_5010_0[1]), .out(far_4_5010_1[1]));
    assign layer_4[930] = ~far_4_5010_1[1]; 
    wire [1:0] far_4_5011_0;    relay_conn far_4_5011_0_a(.in(layer_3[688]), .out(far_4_5011_0[0]));    relay_conn far_4_5011_0_b(.in(layer_3[772]), .out(far_4_5011_0[1]));
    wire [1:0] far_4_5011_1;    relay_conn far_4_5011_1_a(.in(far_4_5011_0[0]), .out(far_4_5011_1[0]));    relay_conn far_4_5011_1_b(.in(far_4_5011_0[1]), .out(far_4_5011_1[1]));
    assign layer_4[931] = ~(far_4_5011_1[0] | far_4_5011_1[1]); 
    wire [1:0] far_4_5012_0;    relay_conn far_4_5012_0_a(.in(layer_3[936]), .out(far_4_5012_0[0]));    relay_conn far_4_5012_0_b(.in(layer_3[972]), .out(far_4_5012_0[1]));
    assign layer_4[932] = ~far_4_5012_0[1]; 
    assign layer_4[933] = ~layer_3[146]; 
    wire [1:0] far_4_5014_0;    relay_conn far_4_5014_0_a(.in(layer_3[777]), .out(far_4_5014_0[0]));    relay_conn far_4_5014_0_b(.in(layer_3[676]), .out(far_4_5014_0[1]));
    wire [1:0] far_4_5014_1;    relay_conn far_4_5014_1_a(.in(far_4_5014_0[0]), .out(far_4_5014_1[0]));    relay_conn far_4_5014_1_b(.in(far_4_5014_0[1]), .out(far_4_5014_1[1]));
    wire [1:0] far_4_5014_2;    relay_conn far_4_5014_2_a(.in(far_4_5014_1[0]), .out(far_4_5014_2[0]));    relay_conn far_4_5014_2_b(.in(far_4_5014_1[1]), .out(far_4_5014_2[1]));
    assign layer_4[934] = far_4_5014_2[0] ^ far_4_5014_2[1]; 
    wire [1:0] far_4_5015_0;    relay_conn far_4_5015_0_a(.in(layer_3[873]), .out(far_4_5015_0[0]));    relay_conn far_4_5015_0_b(.in(layer_3[769]), .out(far_4_5015_0[1]));
    wire [1:0] far_4_5015_1;    relay_conn far_4_5015_1_a(.in(far_4_5015_0[0]), .out(far_4_5015_1[0]));    relay_conn far_4_5015_1_b(.in(far_4_5015_0[1]), .out(far_4_5015_1[1]));
    wire [1:0] far_4_5015_2;    relay_conn far_4_5015_2_a(.in(far_4_5015_1[0]), .out(far_4_5015_2[0]));    relay_conn far_4_5015_2_b(.in(far_4_5015_1[1]), .out(far_4_5015_2[1]));
    assign layer_4[935] = ~far_4_5015_2[1] | (far_4_5015_2[0] & far_4_5015_2[1]); 
    wire [1:0] far_4_5016_0;    relay_conn far_4_5016_0_a(.in(layer_3[50]), .out(far_4_5016_0[0]));    relay_conn far_4_5016_0_b(.in(layer_3[157]), .out(far_4_5016_0[1]));
    wire [1:0] far_4_5016_1;    relay_conn far_4_5016_1_a(.in(far_4_5016_0[0]), .out(far_4_5016_1[0]));    relay_conn far_4_5016_1_b(.in(far_4_5016_0[1]), .out(far_4_5016_1[1]));
    wire [1:0] far_4_5016_2;    relay_conn far_4_5016_2_a(.in(far_4_5016_1[0]), .out(far_4_5016_2[0]));    relay_conn far_4_5016_2_b(.in(far_4_5016_1[1]), .out(far_4_5016_2[1]));
    assign layer_4[936] = ~(far_4_5016_2[0] & far_4_5016_2[1]); 
    wire [1:0] far_4_5017_0;    relay_conn far_4_5017_0_a(.in(layer_3[353]), .out(far_4_5017_0[0]));    relay_conn far_4_5017_0_b(.in(layer_3[426]), .out(far_4_5017_0[1]));
    wire [1:0] far_4_5017_1;    relay_conn far_4_5017_1_a(.in(far_4_5017_0[0]), .out(far_4_5017_1[0]));    relay_conn far_4_5017_1_b(.in(far_4_5017_0[1]), .out(far_4_5017_1[1]));
    assign layer_4[937] = ~far_4_5017_1[0]; 
    wire [1:0] far_4_5018_0;    relay_conn far_4_5018_0_a(.in(layer_3[884]), .out(far_4_5018_0[0]));    relay_conn far_4_5018_0_b(.in(layer_3[802]), .out(far_4_5018_0[1]));
    wire [1:0] far_4_5018_1;    relay_conn far_4_5018_1_a(.in(far_4_5018_0[0]), .out(far_4_5018_1[0]));    relay_conn far_4_5018_1_b(.in(far_4_5018_0[1]), .out(far_4_5018_1[1]));
    assign layer_4[938] = ~far_4_5018_1[1]; 
    wire [1:0] far_4_5019_0;    relay_conn far_4_5019_0_a(.in(layer_3[65]), .out(far_4_5019_0[0]));    relay_conn far_4_5019_0_b(.in(layer_3[192]), .out(far_4_5019_0[1]));
    wire [1:0] far_4_5019_1;    relay_conn far_4_5019_1_a(.in(far_4_5019_0[0]), .out(far_4_5019_1[0]));    relay_conn far_4_5019_1_b(.in(far_4_5019_0[1]), .out(far_4_5019_1[1]));
    wire [1:0] far_4_5019_2;    relay_conn far_4_5019_2_a(.in(far_4_5019_1[0]), .out(far_4_5019_2[0]));    relay_conn far_4_5019_2_b(.in(far_4_5019_1[1]), .out(far_4_5019_2[1]));
    assign layer_4[939] = ~far_4_5019_2[1]; 
    assign layer_4[940] = layer_3[266] & layer_3[289]; 
    wire [1:0] far_4_5021_0;    relay_conn far_4_5021_0_a(.in(layer_3[321]), .out(far_4_5021_0[0]));    relay_conn far_4_5021_0_b(.in(layer_3[382]), .out(far_4_5021_0[1]));
    assign layer_4[941] = far_4_5021_0[1] & ~far_4_5021_0[0]; 
    assign layer_4[942] = layer_3[408] ^ layer_3[384]; 
    assign layer_4[943] = ~layer_3[10]; 
    assign layer_4[944] = layer_3[398] & ~layer_3[420]; 
    wire [1:0] far_4_5025_0;    relay_conn far_4_5025_0_a(.in(layer_3[345]), .out(far_4_5025_0[0]));    relay_conn far_4_5025_0_b(.in(layer_3[431]), .out(far_4_5025_0[1]));
    wire [1:0] far_4_5025_1;    relay_conn far_4_5025_1_a(.in(far_4_5025_0[0]), .out(far_4_5025_1[0]));    relay_conn far_4_5025_1_b(.in(far_4_5025_0[1]), .out(far_4_5025_1[1]));
    assign layer_4[945] = far_4_5025_1[0] & far_4_5025_1[1]; 
    wire [1:0] far_4_5026_0;    relay_conn far_4_5026_0_a(.in(layer_3[819]), .out(far_4_5026_0[0]));    relay_conn far_4_5026_0_b(.in(layer_3[866]), .out(far_4_5026_0[1]));
    assign layer_4[946] = far_4_5026_0[0] & far_4_5026_0[1]; 
    wire [1:0] far_4_5027_0;    relay_conn far_4_5027_0_a(.in(layer_3[719]), .out(far_4_5027_0[0]));    relay_conn far_4_5027_0_b(.in(layer_3[667]), .out(far_4_5027_0[1]));
    assign layer_4[947] = ~far_4_5027_0[0] | (far_4_5027_0[0] & far_4_5027_0[1]); 
    wire [1:0] far_4_5028_0;    relay_conn far_4_5028_0_a(.in(layer_3[885]), .out(far_4_5028_0[0]));    relay_conn far_4_5028_0_b(.in(layer_3[921]), .out(far_4_5028_0[1]));
    assign layer_4[948] = far_4_5028_0[1] & ~far_4_5028_0[0]; 
    assign layer_4[949] = ~(layer_3[625] & layer_3[598]); 
    wire [1:0] far_4_5030_0;    relay_conn far_4_5030_0_a(.in(layer_3[8]), .out(far_4_5030_0[0]));    relay_conn far_4_5030_0_b(.in(layer_3[69]), .out(far_4_5030_0[1]));
    assign layer_4[950] = far_4_5030_0[0] | far_4_5030_0[1]; 
    assign layer_4[951] = ~layer_3[408]; 
    wire [1:0] far_4_5032_0;    relay_conn far_4_5032_0_a(.in(layer_3[774]), .out(far_4_5032_0[0]));    relay_conn far_4_5032_0_b(.in(layer_3[857]), .out(far_4_5032_0[1]));
    wire [1:0] far_4_5032_1;    relay_conn far_4_5032_1_a(.in(far_4_5032_0[0]), .out(far_4_5032_1[0]));    relay_conn far_4_5032_1_b(.in(far_4_5032_0[1]), .out(far_4_5032_1[1]));
    assign layer_4[952] = ~(far_4_5032_1[0] | far_4_5032_1[1]); 
    assign layer_4[953] = layer_3[384] & layer_3[365]; 
    wire [1:0] far_4_5034_0;    relay_conn far_4_5034_0_a(.in(layer_3[748]), .out(far_4_5034_0[0]));    relay_conn far_4_5034_0_b(.in(layer_3[800]), .out(far_4_5034_0[1]));
    assign layer_4[954] = ~far_4_5034_0[1]; 
    wire [1:0] far_4_5035_0;    relay_conn far_4_5035_0_a(.in(layer_3[185]), .out(far_4_5035_0[0]));    relay_conn far_4_5035_0_b(.in(layer_3[279]), .out(far_4_5035_0[1]));
    wire [1:0] far_4_5035_1;    relay_conn far_4_5035_1_a(.in(far_4_5035_0[0]), .out(far_4_5035_1[0]));    relay_conn far_4_5035_1_b(.in(far_4_5035_0[1]), .out(far_4_5035_1[1]));
    assign layer_4[955] = far_4_5035_1[0]; 
    wire [1:0] far_4_5036_0;    relay_conn far_4_5036_0_a(.in(layer_3[335]), .out(far_4_5036_0[0]));    relay_conn far_4_5036_0_b(.in(layer_3[280]), .out(far_4_5036_0[1]));
    assign layer_4[956] = ~(far_4_5036_0[0] | far_4_5036_0[1]); 
    wire [1:0] far_4_5037_0;    relay_conn far_4_5037_0_a(.in(layer_3[105]), .out(far_4_5037_0[0]));    relay_conn far_4_5037_0_b(.in(layer_3[137]), .out(far_4_5037_0[1]));
    assign layer_4[957] = ~far_4_5037_0[0]; 
    wire [1:0] far_4_5038_0;    relay_conn far_4_5038_0_a(.in(layer_3[185]), .out(far_4_5038_0[0]));    relay_conn far_4_5038_0_b(.in(layer_3[274]), .out(far_4_5038_0[1]));
    wire [1:0] far_4_5038_1;    relay_conn far_4_5038_1_a(.in(far_4_5038_0[0]), .out(far_4_5038_1[0]));    relay_conn far_4_5038_1_b(.in(far_4_5038_0[1]), .out(far_4_5038_1[1]));
    assign layer_4[958] = far_4_5038_1[0] & far_4_5038_1[1]; 
    wire [1:0] far_4_5039_0;    relay_conn far_4_5039_0_a(.in(layer_3[274]), .out(far_4_5039_0[0]));    relay_conn far_4_5039_0_b(.in(layer_3[383]), .out(far_4_5039_0[1]));
    wire [1:0] far_4_5039_1;    relay_conn far_4_5039_1_a(.in(far_4_5039_0[0]), .out(far_4_5039_1[0]));    relay_conn far_4_5039_1_b(.in(far_4_5039_0[1]), .out(far_4_5039_1[1]));
    wire [1:0] far_4_5039_2;    relay_conn far_4_5039_2_a(.in(far_4_5039_1[0]), .out(far_4_5039_2[0]));    relay_conn far_4_5039_2_b(.in(far_4_5039_1[1]), .out(far_4_5039_2[1]));
    assign layer_4[959] = far_4_5039_2[0] & ~far_4_5039_2[1]; 
    wire [1:0] far_4_5040_0;    relay_conn far_4_5040_0_a(.in(layer_3[846]), .out(far_4_5040_0[0]));    relay_conn far_4_5040_0_b(.in(layer_3[788]), .out(far_4_5040_0[1]));
    assign layer_4[960] = ~far_4_5040_0[1] | (far_4_5040_0[0] & far_4_5040_0[1]); 
    wire [1:0] far_4_5041_0;    relay_conn far_4_5041_0_a(.in(layer_3[95]), .out(far_4_5041_0[0]));    relay_conn far_4_5041_0_b(.in(layer_3[178]), .out(far_4_5041_0[1]));
    wire [1:0] far_4_5041_1;    relay_conn far_4_5041_1_a(.in(far_4_5041_0[0]), .out(far_4_5041_1[0]));    relay_conn far_4_5041_1_b(.in(far_4_5041_0[1]), .out(far_4_5041_1[1]));
    assign layer_4[961] = ~far_4_5041_1[1] | (far_4_5041_1[0] & far_4_5041_1[1]); 
    assign layer_4[962] = ~layer_3[593]; 
    wire [1:0] far_4_5043_0;    relay_conn far_4_5043_0_a(.in(layer_3[532]), .out(far_4_5043_0[0]));    relay_conn far_4_5043_0_b(.in(layer_3[428]), .out(far_4_5043_0[1]));
    wire [1:0] far_4_5043_1;    relay_conn far_4_5043_1_a(.in(far_4_5043_0[0]), .out(far_4_5043_1[0]));    relay_conn far_4_5043_1_b(.in(far_4_5043_0[1]), .out(far_4_5043_1[1]));
    wire [1:0] far_4_5043_2;    relay_conn far_4_5043_2_a(.in(far_4_5043_1[0]), .out(far_4_5043_2[0]));    relay_conn far_4_5043_2_b(.in(far_4_5043_1[1]), .out(far_4_5043_2[1]));
    assign layer_4[963] = ~(far_4_5043_2[0] & far_4_5043_2[1]); 
    assign layer_4[964] = ~layer_3[874] | (layer_3[865] & layer_3[874]); 
    wire [1:0] far_4_5045_0;    relay_conn far_4_5045_0_a(.in(layer_3[898]), .out(far_4_5045_0[0]));    relay_conn far_4_5045_0_b(.in(layer_3[807]), .out(far_4_5045_0[1]));
    wire [1:0] far_4_5045_1;    relay_conn far_4_5045_1_a(.in(far_4_5045_0[0]), .out(far_4_5045_1[0]));    relay_conn far_4_5045_1_b(.in(far_4_5045_0[1]), .out(far_4_5045_1[1]));
    assign layer_4[965] = ~far_4_5045_1[0] | (far_4_5045_1[0] & far_4_5045_1[1]); 
    assign layer_4[966] = ~layer_3[781] | (layer_3[758] & layer_3[781]); 
    wire [1:0] far_4_5047_0;    relay_conn far_4_5047_0_a(.in(layer_3[710]), .out(far_4_5047_0[0]));    relay_conn far_4_5047_0_b(.in(layer_3[807]), .out(far_4_5047_0[1]));
    wire [1:0] far_4_5047_1;    relay_conn far_4_5047_1_a(.in(far_4_5047_0[0]), .out(far_4_5047_1[0]));    relay_conn far_4_5047_1_b(.in(far_4_5047_0[1]), .out(far_4_5047_1[1]));
    wire [1:0] far_4_5047_2;    relay_conn far_4_5047_2_a(.in(far_4_5047_1[0]), .out(far_4_5047_2[0]));    relay_conn far_4_5047_2_b(.in(far_4_5047_1[1]), .out(far_4_5047_2[1]));
    assign layer_4[967] = ~far_4_5047_2[1] | (far_4_5047_2[0] & far_4_5047_2[1]); 
    wire [1:0] far_4_5048_0;    relay_conn far_4_5048_0_a(.in(layer_3[394]), .out(far_4_5048_0[0]));    relay_conn far_4_5048_0_b(.in(layer_3[438]), .out(far_4_5048_0[1]));
    assign layer_4[968] = ~(far_4_5048_0[0] & far_4_5048_0[1]); 
    wire [1:0] far_4_5049_0;    relay_conn far_4_5049_0_a(.in(layer_3[527]), .out(far_4_5049_0[0]));    relay_conn far_4_5049_0_b(.in(layer_3[466]), .out(far_4_5049_0[1]));
    assign layer_4[969] = ~(far_4_5049_0[0] | far_4_5049_0[1]); 
    wire [1:0] far_4_5050_0;    relay_conn far_4_5050_0_a(.in(layer_3[376]), .out(far_4_5050_0[0]));    relay_conn far_4_5050_0_b(.in(layer_3[477]), .out(far_4_5050_0[1]));
    wire [1:0] far_4_5050_1;    relay_conn far_4_5050_1_a(.in(far_4_5050_0[0]), .out(far_4_5050_1[0]));    relay_conn far_4_5050_1_b(.in(far_4_5050_0[1]), .out(far_4_5050_1[1]));
    wire [1:0] far_4_5050_2;    relay_conn far_4_5050_2_a(.in(far_4_5050_1[0]), .out(far_4_5050_2[0]));    relay_conn far_4_5050_2_b(.in(far_4_5050_1[1]), .out(far_4_5050_2[1]));
    assign layer_4[970] = far_4_5050_2[1] & ~far_4_5050_2[0]; 
    assign layer_4[971] = ~layer_3[438]; 
    wire [1:0] far_4_5052_0;    relay_conn far_4_5052_0_a(.in(layer_3[644]), .out(far_4_5052_0[0]));    relay_conn far_4_5052_0_b(.in(layer_3[739]), .out(far_4_5052_0[1]));
    wire [1:0] far_4_5052_1;    relay_conn far_4_5052_1_a(.in(far_4_5052_0[0]), .out(far_4_5052_1[0]));    relay_conn far_4_5052_1_b(.in(far_4_5052_0[1]), .out(far_4_5052_1[1]));
    assign layer_4[972] = ~far_4_5052_1[0]; 
    wire [1:0] far_4_5053_0;    relay_conn far_4_5053_0_a(.in(layer_3[210]), .out(far_4_5053_0[0]));    relay_conn far_4_5053_0_b(.in(layer_3[321]), .out(far_4_5053_0[1]));
    wire [1:0] far_4_5053_1;    relay_conn far_4_5053_1_a(.in(far_4_5053_0[0]), .out(far_4_5053_1[0]));    relay_conn far_4_5053_1_b(.in(far_4_5053_0[1]), .out(far_4_5053_1[1]));
    wire [1:0] far_4_5053_2;    relay_conn far_4_5053_2_a(.in(far_4_5053_1[0]), .out(far_4_5053_2[0]));    relay_conn far_4_5053_2_b(.in(far_4_5053_1[1]), .out(far_4_5053_2[1]));
    assign layer_4[973] = ~far_4_5053_2[0]; 
    wire [1:0] far_4_5054_0;    relay_conn far_4_5054_0_a(.in(layer_3[380]), .out(far_4_5054_0[0]));    relay_conn far_4_5054_0_b(.in(layer_3[478]), .out(far_4_5054_0[1]));
    wire [1:0] far_4_5054_1;    relay_conn far_4_5054_1_a(.in(far_4_5054_0[0]), .out(far_4_5054_1[0]));    relay_conn far_4_5054_1_b(.in(far_4_5054_0[1]), .out(far_4_5054_1[1]));
    wire [1:0] far_4_5054_2;    relay_conn far_4_5054_2_a(.in(far_4_5054_1[0]), .out(far_4_5054_2[0]));    relay_conn far_4_5054_2_b(.in(far_4_5054_1[1]), .out(far_4_5054_2[1]));
    assign layer_4[974] = ~(far_4_5054_2[0] | far_4_5054_2[1]); 
    wire [1:0] far_4_5055_0;    relay_conn far_4_5055_0_a(.in(layer_3[431]), .out(far_4_5055_0[0]));    relay_conn far_4_5055_0_b(.in(layer_3[481]), .out(far_4_5055_0[1]));
    assign layer_4[975] = ~far_4_5055_0[1] | (far_4_5055_0[0] & far_4_5055_0[1]); 
    wire [1:0] far_4_5056_0;    relay_conn far_4_5056_0_a(.in(layer_3[398]), .out(far_4_5056_0[0]));    relay_conn far_4_5056_0_b(.in(layer_3[481]), .out(far_4_5056_0[1]));
    wire [1:0] far_4_5056_1;    relay_conn far_4_5056_1_a(.in(far_4_5056_0[0]), .out(far_4_5056_1[0]));    relay_conn far_4_5056_1_b(.in(far_4_5056_0[1]), .out(far_4_5056_1[1]));
    assign layer_4[976] = ~(far_4_5056_1[0] | far_4_5056_1[1]); 
    wire [1:0] far_4_5057_0;    relay_conn far_4_5057_0_a(.in(layer_3[916]), .out(far_4_5057_0[0]));    relay_conn far_4_5057_0_b(.in(layer_3[952]), .out(far_4_5057_0[1]));
    assign layer_4[977] = far_4_5057_0[1]; 
    wire [1:0] far_4_5058_0;    relay_conn far_4_5058_0_a(.in(layer_3[775]), .out(far_4_5058_0[0]));    relay_conn far_4_5058_0_b(.in(layer_3[837]), .out(far_4_5058_0[1]));
    assign layer_4[978] = ~far_4_5058_0[1]; 
    wire [1:0] far_4_5059_0;    relay_conn far_4_5059_0_a(.in(layer_3[544]), .out(far_4_5059_0[0]));    relay_conn far_4_5059_0_b(.in(layer_3[466]), .out(far_4_5059_0[1]));
    wire [1:0] far_4_5059_1;    relay_conn far_4_5059_1_a(.in(far_4_5059_0[0]), .out(far_4_5059_1[0]));    relay_conn far_4_5059_1_b(.in(far_4_5059_0[1]), .out(far_4_5059_1[1]));
    assign layer_4[979] = far_4_5059_1[0] & ~far_4_5059_1[1]; 
    wire [1:0] far_4_5060_0;    relay_conn far_4_5060_0_a(.in(layer_3[896]), .out(far_4_5060_0[0]));    relay_conn far_4_5060_0_b(.in(layer_3[807]), .out(far_4_5060_0[1]));
    wire [1:0] far_4_5060_1;    relay_conn far_4_5060_1_a(.in(far_4_5060_0[0]), .out(far_4_5060_1[0]));    relay_conn far_4_5060_1_b(.in(far_4_5060_0[1]), .out(far_4_5060_1[1]));
    assign layer_4[980] = ~far_4_5060_1[1]; 
    assign layer_4[981] = layer_3[342] & layer_3[314]; 
    wire [1:0] far_4_5062_0;    relay_conn far_4_5062_0_a(.in(layer_3[790]), .out(far_4_5062_0[0]));    relay_conn far_4_5062_0_b(.in(layer_3[880]), .out(far_4_5062_0[1]));
    wire [1:0] far_4_5062_1;    relay_conn far_4_5062_1_a(.in(far_4_5062_0[0]), .out(far_4_5062_1[0]));    relay_conn far_4_5062_1_b(.in(far_4_5062_0[1]), .out(far_4_5062_1[1]));
    assign layer_4[982] = far_4_5062_1[0]; 
    wire [1:0] far_4_5063_0;    relay_conn far_4_5063_0_a(.in(layer_3[615]), .out(far_4_5063_0[0]));    relay_conn far_4_5063_0_b(.in(layer_3[568]), .out(far_4_5063_0[1]));
    assign layer_4[983] = ~far_4_5063_0[0]; 
    wire [1:0] far_4_5064_0;    relay_conn far_4_5064_0_a(.in(layer_3[154]), .out(far_4_5064_0[0]));    relay_conn far_4_5064_0_b(.in(layer_3[278]), .out(far_4_5064_0[1]));
    wire [1:0] far_4_5064_1;    relay_conn far_4_5064_1_a(.in(far_4_5064_0[0]), .out(far_4_5064_1[0]));    relay_conn far_4_5064_1_b(.in(far_4_5064_0[1]), .out(far_4_5064_1[1]));
    wire [1:0] far_4_5064_2;    relay_conn far_4_5064_2_a(.in(far_4_5064_1[0]), .out(far_4_5064_2[0]));    relay_conn far_4_5064_2_b(.in(far_4_5064_1[1]), .out(far_4_5064_2[1]));
    assign layer_4[984] = far_4_5064_2[0] | far_4_5064_2[1]; 
    wire [1:0] far_4_5065_0;    relay_conn far_4_5065_0_a(.in(layer_3[552]), .out(far_4_5065_0[0]));    relay_conn far_4_5065_0_b(.in(layer_3[480]), .out(far_4_5065_0[1]));
    wire [1:0] far_4_5065_1;    relay_conn far_4_5065_1_a(.in(far_4_5065_0[0]), .out(far_4_5065_1[0]));    relay_conn far_4_5065_1_b(.in(far_4_5065_0[1]), .out(far_4_5065_1[1]));
    assign layer_4[985] = ~far_4_5065_1[1] | (far_4_5065_1[0] & far_4_5065_1[1]); 
    wire [1:0] far_4_5066_0;    relay_conn far_4_5066_0_a(.in(layer_3[391]), .out(far_4_5066_0[0]));    relay_conn far_4_5066_0_b(.in(layer_3[477]), .out(far_4_5066_0[1]));
    wire [1:0] far_4_5066_1;    relay_conn far_4_5066_1_a(.in(far_4_5066_0[0]), .out(far_4_5066_1[0]));    relay_conn far_4_5066_1_b(.in(far_4_5066_0[1]), .out(far_4_5066_1[1]));
    assign layer_4[986] = far_4_5066_1[1] & ~far_4_5066_1[0]; 
    wire [1:0] far_4_5067_0;    relay_conn far_4_5067_0_a(.in(layer_3[844]), .out(far_4_5067_0[0]));    relay_conn far_4_5067_0_b(.in(layer_3[807]), .out(far_4_5067_0[1]));
    assign layer_4[987] = ~far_4_5067_0[0]; 
    wire [1:0] far_4_5068_0;    relay_conn far_4_5068_0_a(.in(layer_3[718]), .out(far_4_5068_0[0]));    relay_conn far_4_5068_0_b(.in(layer_3[807]), .out(far_4_5068_0[1]));
    wire [1:0] far_4_5068_1;    relay_conn far_4_5068_1_a(.in(far_4_5068_0[0]), .out(far_4_5068_1[0]));    relay_conn far_4_5068_1_b(.in(far_4_5068_0[1]), .out(far_4_5068_1[1]));
    assign layer_4[988] = ~(far_4_5068_1[0] & far_4_5068_1[1]); 
    assign layer_4[989] = ~layer_3[625]; 
    wire [1:0] far_4_5070_0;    relay_conn far_4_5070_0_a(.in(layer_3[809]), .out(far_4_5070_0[0]));    relay_conn far_4_5070_0_b(.in(layer_3[868]), .out(far_4_5070_0[1]));
    assign layer_4[990] = far_4_5070_0[0] | far_4_5070_0[1]; 
    wire [1:0] far_4_5071_0;    relay_conn far_4_5071_0_a(.in(layer_3[576]), .out(far_4_5071_0[0]));    relay_conn far_4_5071_0_b(.in(layer_3[475]), .out(far_4_5071_0[1]));
    wire [1:0] far_4_5071_1;    relay_conn far_4_5071_1_a(.in(far_4_5071_0[0]), .out(far_4_5071_1[0]));    relay_conn far_4_5071_1_b(.in(far_4_5071_0[1]), .out(far_4_5071_1[1]));
    wire [1:0] far_4_5071_2;    relay_conn far_4_5071_2_a(.in(far_4_5071_1[0]), .out(far_4_5071_2[0]));    relay_conn far_4_5071_2_b(.in(far_4_5071_1[1]), .out(far_4_5071_2[1]));
    assign layer_4[991] = far_4_5071_2[0] & far_4_5071_2[1]; 
    assign layer_4[992] = layer_3[950]; 
    wire [1:0] far_4_5073_0;    relay_conn far_4_5073_0_a(.in(layer_3[504]), .out(far_4_5073_0[0]));    relay_conn far_4_5073_0_b(.in(layer_3[576]), .out(far_4_5073_0[1]));
    wire [1:0] far_4_5073_1;    relay_conn far_4_5073_1_a(.in(far_4_5073_0[0]), .out(far_4_5073_1[0]));    relay_conn far_4_5073_1_b(.in(far_4_5073_0[1]), .out(far_4_5073_1[1]));
    assign layer_4[993] = ~(far_4_5073_1[0] ^ far_4_5073_1[1]); 
    wire [1:0] far_4_5074_0;    relay_conn far_4_5074_0_a(.in(layer_3[857]), .out(far_4_5074_0[0]));    relay_conn far_4_5074_0_b(.in(layer_3[916]), .out(far_4_5074_0[1]));
    assign layer_4[994] = far_4_5074_0[0] & ~far_4_5074_0[1]; 
    wire [1:0] far_4_5075_0;    relay_conn far_4_5075_0_a(.in(layer_3[478]), .out(far_4_5075_0[0]));    relay_conn far_4_5075_0_b(.in(layer_3[428]), .out(far_4_5075_0[1]));
    assign layer_4[995] = ~far_4_5075_0[1]; 
    assign layer_4[996] = ~layer_3[302]; 
    assign layer_4[997] = ~layer_3[317] | (layer_3[329] & layer_3[317]); 
    wire [1:0] far_4_5078_0;    relay_conn far_4_5078_0_a(.in(layer_3[664]), .out(far_4_5078_0[0]));    relay_conn far_4_5078_0_b(.in(layer_3[570]), .out(far_4_5078_0[1]));
    wire [1:0] far_4_5078_1;    relay_conn far_4_5078_1_a(.in(far_4_5078_0[0]), .out(far_4_5078_1[0]));    relay_conn far_4_5078_1_b(.in(far_4_5078_0[1]), .out(far_4_5078_1[1]));
    assign layer_4[998] = ~far_4_5078_1[0]; 
    wire [1:0] far_4_5079_0;    relay_conn far_4_5079_0_a(.in(layer_3[592]), .out(far_4_5079_0[0]));    relay_conn far_4_5079_0_b(.in(layer_3[664]), .out(far_4_5079_0[1]));
    wire [1:0] far_4_5079_1;    relay_conn far_4_5079_1_a(.in(far_4_5079_0[0]), .out(far_4_5079_1[0]));    relay_conn far_4_5079_1_b(.in(far_4_5079_0[1]), .out(far_4_5079_1[1]));
    assign layer_4[999] = ~far_4_5079_1[1]; 
    wire [1:0] far_4_5080_0;    relay_conn far_4_5080_0_a(.in(layer_3[274]), .out(far_4_5080_0[0]));    relay_conn far_4_5080_0_b(.in(layer_3[334]), .out(far_4_5080_0[1]));
    assign layer_4[1000] = ~far_4_5080_0[1]; 
    wire [1:0] far_4_5081_0;    relay_conn far_4_5081_0_a(.in(layer_3[373]), .out(far_4_5081_0[0]));    relay_conn far_4_5081_0_b(.in(layer_3[475]), .out(far_4_5081_0[1]));
    wire [1:0] far_4_5081_1;    relay_conn far_4_5081_1_a(.in(far_4_5081_0[0]), .out(far_4_5081_1[0]));    relay_conn far_4_5081_1_b(.in(far_4_5081_0[1]), .out(far_4_5081_1[1]));
    wire [1:0] far_4_5081_2;    relay_conn far_4_5081_2_a(.in(far_4_5081_1[0]), .out(far_4_5081_2[0]));    relay_conn far_4_5081_2_b(.in(far_4_5081_1[1]), .out(far_4_5081_2[1]));
    assign layer_4[1001] = ~far_4_5081_2[1]; 
    wire [1:0] far_4_5082_0;    relay_conn far_4_5082_0_a(.in(layer_3[35]), .out(far_4_5082_0[0]));    relay_conn far_4_5082_0_b(.in(layer_3[104]), .out(far_4_5082_0[1]));
    wire [1:0] far_4_5082_1;    relay_conn far_4_5082_1_a(.in(far_4_5082_0[0]), .out(far_4_5082_1[0]));    relay_conn far_4_5082_1_b(.in(far_4_5082_0[1]), .out(far_4_5082_1[1]));
    assign layer_4[1002] = far_4_5082_1[0] | far_4_5082_1[1]; 
    wire [1:0] far_4_5083_0;    relay_conn far_4_5083_0_a(.in(layer_3[402]), .out(far_4_5083_0[0]));    relay_conn far_4_5083_0_b(.in(layer_3[318]), .out(far_4_5083_0[1]));
    wire [1:0] far_4_5083_1;    relay_conn far_4_5083_1_a(.in(far_4_5083_0[0]), .out(far_4_5083_1[0]));    relay_conn far_4_5083_1_b(.in(far_4_5083_0[1]), .out(far_4_5083_1[1]));
    assign layer_4[1003] = ~(far_4_5083_1[0] | far_4_5083_1[1]); 
    wire [1:0] far_4_5084_0;    relay_conn far_4_5084_0_a(.in(layer_3[859]), .out(far_4_5084_0[0]));    relay_conn far_4_5084_0_b(.in(layer_3[962]), .out(far_4_5084_0[1]));
    wire [1:0] far_4_5084_1;    relay_conn far_4_5084_1_a(.in(far_4_5084_0[0]), .out(far_4_5084_1[0]));    relay_conn far_4_5084_1_b(.in(far_4_5084_0[1]), .out(far_4_5084_1[1]));
    wire [1:0] far_4_5084_2;    relay_conn far_4_5084_2_a(.in(far_4_5084_1[0]), .out(far_4_5084_2[0]));    relay_conn far_4_5084_2_b(.in(far_4_5084_1[1]), .out(far_4_5084_2[1]));
    assign layer_4[1004] = ~far_4_5084_2[1]; 
    wire [1:0] far_4_5085_0;    relay_conn far_4_5085_0_a(.in(layer_3[256]), .out(far_4_5085_0[0]));    relay_conn far_4_5085_0_b(.in(layer_3[200]), .out(far_4_5085_0[1]));
    assign layer_4[1005] = ~(far_4_5085_0[0] | far_4_5085_0[1]); 
    wire [1:0] far_4_5086_0;    relay_conn far_4_5086_0_a(.in(layer_3[0]), .out(far_4_5086_0[0]));    relay_conn far_4_5086_0_b(.in(layer_3[110]), .out(far_4_5086_0[1]));
    wire [1:0] far_4_5086_1;    relay_conn far_4_5086_1_a(.in(far_4_5086_0[0]), .out(far_4_5086_1[0]));    relay_conn far_4_5086_1_b(.in(far_4_5086_0[1]), .out(far_4_5086_1[1]));
    wire [1:0] far_4_5086_2;    relay_conn far_4_5086_2_a(.in(far_4_5086_1[0]), .out(far_4_5086_2[0]));    relay_conn far_4_5086_2_b(.in(far_4_5086_1[1]), .out(far_4_5086_2[1]));
    assign layer_4[1006] = ~far_4_5086_2[1]; 
    wire [1:0] far_4_5087_0;    relay_conn far_4_5087_0_a(.in(layer_3[331]), .out(far_4_5087_0[0]));    relay_conn far_4_5087_0_b(.in(layer_3[398]), .out(far_4_5087_0[1]));
    wire [1:0] far_4_5087_1;    relay_conn far_4_5087_1_a(.in(far_4_5087_0[0]), .out(far_4_5087_1[0]));    relay_conn far_4_5087_1_b(.in(far_4_5087_0[1]), .out(far_4_5087_1[1]));
    assign layer_4[1007] = far_4_5087_1[0] ^ far_4_5087_1[1]; 
    assign layer_4[1008] = layer_3[667] | layer_3[674]; 
    wire [1:0] far_4_5089_0;    relay_conn far_4_5089_0_a(.in(layer_3[323]), .out(far_4_5089_0[0]));    relay_conn far_4_5089_0_b(.in(layer_3[271]), .out(far_4_5089_0[1]));
    assign layer_4[1009] = ~(far_4_5089_0[0] | far_4_5089_0[1]); 
    wire [1:0] far_4_5090_0;    relay_conn far_4_5090_0_a(.in(layer_3[408]), .out(far_4_5090_0[0]));    relay_conn far_4_5090_0_b(.in(layer_3[504]), .out(far_4_5090_0[1]));
    wire [1:0] far_4_5090_1;    relay_conn far_4_5090_1_a(.in(far_4_5090_0[0]), .out(far_4_5090_1[0]));    relay_conn far_4_5090_1_b(.in(far_4_5090_0[1]), .out(far_4_5090_1[1]));
    wire [1:0] far_4_5090_2;    relay_conn far_4_5090_2_a(.in(far_4_5090_1[0]), .out(far_4_5090_2[0]));    relay_conn far_4_5090_2_b(.in(far_4_5090_1[1]), .out(far_4_5090_2[1]));
    assign layer_4[1010] = ~far_4_5090_2[1]; 
    wire [1:0] far_4_5091_0;    relay_conn far_4_5091_0_a(.in(layer_3[466]), .out(far_4_5091_0[0]));    relay_conn far_4_5091_0_b(.in(layer_3[498]), .out(far_4_5091_0[1]));
    assign layer_4[1011] = far_4_5091_0[1] & ~far_4_5091_0[0]; 
    assign layer_4[1012] = ~layer_3[454]; 
    wire [1:0] far_4_5093_0;    relay_conn far_4_5093_0_a(.in(layer_3[362]), .out(far_4_5093_0[0]));    relay_conn far_4_5093_0_b(.in(layer_3[424]), .out(far_4_5093_0[1]));
    assign layer_4[1013] = far_4_5093_0[0] & ~far_4_5093_0[1]; 
    wire [1:0] far_4_5094_0;    relay_conn far_4_5094_0_a(.in(layer_3[353]), .out(far_4_5094_0[0]));    relay_conn far_4_5094_0_b(.in(layer_3[393]), .out(far_4_5094_0[1]));
    assign layer_4[1014] = far_4_5094_0[1] & ~far_4_5094_0[0]; 
    wire [1:0] far_4_5095_0;    relay_conn far_4_5095_0_a(.in(layer_3[949]), .out(far_4_5095_0[0]));    relay_conn far_4_5095_0_b(.in(layer_3[843]), .out(far_4_5095_0[1]));
    wire [1:0] far_4_5095_1;    relay_conn far_4_5095_1_a(.in(far_4_5095_0[0]), .out(far_4_5095_1[0]));    relay_conn far_4_5095_1_b(.in(far_4_5095_0[1]), .out(far_4_5095_1[1]));
    wire [1:0] far_4_5095_2;    relay_conn far_4_5095_2_a(.in(far_4_5095_1[0]), .out(far_4_5095_2[0]));    relay_conn far_4_5095_2_b(.in(far_4_5095_1[1]), .out(far_4_5095_2[1]));
    assign layer_4[1015] = ~(far_4_5095_2[0] | far_4_5095_2[1]); 
    wire [1:0] far_4_5096_0;    relay_conn far_4_5096_0_a(.in(layer_3[576]), .out(far_4_5096_0[0]));    relay_conn far_4_5096_0_b(.in(layer_3[542]), .out(far_4_5096_0[1]));
    assign layer_4[1016] = far_4_5096_0[0]; 
    wire [1:0] far_4_5097_0;    relay_conn far_4_5097_0_a(.in(layer_3[143]), .out(far_4_5097_0[0]));    relay_conn far_4_5097_0_b(.in(layer_3[200]), .out(far_4_5097_0[1]));
    assign layer_4[1017] = far_4_5097_0[0] | far_4_5097_0[1]; 
    wire [1:0] far_4_5098_0;    relay_conn far_4_5098_0_a(.in(layer_3[653]), .out(far_4_5098_0[0]));    relay_conn far_4_5098_0_b(.in(layer_3[568]), .out(far_4_5098_0[1]));
    wire [1:0] far_4_5098_1;    relay_conn far_4_5098_1_a(.in(far_4_5098_0[0]), .out(far_4_5098_1[0]));    relay_conn far_4_5098_1_b(.in(far_4_5098_0[1]), .out(far_4_5098_1[1]));
    assign layer_4[1018] = ~far_4_5098_1[1]; 
    wire [1:0] far_4_5099_0;    relay_conn far_4_5099_0_a(.in(layer_3[831]), .out(far_4_5099_0[0]));    relay_conn far_4_5099_0_b(.in(layer_3[958]), .out(far_4_5099_0[1]));
    wire [1:0] far_4_5099_1;    relay_conn far_4_5099_1_a(.in(far_4_5099_0[0]), .out(far_4_5099_1[0]));    relay_conn far_4_5099_1_b(.in(far_4_5099_0[1]), .out(far_4_5099_1[1]));
    wire [1:0] far_4_5099_2;    relay_conn far_4_5099_2_a(.in(far_4_5099_1[0]), .out(far_4_5099_2[0]));    relay_conn far_4_5099_2_b(.in(far_4_5099_1[1]), .out(far_4_5099_2[1]));
    assign layer_4[1019] = ~(far_4_5099_2[0] | far_4_5099_2[1]); 
    // Layer 5 ============================================================
    wire [1:0] far_5_5100_0;    relay_conn far_5_5100_0_a(.in(layer_4[392]), .out(far_5_5100_0[0]));    relay_conn far_5_5100_0_b(.in(layer_4[451]), .out(far_5_5100_0[1]));
    assign layer_5[0] = far_5_5100_0[1] & ~far_5_5100_0[0]; 
    wire [1:0] far_5_5101_0;    relay_conn far_5_5101_0_a(.in(layer_4[284]), .out(far_5_5101_0[0]));    relay_conn far_5_5101_0_b(.in(layer_4[324]), .out(far_5_5101_0[1]));
    assign layer_5[1] = ~far_5_5101_0[0] | (far_5_5101_0[0] & far_5_5101_0[1]); 
    wire [1:0] far_5_5102_0;    relay_conn far_5_5102_0_a(.in(layer_4[620]), .out(far_5_5102_0[0]));    relay_conn far_5_5102_0_b(.in(layer_4[692]), .out(far_5_5102_0[1]));
    wire [1:0] far_5_5102_1;    relay_conn far_5_5102_1_a(.in(far_5_5102_0[0]), .out(far_5_5102_1[0]));    relay_conn far_5_5102_1_b(.in(far_5_5102_0[1]), .out(far_5_5102_1[1]));
    assign layer_5[2] = ~far_5_5102_1[0]; 
    wire [1:0] far_5_5103_0;    relay_conn far_5_5103_0_a(.in(layer_4[212]), .out(far_5_5103_0[0]));    relay_conn far_5_5103_0_b(.in(layer_4[168]), .out(far_5_5103_0[1]));
    assign layer_5[3] = far_5_5103_0[1]; 
    wire [1:0] far_5_5104_0;    relay_conn far_5_5104_0_a(.in(layer_4[127]), .out(far_5_5104_0[0]));    relay_conn far_5_5104_0_b(.in(layer_4[8]), .out(far_5_5104_0[1]));
    wire [1:0] far_5_5104_1;    relay_conn far_5_5104_1_a(.in(far_5_5104_0[0]), .out(far_5_5104_1[0]));    relay_conn far_5_5104_1_b(.in(far_5_5104_0[1]), .out(far_5_5104_1[1]));
    wire [1:0] far_5_5104_2;    relay_conn far_5_5104_2_a(.in(far_5_5104_1[0]), .out(far_5_5104_2[0]));    relay_conn far_5_5104_2_b(.in(far_5_5104_1[1]), .out(far_5_5104_2[1]));
    assign layer_5[4] = ~(far_5_5104_2[0] | far_5_5104_2[1]); 
    wire [1:0] far_5_5105_0;    relay_conn far_5_5105_0_a(.in(layer_4[898]), .out(far_5_5105_0[0]));    relay_conn far_5_5105_0_b(.in(layer_4[932]), .out(far_5_5105_0[1]));
    assign layer_5[5] = far_5_5105_0[0] & ~far_5_5105_0[1]; 
    wire [1:0] far_5_5106_0;    relay_conn far_5_5106_0_a(.in(layer_4[650]), .out(far_5_5106_0[0]));    relay_conn far_5_5106_0_b(.in(layer_4[542]), .out(far_5_5106_0[1]));
    wire [1:0] far_5_5106_1;    relay_conn far_5_5106_1_a(.in(far_5_5106_0[0]), .out(far_5_5106_1[0]));    relay_conn far_5_5106_1_b(.in(far_5_5106_0[1]), .out(far_5_5106_1[1]));
    wire [1:0] far_5_5106_2;    relay_conn far_5_5106_2_a(.in(far_5_5106_1[0]), .out(far_5_5106_2[0]));    relay_conn far_5_5106_2_b(.in(far_5_5106_1[1]), .out(far_5_5106_2[1]));
    assign layer_5[6] = ~far_5_5106_2[1]; 
    assign layer_5[7] = ~layer_4[995] | (layer_4[995] & layer_4[977]); 
    wire [1:0] far_5_5108_0;    relay_conn far_5_5108_0_a(.in(layer_4[521]), .out(far_5_5108_0[0]));    relay_conn far_5_5108_0_b(.in(layer_4[585]), .out(far_5_5108_0[1]));
    wire [1:0] far_5_5108_1;    relay_conn far_5_5108_1_a(.in(far_5_5108_0[0]), .out(far_5_5108_1[0]));    relay_conn far_5_5108_1_b(.in(far_5_5108_0[1]), .out(far_5_5108_1[1]));
    assign layer_5[8] = ~(far_5_5108_1[0] & far_5_5108_1[1]); 
    wire [1:0] far_5_5109_0;    relay_conn far_5_5109_0_a(.in(layer_4[736]), .out(far_5_5109_0[0]));    relay_conn far_5_5109_0_b(.in(layer_4[675]), .out(far_5_5109_0[1]));
    assign layer_5[9] = ~(far_5_5109_0[0] ^ far_5_5109_0[1]); 
    wire [1:0] far_5_5110_0;    relay_conn far_5_5110_0_a(.in(layer_4[602]), .out(far_5_5110_0[0]));    relay_conn far_5_5110_0_b(.in(layer_4[728]), .out(far_5_5110_0[1]));
    wire [1:0] far_5_5110_1;    relay_conn far_5_5110_1_a(.in(far_5_5110_0[0]), .out(far_5_5110_1[0]));    relay_conn far_5_5110_1_b(.in(far_5_5110_0[1]), .out(far_5_5110_1[1]));
    wire [1:0] far_5_5110_2;    relay_conn far_5_5110_2_a(.in(far_5_5110_1[0]), .out(far_5_5110_2[0]));    relay_conn far_5_5110_2_b(.in(far_5_5110_1[1]), .out(far_5_5110_2[1]));
    assign layer_5[10] = far_5_5110_2[0] & far_5_5110_2[1]; 
    wire [1:0] far_5_5111_0;    relay_conn far_5_5111_0_a(.in(layer_4[632]), .out(far_5_5111_0[0]));    relay_conn far_5_5111_0_b(.in(layer_4[742]), .out(far_5_5111_0[1]));
    wire [1:0] far_5_5111_1;    relay_conn far_5_5111_1_a(.in(far_5_5111_0[0]), .out(far_5_5111_1[0]));    relay_conn far_5_5111_1_b(.in(far_5_5111_0[1]), .out(far_5_5111_1[1]));
    wire [1:0] far_5_5111_2;    relay_conn far_5_5111_2_a(.in(far_5_5111_1[0]), .out(far_5_5111_2[0]));    relay_conn far_5_5111_2_b(.in(far_5_5111_1[1]), .out(far_5_5111_2[1]));
    assign layer_5[11] = far_5_5111_2[1]; 
    wire [1:0] far_5_5112_0;    relay_conn far_5_5112_0_a(.in(layer_4[654]), .out(far_5_5112_0[0]));    relay_conn far_5_5112_0_b(.in(layer_4[597]), .out(far_5_5112_0[1]));
    assign layer_5[12] = far_5_5112_0[0] & far_5_5112_0[1]; 
    assign layer_5[13] = ~layer_4[499] | (layer_4[499] & layer_4[475]); 
    wire [1:0] far_5_5114_0;    relay_conn far_5_5114_0_a(.in(layer_4[845]), .out(far_5_5114_0[0]));    relay_conn far_5_5114_0_b(.in(layer_4[930]), .out(far_5_5114_0[1]));
    wire [1:0] far_5_5114_1;    relay_conn far_5_5114_1_a(.in(far_5_5114_0[0]), .out(far_5_5114_1[0]));    relay_conn far_5_5114_1_b(.in(far_5_5114_0[1]), .out(far_5_5114_1[1]));
    assign layer_5[14] = ~(far_5_5114_1[0] | far_5_5114_1[1]); 
    assign layer_5[15] = ~layer_4[266] | (layer_4[266] & layer_4[286]); 
    assign layer_5[16] = layer_4[759] ^ layer_4[778]; 
    wire [1:0] far_5_5117_0;    relay_conn far_5_5117_0_a(.in(layer_4[697]), .out(far_5_5117_0[0]));    relay_conn far_5_5117_0_b(.in(layer_4[812]), .out(far_5_5117_0[1]));
    wire [1:0] far_5_5117_1;    relay_conn far_5_5117_1_a(.in(far_5_5117_0[0]), .out(far_5_5117_1[0]));    relay_conn far_5_5117_1_b(.in(far_5_5117_0[1]), .out(far_5_5117_1[1]));
    wire [1:0] far_5_5117_2;    relay_conn far_5_5117_2_a(.in(far_5_5117_1[0]), .out(far_5_5117_2[0]));    relay_conn far_5_5117_2_b(.in(far_5_5117_1[1]), .out(far_5_5117_2[1]));
    assign layer_5[17] = ~far_5_5117_2[1]; 
    wire [1:0] far_5_5118_0;    relay_conn far_5_5118_0_a(.in(layer_4[94]), .out(far_5_5118_0[0]));    relay_conn far_5_5118_0_b(.in(layer_4[170]), .out(far_5_5118_0[1]));
    wire [1:0] far_5_5118_1;    relay_conn far_5_5118_1_a(.in(far_5_5118_0[0]), .out(far_5_5118_1[0]));    relay_conn far_5_5118_1_b(.in(far_5_5118_0[1]), .out(far_5_5118_1[1]));
    assign layer_5[18] = ~(far_5_5118_1[0] & far_5_5118_1[1]); 
    wire [1:0] far_5_5119_0;    relay_conn far_5_5119_0_a(.in(layer_4[65]), .out(far_5_5119_0[0]));    relay_conn far_5_5119_0_b(.in(layer_4[175]), .out(far_5_5119_0[1]));
    wire [1:0] far_5_5119_1;    relay_conn far_5_5119_1_a(.in(far_5_5119_0[0]), .out(far_5_5119_1[0]));    relay_conn far_5_5119_1_b(.in(far_5_5119_0[1]), .out(far_5_5119_1[1]));
    wire [1:0] far_5_5119_2;    relay_conn far_5_5119_2_a(.in(far_5_5119_1[0]), .out(far_5_5119_2[0]));    relay_conn far_5_5119_2_b(.in(far_5_5119_1[1]), .out(far_5_5119_2[1]));
    assign layer_5[19] = ~(far_5_5119_2[0] ^ far_5_5119_2[1]); 
    wire [1:0] far_5_5120_0;    relay_conn far_5_5120_0_a(.in(layer_4[516]), .out(far_5_5120_0[0]));    relay_conn far_5_5120_0_b(.in(layer_4[616]), .out(far_5_5120_0[1]));
    wire [1:0] far_5_5120_1;    relay_conn far_5_5120_1_a(.in(far_5_5120_0[0]), .out(far_5_5120_1[0]));    relay_conn far_5_5120_1_b(.in(far_5_5120_0[1]), .out(far_5_5120_1[1]));
    wire [1:0] far_5_5120_2;    relay_conn far_5_5120_2_a(.in(far_5_5120_1[0]), .out(far_5_5120_2[0]));    relay_conn far_5_5120_2_b(.in(far_5_5120_1[1]), .out(far_5_5120_2[1]));
    assign layer_5[20] = far_5_5120_2[0] ^ far_5_5120_2[1]; 
    wire [1:0] far_5_5121_0;    relay_conn far_5_5121_0_a(.in(layer_4[325]), .out(far_5_5121_0[0]));    relay_conn far_5_5121_0_b(.in(layer_4[419]), .out(far_5_5121_0[1]));
    wire [1:0] far_5_5121_1;    relay_conn far_5_5121_1_a(.in(far_5_5121_0[0]), .out(far_5_5121_1[0]));    relay_conn far_5_5121_1_b(.in(far_5_5121_0[1]), .out(far_5_5121_1[1]));
    assign layer_5[21] = far_5_5121_1[0]; 
    wire [1:0] far_5_5122_0;    relay_conn far_5_5122_0_a(.in(layer_4[478]), .out(far_5_5122_0[0]));    relay_conn far_5_5122_0_b(.in(layer_4[516]), .out(far_5_5122_0[1]));
    assign layer_5[22] = ~far_5_5122_0[1] | (far_5_5122_0[0] & far_5_5122_0[1]); 
    assign layer_5[23] = ~layer_4[983] | (layer_4[974] & layer_4[983]); 
    wire [1:0] far_5_5124_0;    relay_conn far_5_5124_0_a(.in(layer_4[546]), .out(far_5_5124_0[0]));    relay_conn far_5_5124_0_b(.in(layer_4[633]), .out(far_5_5124_0[1]));
    wire [1:0] far_5_5124_1;    relay_conn far_5_5124_1_a(.in(far_5_5124_0[0]), .out(far_5_5124_1[0]));    relay_conn far_5_5124_1_b(.in(far_5_5124_0[1]), .out(far_5_5124_1[1]));
    assign layer_5[24] = far_5_5124_1[0] | far_5_5124_1[1]; 
    wire [1:0] far_5_5125_0;    relay_conn far_5_5125_0_a(.in(layer_4[357]), .out(far_5_5125_0[0]));    relay_conn far_5_5125_0_b(.in(layer_4[261]), .out(far_5_5125_0[1]));
    wire [1:0] far_5_5125_1;    relay_conn far_5_5125_1_a(.in(far_5_5125_0[0]), .out(far_5_5125_1[0]));    relay_conn far_5_5125_1_b(.in(far_5_5125_0[1]), .out(far_5_5125_1[1]));
    wire [1:0] far_5_5125_2;    relay_conn far_5_5125_2_a(.in(far_5_5125_1[0]), .out(far_5_5125_2[0]));    relay_conn far_5_5125_2_b(.in(far_5_5125_1[1]), .out(far_5_5125_2[1]));
    assign layer_5[25] = ~far_5_5125_2[1] | (far_5_5125_2[0] & far_5_5125_2[1]); 
    assign layer_5[26] = layer_4[656]; 
    wire [1:0] far_5_5127_0;    relay_conn far_5_5127_0_a(.in(layer_4[559]), .out(far_5_5127_0[0]));    relay_conn far_5_5127_0_b(.in(layer_4[665]), .out(far_5_5127_0[1]));
    wire [1:0] far_5_5127_1;    relay_conn far_5_5127_1_a(.in(far_5_5127_0[0]), .out(far_5_5127_1[0]));    relay_conn far_5_5127_1_b(.in(far_5_5127_0[1]), .out(far_5_5127_1[1]));
    wire [1:0] far_5_5127_2;    relay_conn far_5_5127_2_a(.in(far_5_5127_1[0]), .out(far_5_5127_2[0]));    relay_conn far_5_5127_2_b(.in(far_5_5127_1[1]), .out(far_5_5127_2[1]));
    assign layer_5[27] = ~far_5_5127_2[0] | (far_5_5127_2[0] & far_5_5127_2[1]); 
    wire [1:0] far_5_5128_0;    relay_conn far_5_5128_0_a(.in(layer_4[650]), .out(far_5_5128_0[0]));    relay_conn far_5_5128_0_b(.in(layer_4[752]), .out(far_5_5128_0[1]));
    wire [1:0] far_5_5128_1;    relay_conn far_5_5128_1_a(.in(far_5_5128_0[0]), .out(far_5_5128_1[0]));    relay_conn far_5_5128_1_b(.in(far_5_5128_0[1]), .out(far_5_5128_1[1]));
    wire [1:0] far_5_5128_2;    relay_conn far_5_5128_2_a(.in(far_5_5128_1[0]), .out(far_5_5128_2[0]));    relay_conn far_5_5128_2_b(.in(far_5_5128_1[1]), .out(far_5_5128_2[1]));
    assign layer_5[28] = ~(far_5_5128_2[0] & far_5_5128_2[1]); 
    wire [1:0] far_5_5129_0;    relay_conn far_5_5129_0_a(.in(layer_4[397]), .out(far_5_5129_0[0]));    relay_conn far_5_5129_0_b(.in(layer_4[497]), .out(far_5_5129_0[1]));
    wire [1:0] far_5_5129_1;    relay_conn far_5_5129_1_a(.in(far_5_5129_0[0]), .out(far_5_5129_1[0]));    relay_conn far_5_5129_1_b(.in(far_5_5129_0[1]), .out(far_5_5129_1[1]));
    wire [1:0] far_5_5129_2;    relay_conn far_5_5129_2_a(.in(far_5_5129_1[0]), .out(far_5_5129_2[0]));    relay_conn far_5_5129_2_b(.in(far_5_5129_1[1]), .out(far_5_5129_2[1]));
    assign layer_5[29] = far_5_5129_2[0] & ~far_5_5129_2[1]; 
    assign layer_5[30] = layer_4[528] & ~layer_4[525]; 
    wire [1:0] far_5_5131_0;    relay_conn far_5_5131_0_a(.in(layer_4[455]), .out(far_5_5131_0[0]));    relay_conn far_5_5131_0_b(.in(layer_4[331]), .out(far_5_5131_0[1]));
    wire [1:0] far_5_5131_1;    relay_conn far_5_5131_1_a(.in(far_5_5131_0[0]), .out(far_5_5131_1[0]));    relay_conn far_5_5131_1_b(.in(far_5_5131_0[1]), .out(far_5_5131_1[1]));
    wire [1:0] far_5_5131_2;    relay_conn far_5_5131_2_a(.in(far_5_5131_1[0]), .out(far_5_5131_2[0]));    relay_conn far_5_5131_2_b(.in(far_5_5131_1[1]), .out(far_5_5131_2[1]));
    assign layer_5[31] = far_5_5131_2[1]; 
    wire [1:0] far_5_5132_0;    relay_conn far_5_5132_0_a(.in(layer_4[363]), .out(far_5_5132_0[0]));    relay_conn far_5_5132_0_b(.in(layer_4[422]), .out(far_5_5132_0[1]));
    assign layer_5[32] = far_5_5132_0[0] ^ far_5_5132_0[1]; 
    wire [1:0] far_5_5133_0;    relay_conn far_5_5133_0_a(.in(layer_4[571]), .out(far_5_5133_0[0]));    relay_conn far_5_5133_0_b(.in(layer_4[656]), .out(far_5_5133_0[1]));
    wire [1:0] far_5_5133_1;    relay_conn far_5_5133_1_a(.in(far_5_5133_0[0]), .out(far_5_5133_1[0]));    relay_conn far_5_5133_1_b(.in(far_5_5133_0[1]), .out(far_5_5133_1[1]));
    assign layer_5[33] = ~far_5_5133_1[0] | (far_5_5133_1[0] & far_5_5133_1[1]); 
    wire [1:0] far_5_5134_0;    relay_conn far_5_5134_0_a(.in(layer_4[616]), .out(far_5_5134_0[0]));    relay_conn far_5_5134_0_b(.in(layer_4[538]), .out(far_5_5134_0[1]));
    wire [1:0] far_5_5134_1;    relay_conn far_5_5134_1_a(.in(far_5_5134_0[0]), .out(far_5_5134_1[0]));    relay_conn far_5_5134_1_b(.in(far_5_5134_0[1]), .out(far_5_5134_1[1]));
    assign layer_5[34] = far_5_5134_1[0] & far_5_5134_1[1]; 
    wire [1:0] far_5_5135_0;    relay_conn far_5_5135_0_a(.in(layer_4[589]), .out(far_5_5135_0[0]));    relay_conn far_5_5135_0_b(.in(layer_4[526]), .out(far_5_5135_0[1]));
    assign layer_5[35] = ~far_5_5135_0[1] | (far_5_5135_0[0] & far_5_5135_0[1]); 
    assign layer_5[36] = layer_4[958] | layer_4[986]; 
    assign layer_5[37] = layer_4[442] & ~layer_4[428]; 
    wire [1:0] far_5_5138_0;    relay_conn far_5_5138_0_a(.in(layer_4[952]), .out(far_5_5138_0[0]));    relay_conn far_5_5138_0_b(.in(layer_4[893]), .out(far_5_5138_0[1]));
    assign layer_5[38] = far_5_5138_0[0] | far_5_5138_0[1]; 
    wire [1:0] far_5_5139_0;    relay_conn far_5_5139_0_a(.in(layer_4[204]), .out(far_5_5139_0[0]));    relay_conn far_5_5139_0_b(.in(layer_4[106]), .out(far_5_5139_0[1]));
    wire [1:0] far_5_5139_1;    relay_conn far_5_5139_1_a(.in(far_5_5139_0[0]), .out(far_5_5139_1[0]));    relay_conn far_5_5139_1_b(.in(far_5_5139_0[1]), .out(far_5_5139_1[1]));
    wire [1:0] far_5_5139_2;    relay_conn far_5_5139_2_a(.in(far_5_5139_1[0]), .out(far_5_5139_2[0]));    relay_conn far_5_5139_2_b(.in(far_5_5139_1[1]), .out(far_5_5139_2[1]));
    assign layer_5[39] = far_5_5139_2[0] & ~far_5_5139_2[1]; 
    wire [1:0] far_5_5140_0;    relay_conn far_5_5140_0_a(.in(layer_4[526]), .out(far_5_5140_0[0]));    relay_conn far_5_5140_0_b(.in(layer_4[424]), .out(far_5_5140_0[1]));
    wire [1:0] far_5_5140_1;    relay_conn far_5_5140_1_a(.in(far_5_5140_0[0]), .out(far_5_5140_1[0]));    relay_conn far_5_5140_1_b(.in(far_5_5140_0[1]), .out(far_5_5140_1[1]));
    wire [1:0] far_5_5140_2;    relay_conn far_5_5140_2_a(.in(far_5_5140_1[0]), .out(far_5_5140_2[0]));    relay_conn far_5_5140_2_b(.in(far_5_5140_1[1]), .out(far_5_5140_2[1]));
    assign layer_5[40] = ~far_5_5140_2[1] | (far_5_5140_2[0] & far_5_5140_2[1]); 
    wire [1:0] far_5_5141_0;    relay_conn far_5_5141_0_a(.in(layer_4[107]), .out(far_5_5141_0[0]));    relay_conn far_5_5141_0_b(.in(layer_4[174]), .out(far_5_5141_0[1]));
    wire [1:0] far_5_5141_1;    relay_conn far_5_5141_1_a(.in(far_5_5141_0[0]), .out(far_5_5141_1[0]));    relay_conn far_5_5141_1_b(.in(far_5_5141_0[1]), .out(far_5_5141_1[1]));
    assign layer_5[41] = far_5_5141_1[0] & far_5_5141_1[1]; 
    assign layer_5[42] = layer_4[300]; 
    wire [1:0] far_5_5143_0;    relay_conn far_5_5143_0_a(.in(layer_4[527]), .out(far_5_5143_0[0]));    relay_conn far_5_5143_0_b(.in(layer_4[443]), .out(far_5_5143_0[1]));
    wire [1:0] far_5_5143_1;    relay_conn far_5_5143_1_a(.in(far_5_5143_0[0]), .out(far_5_5143_1[0]));    relay_conn far_5_5143_1_b(.in(far_5_5143_0[1]), .out(far_5_5143_1[1]));
    assign layer_5[43] = far_5_5143_1[1] & ~far_5_5143_1[0]; 
    wire [1:0] far_5_5144_0;    relay_conn far_5_5144_0_a(.in(layer_4[226]), .out(far_5_5144_0[0]));    relay_conn far_5_5144_0_b(.in(layer_4[167]), .out(far_5_5144_0[1]));
    assign layer_5[44] = far_5_5144_0[1] & ~far_5_5144_0[0]; 
    wire [1:0] far_5_5145_0;    relay_conn far_5_5145_0_a(.in(layer_4[358]), .out(far_5_5145_0[0]));    relay_conn far_5_5145_0_b(.in(layer_4[437]), .out(far_5_5145_0[1]));
    wire [1:0] far_5_5145_1;    relay_conn far_5_5145_1_a(.in(far_5_5145_0[0]), .out(far_5_5145_1[0]));    relay_conn far_5_5145_1_b(.in(far_5_5145_0[1]), .out(far_5_5145_1[1]));
    assign layer_5[45] = ~far_5_5145_1[1] | (far_5_5145_1[0] & far_5_5145_1[1]); 
    wire [1:0] far_5_5146_0;    relay_conn far_5_5146_0_a(.in(layer_4[813]), .out(far_5_5146_0[0]));    relay_conn far_5_5146_0_b(.in(layer_4[941]), .out(far_5_5146_0[1]));
    wire [1:0] far_5_5146_1;    relay_conn far_5_5146_1_a(.in(far_5_5146_0[0]), .out(far_5_5146_1[0]));    relay_conn far_5_5146_1_b(.in(far_5_5146_0[1]), .out(far_5_5146_1[1]));
    wire [1:0] far_5_5146_2;    relay_conn far_5_5146_2_a(.in(far_5_5146_1[0]), .out(far_5_5146_2[0]));    relay_conn far_5_5146_2_b(.in(far_5_5146_1[1]), .out(far_5_5146_2[1]));
    wire [1:0] far_5_5146_3;    relay_conn far_5_5146_3_a(.in(far_5_5146_2[0]), .out(far_5_5146_3[0]));    relay_conn far_5_5146_3_b(.in(far_5_5146_2[1]), .out(far_5_5146_3[1]));
    assign layer_5[46] = far_5_5146_3[1]; 
    wire [1:0] far_5_5147_0;    relay_conn far_5_5147_0_a(.in(layer_4[692]), .out(far_5_5147_0[0]));    relay_conn far_5_5147_0_b(.in(layer_4[643]), .out(far_5_5147_0[1]));
    assign layer_5[47] = ~far_5_5147_0[1] | (far_5_5147_0[0] & far_5_5147_0[1]); 
    wire [1:0] far_5_5148_0;    relay_conn far_5_5148_0_a(.in(layer_4[636]), .out(far_5_5148_0[0]));    relay_conn far_5_5148_0_b(.in(layer_4[707]), .out(far_5_5148_0[1]));
    wire [1:0] far_5_5148_1;    relay_conn far_5_5148_1_a(.in(far_5_5148_0[0]), .out(far_5_5148_1[0]));    relay_conn far_5_5148_1_b(.in(far_5_5148_0[1]), .out(far_5_5148_1[1]));
    assign layer_5[48] = ~(far_5_5148_1[0] | far_5_5148_1[1]); 
    wire [1:0] far_5_5149_0;    relay_conn far_5_5149_0_a(.in(layer_4[500]), .out(far_5_5149_0[0]));    relay_conn far_5_5149_0_b(.in(layer_4[556]), .out(far_5_5149_0[1]));
    assign layer_5[49] = ~far_5_5149_0[1]; 
    assign layer_5[50] = layer_4[632]; 
    wire [1:0] far_5_5151_0;    relay_conn far_5_5151_0_a(.in(layer_4[542]), .out(far_5_5151_0[0]));    relay_conn far_5_5151_0_b(.in(layer_4[654]), .out(far_5_5151_0[1]));
    wire [1:0] far_5_5151_1;    relay_conn far_5_5151_1_a(.in(far_5_5151_0[0]), .out(far_5_5151_1[0]));    relay_conn far_5_5151_1_b(.in(far_5_5151_0[1]), .out(far_5_5151_1[1]));
    wire [1:0] far_5_5151_2;    relay_conn far_5_5151_2_a(.in(far_5_5151_1[0]), .out(far_5_5151_2[0]));    relay_conn far_5_5151_2_b(.in(far_5_5151_1[1]), .out(far_5_5151_2[1]));
    assign layer_5[51] = ~far_5_5151_2[1]; 
    assign layer_5[52] = ~(layer_4[811] & layer_4[787]); 
    wire [1:0] far_5_5153_0;    relay_conn far_5_5153_0_a(.in(layer_4[4]), .out(far_5_5153_0[0]));    relay_conn far_5_5153_0_b(.in(layer_4[131]), .out(far_5_5153_0[1]));
    wire [1:0] far_5_5153_1;    relay_conn far_5_5153_1_a(.in(far_5_5153_0[0]), .out(far_5_5153_1[0]));    relay_conn far_5_5153_1_b(.in(far_5_5153_0[1]), .out(far_5_5153_1[1]));
    wire [1:0] far_5_5153_2;    relay_conn far_5_5153_2_a(.in(far_5_5153_1[0]), .out(far_5_5153_2[0]));    relay_conn far_5_5153_2_b(.in(far_5_5153_1[1]), .out(far_5_5153_2[1]));
    assign layer_5[53] = ~(far_5_5153_2[0] | far_5_5153_2[1]); 
    wire [1:0] far_5_5154_0;    relay_conn far_5_5154_0_a(.in(layer_4[158]), .out(far_5_5154_0[0]));    relay_conn far_5_5154_0_b(.in(layer_4[67]), .out(far_5_5154_0[1]));
    wire [1:0] far_5_5154_1;    relay_conn far_5_5154_1_a(.in(far_5_5154_0[0]), .out(far_5_5154_1[0]));    relay_conn far_5_5154_1_b(.in(far_5_5154_0[1]), .out(far_5_5154_1[1]));
    assign layer_5[54] = ~far_5_5154_1[0] | (far_5_5154_1[0] & far_5_5154_1[1]); 
    wire [1:0] far_5_5155_0;    relay_conn far_5_5155_0_a(.in(layer_4[104]), .out(far_5_5155_0[0]));    relay_conn far_5_5155_0_b(.in(layer_4[215]), .out(far_5_5155_0[1]));
    wire [1:0] far_5_5155_1;    relay_conn far_5_5155_1_a(.in(far_5_5155_0[0]), .out(far_5_5155_1[0]));    relay_conn far_5_5155_1_b(.in(far_5_5155_0[1]), .out(far_5_5155_1[1]));
    wire [1:0] far_5_5155_2;    relay_conn far_5_5155_2_a(.in(far_5_5155_1[0]), .out(far_5_5155_2[0]));    relay_conn far_5_5155_2_b(.in(far_5_5155_1[1]), .out(far_5_5155_2[1]));
    assign layer_5[55] = ~far_5_5155_2[1] | (far_5_5155_2[0] & far_5_5155_2[1]); 
    wire [1:0] far_5_5156_0;    relay_conn far_5_5156_0_a(.in(layer_4[669]), .out(far_5_5156_0[0]));    relay_conn far_5_5156_0_b(.in(layer_4[580]), .out(far_5_5156_0[1]));
    wire [1:0] far_5_5156_1;    relay_conn far_5_5156_1_a(.in(far_5_5156_0[0]), .out(far_5_5156_1[0]));    relay_conn far_5_5156_1_b(.in(far_5_5156_0[1]), .out(far_5_5156_1[1]));
    assign layer_5[56] = ~(far_5_5156_1[0] | far_5_5156_1[1]); 
    wire [1:0] far_5_5157_0;    relay_conn far_5_5157_0_a(.in(layer_4[573]), .out(far_5_5157_0[0]));    relay_conn far_5_5157_0_b(.in(layer_4[614]), .out(far_5_5157_0[1]));
    assign layer_5[57] = ~(far_5_5157_0[0] & far_5_5157_0[1]); 
    wire [1:0] far_5_5158_0;    relay_conn far_5_5158_0_a(.in(layer_4[559]), .out(far_5_5158_0[0]));    relay_conn far_5_5158_0_b(.in(layer_4[654]), .out(far_5_5158_0[1]));
    wire [1:0] far_5_5158_1;    relay_conn far_5_5158_1_a(.in(far_5_5158_0[0]), .out(far_5_5158_1[0]));    relay_conn far_5_5158_1_b(.in(far_5_5158_0[1]), .out(far_5_5158_1[1]));
    assign layer_5[58] = ~far_5_5158_1[0]; 
    wire [1:0] far_5_5159_0;    relay_conn far_5_5159_0_a(.in(layer_4[625]), .out(far_5_5159_0[0]));    relay_conn far_5_5159_0_b(.in(layer_4[676]), .out(far_5_5159_0[1]));
    assign layer_5[59] = ~far_5_5159_0[0]; 
    wire [1:0] far_5_5160_0;    relay_conn far_5_5160_0_a(.in(layer_4[901]), .out(far_5_5160_0[0]));    relay_conn far_5_5160_0_b(.in(layer_4[955]), .out(far_5_5160_0[1]));
    assign layer_5[60] = far_5_5160_0[0] & far_5_5160_0[1]; 
    wire [1:0] far_5_5161_0;    relay_conn far_5_5161_0_a(.in(layer_4[713]), .out(far_5_5161_0[0]));    relay_conn far_5_5161_0_b(.in(layer_4[666]), .out(far_5_5161_0[1]));
    assign layer_5[61] = ~far_5_5161_0[1]; 
    assign layer_5[62] = layer_4[772] | layer_4[789]; 
    wire [1:0] far_5_5163_0;    relay_conn far_5_5163_0_a(.in(layer_4[997]), .out(far_5_5163_0[0]));    relay_conn far_5_5163_0_b(.in(layer_4[947]), .out(far_5_5163_0[1]));
    assign layer_5[63] = ~far_5_5163_0[0]; 
    wire [1:0] far_5_5164_0;    relay_conn far_5_5164_0_a(.in(layer_4[874]), .out(far_5_5164_0[0]));    relay_conn far_5_5164_0_b(.in(layer_4[954]), .out(far_5_5164_0[1]));
    wire [1:0] far_5_5164_1;    relay_conn far_5_5164_1_a(.in(far_5_5164_0[0]), .out(far_5_5164_1[0]));    relay_conn far_5_5164_1_b(.in(far_5_5164_0[1]), .out(far_5_5164_1[1]));
    assign layer_5[64] = far_5_5164_1[0] & ~far_5_5164_1[1]; 
    wire [1:0] far_5_5165_0;    relay_conn far_5_5165_0_a(.in(layer_4[619]), .out(far_5_5165_0[0]));    relay_conn far_5_5165_0_b(.in(layer_4[580]), .out(far_5_5165_0[1]));
    assign layer_5[65] = ~far_5_5165_0[1]; 
    wire [1:0] far_5_5166_0;    relay_conn far_5_5166_0_a(.in(layer_4[787]), .out(far_5_5166_0[0]));    relay_conn far_5_5166_0_b(.in(layer_4[910]), .out(far_5_5166_0[1]));
    wire [1:0] far_5_5166_1;    relay_conn far_5_5166_1_a(.in(far_5_5166_0[0]), .out(far_5_5166_1[0]));    relay_conn far_5_5166_1_b(.in(far_5_5166_0[1]), .out(far_5_5166_1[1]));
    wire [1:0] far_5_5166_2;    relay_conn far_5_5166_2_a(.in(far_5_5166_1[0]), .out(far_5_5166_2[0]));    relay_conn far_5_5166_2_b(.in(far_5_5166_1[1]), .out(far_5_5166_2[1]));
    assign layer_5[66] = ~far_5_5166_2[1]; 
    wire [1:0] far_5_5167_0;    relay_conn far_5_5167_0_a(.in(layer_4[658]), .out(far_5_5167_0[0]));    relay_conn far_5_5167_0_b(.in(layer_4[743]), .out(far_5_5167_0[1]));
    wire [1:0] far_5_5167_1;    relay_conn far_5_5167_1_a(.in(far_5_5167_0[0]), .out(far_5_5167_1[0]));    relay_conn far_5_5167_1_b(.in(far_5_5167_0[1]), .out(far_5_5167_1[1]));
    assign layer_5[67] = far_5_5167_1[0]; 
    wire [1:0] far_5_5168_0;    relay_conn far_5_5168_0_a(.in(layer_4[928]), .out(far_5_5168_0[0]));    relay_conn far_5_5168_0_b(.in(layer_4[964]), .out(far_5_5168_0[1]));
    assign layer_5[68] = ~(far_5_5168_0[0] ^ far_5_5168_0[1]); 
    wire [1:0] far_5_5169_0;    relay_conn far_5_5169_0_a(.in(layer_4[381]), .out(far_5_5169_0[0]));    relay_conn far_5_5169_0_b(.in(layer_4[318]), .out(far_5_5169_0[1]));
    assign layer_5[69] = far_5_5169_0[1]; 
    wire [1:0] far_5_5170_0;    relay_conn far_5_5170_0_a(.in(layer_4[802]), .out(far_5_5170_0[0]));    relay_conn far_5_5170_0_b(.in(layer_4[726]), .out(far_5_5170_0[1]));
    wire [1:0] far_5_5170_1;    relay_conn far_5_5170_1_a(.in(far_5_5170_0[0]), .out(far_5_5170_1[0]));    relay_conn far_5_5170_1_b(.in(far_5_5170_0[1]), .out(far_5_5170_1[1]));
    assign layer_5[70] = ~far_5_5170_1[1] | (far_5_5170_1[0] & far_5_5170_1[1]); 
    wire [1:0] far_5_5171_0;    relay_conn far_5_5171_0_a(.in(layer_4[273]), .out(far_5_5171_0[0]));    relay_conn far_5_5171_0_b(.in(layer_4[219]), .out(far_5_5171_0[1]));
    assign layer_5[71] = ~(far_5_5171_0[0] & far_5_5171_0[1]); 
    wire [1:0] far_5_5172_0;    relay_conn far_5_5172_0_a(.in(layer_4[190]), .out(far_5_5172_0[0]));    relay_conn far_5_5172_0_b(.in(layer_4[127]), .out(far_5_5172_0[1]));
    assign layer_5[72] = far_5_5172_0[0] & ~far_5_5172_0[1]; 
    wire [1:0] far_5_5173_0;    relay_conn far_5_5173_0_a(.in(layer_4[789]), .out(far_5_5173_0[0]));    relay_conn far_5_5173_0_b(.in(layer_4[699]), .out(far_5_5173_0[1]));
    wire [1:0] far_5_5173_1;    relay_conn far_5_5173_1_a(.in(far_5_5173_0[0]), .out(far_5_5173_1[0]));    relay_conn far_5_5173_1_b(.in(far_5_5173_0[1]), .out(far_5_5173_1[1]));
    assign layer_5[73] = ~(far_5_5173_1[0] & far_5_5173_1[1]); 
    assign layer_5[74] = ~(layer_4[23] | layer_4[42]); 
    assign layer_5[75] = layer_4[386]; 
    assign layer_5[76] = ~(layer_4[18] | layer_4[45]); 
    wire [1:0] far_5_5177_0;    relay_conn far_5_5177_0_a(.in(layer_4[628]), .out(far_5_5177_0[0]));    relay_conn far_5_5177_0_b(.in(layer_4[713]), .out(far_5_5177_0[1]));
    wire [1:0] far_5_5177_1;    relay_conn far_5_5177_1_a(.in(far_5_5177_0[0]), .out(far_5_5177_1[0]));    relay_conn far_5_5177_1_b(.in(far_5_5177_0[1]), .out(far_5_5177_1[1]));
    assign layer_5[77] = far_5_5177_1[0] | far_5_5177_1[1]; 
    wire [1:0] far_5_5178_0;    relay_conn far_5_5178_0_a(.in(layer_4[92]), .out(far_5_5178_0[0]));    relay_conn far_5_5178_0_b(.in(layer_4[176]), .out(far_5_5178_0[1]));
    wire [1:0] far_5_5178_1;    relay_conn far_5_5178_1_a(.in(far_5_5178_0[0]), .out(far_5_5178_1[0]));    relay_conn far_5_5178_1_b(.in(far_5_5178_0[1]), .out(far_5_5178_1[1]));
    assign layer_5[78] = ~far_5_5178_1[0]; 
    assign layer_5[79] = ~layer_4[902] | (layer_4[928] & layer_4[902]); 
    assign layer_5[80] = layer_4[424]; 
    assign layer_5[81] = layer_4[921] | layer_4[941]; 
    assign layer_5[82] = ~layer_4[407]; 
    assign layer_5[83] = ~(layer_4[248] & layer_4[228]); 
    wire [1:0] far_5_5184_0;    relay_conn far_5_5184_0_a(.in(layer_4[836]), .out(far_5_5184_0[0]));    relay_conn far_5_5184_0_b(.in(layer_4[900]), .out(far_5_5184_0[1]));
    wire [1:0] far_5_5184_1;    relay_conn far_5_5184_1_a(.in(far_5_5184_0[0]), .out(far_5_5184_1[0]));    relay_conn far_5_5184_1_b(.in(far_5_5184_0[1]), .out(far_5_5184_1[1]));
    assign layer_5[84] = ~far_5_5184_1[1]; 
    wire [1:0] far_5_5185_0;    relay_conn far_5_5185_0_a(.in(layer_4[839]), .out(far_5_5185_0[0]));    relay_conn far_5_5185_0_b(.in(layer_4[875]), .out(far_5_5185_0[1]));
    assign layer_5[85] = far_5_5185_0[0] & ~far_5_5185_0[1]; 
    wire [1:0] far_5_5186_0;    relay_conn far_5_5186_0_a(.in(layer_4[330]), .out(far_5_5186_0[0]));    relay_conn far_5_5186_0_b(.in(layer_4[253]), .out(far_5_5186_0[1]));
    wire [1:0] far_5_5186_1;    relay_conn far_5_5186_1_a(.in(far_5_5186_0[0]), .out(far_5_5186_1[0]));    relay_conn far_5_5186_1_b(.in(far_5_5186_0[1]), .out(far_5_5186_1[1]));
    assign layer_5[86] = far_5_5186_1[0] | far_5_5186_1[1]; 
    wire [1:0] far_5_5187_0;    relay_conn far_5_5187_0_a(.in(layer_4[106]), .out(far_5_5187_0[0]));    relay_conn far_5_5187_0_b(.in(layer_4[12]), .out(far_5_5187_0[1]));
    wire [1:0] far_5_5187_1;    relay_conn far_5_5187_1_a(.in(far_5_5187_0[0]), .out(far_5_5187_1[0]));    relay_conn far_5_5187_1_b(.in(far_5_5187_0[1]), .out(far_5_5187_1[1]));
    assign layer_5[87] = ~(far_5_5187_1[0] ^ far_5_5187_1[1]); 
    wire [1:0] far_5_5188_0;    relay_conn far_5_5188_0_a(.in(layer_4[704]), .out(far_5_5188_0[0]));    relay_conn far_5_5188_0_b(.in(layer_4[787]), .out(far_5_5188_0[1]));
    wire [1:0] far_5_5188_1;    relay_conn far_5_5188_1_a(.in(far_5_5188_0[0]), .out(far_5_5188_1[0]));    relay_conn far_5_5188_1_b(.in(far_5_5188_0[1]), .out(far_5_5188_1[1]));
    assign layer_5[88] = ~(far_5_5188_1[0] | far_5_5188_1[1]); 
    assign layer_5[89] = layer_4[657]; 
    wire [1:0] far_5_5190_0;    relay_conn far_5_5190_0_a(.in(layer_4[894]), .out(far_5_5190_0[0]));    relay_conn far_5_5190_0_b(.in(layer_4[995]), .out(far_5_5190_0[1]));
    wire [1:0] far_5_5190_1;    relay_conn far_5_5190_1_a(.in(far_5_5190_0[0]), .out(far_5_5190_1[0]));    relay_conn far_5_5190_1_b(.in(far_5_5190_0[1]), .out(far_5_5190_1[1]));
    wire [1:0] far_5_5190_2;    relay_conn far_5_5190_2_a(.in(far_5_5190_1[0]), .out(far_5_5190_2[0]));    relay_conn far_5_5190_2_b(.in(far_5_5190_1[1]), .out(far_5_5190_2[1]));
    assign layer_5[90] = far_5_5190_2[0] | far_5_5190_2[1]; 
    wire [1:0] far_5_5191_0;    relay_conn far_5_5191_0_a(.in(layer_4[656]), .out(far_5_5191_0[0]));    relay_conn far_5_5191_0_b(.in(layer_4[606]), .out(far_5_5191_0[1]));
    assign layer_5[91] = ~(far_5_5191_0[0] | far_5_5191_0[1]); 
    wire [1:0] far_5_5192_0;    relay_conn far_5_5192_0_a(.in(layer_4[719]), .out(far_5_5192_0[0]));    relay_conn far_5_5192_0_b(.in(layer_4[672]), .out(far_5_5192_0[1]));
    assign layer_5[92] = far_5_5192_0[0]; 
    wire [1:0] far_5_5193_0;    relay_conn far_5_5193_0_a(.in(layer_4[900]), .out(far_5_5193_0[0]));    relay_conn far_5_5193_0_b(.in(layer_4[954]), .out(far_5_5193_0[1]));
    assign layer_5[93] = ~far_5_5193_0[1] | (far_5_5193_0[0] & far_5_5193_0[1]); 
    assign layer_5[94] = layer_4[107] & ~layer_4[129]; 
    wire [1:0] far_5_5195_0;    relay_conn far_5_5195_0_a(.in(layer_4[145]), .out(far_5_5195_0[0]));    relay_conn far_5_5195_0_b(.in(layer_4[223]), .out(far_5_5195_0[1]));
    wire [1:0] far_5_5195_1;    relay_conn far_5_5195_1_a(.in(far_5_5195_0[0]), .out(far_5_5195_1[0]));    relay_conn far_5_5195_1_b(.in(far_5_5195_0[1]), .out(far_5_5195_1[1]));
    assign layer_5[95] = far_5_5195_1[1]; 
    wire [1:0] far_5_5196_0;    relay_conn far_5_5196_0_a(.in(layer_4[728]), .out(far_5_5196_0[0]));    relay_conn far_5_5196_0_b(.in(layer_4[620]), .out(far_5_5196_0[1]));
    wire [1:0] far_5_5196_1;    relay_conn far_5_5196_1_a(.in(far_5_5196_0[0]), .out(far_5_5196_1[0]));    relay_conn far_5_5196_1_b(.in(far_5_5196_0[1]), .out(far_5_5196_1[1]));
    wire [1:0] far_5_5196_2;    relay_conn far_5_5196_2_a(.in(far_5_5196_1[0]), .out(far_5_5196_2[0]));    relay_conn far_5_5196_2_b(.in(far_5_5196_1[1]), .out(far_5_5196_2[1]));
    assign layer_5[96] = ~far_5_5196_2[1]; 
    wire [1:0] far_5_5197_0;    relay_conn far_5_5197_0_a(.in(layer_4[107]), .out(far_5_5197_0[0]));    relay_conn far_5_5197_0_b(.in(layer_4[158]), .out(far_5_5197_0[1]));
    assign layer_5[97] = ~far_5_5197_0[0]; 
    wire [1:0] far_5_5198_0;    relay_conn far_5_5198_0_a(.in(layer_4[754]), .out(far_5_5198_0[0]));    relay_conn far_5_5198_0_b(.in(layer_4[670]), .out(far_5_5198_0[1]));
    wire [1:0] far_5_5198_1;    relay_conn far_5_5198_1_a(.in(far_5_5198_0[0]), .out(far_5_5198_1[0]));    relay_conn far_5_5198_1_b(.in(far_5_5198_0[1]), .out(far_5_5198_1[1]));
    assign layer_5[98] = far_5_5198_1[0] & ~far_5_5198_1[1]; 
    assign layer_5[99] = ~layer_4[994]; 
    assign layer_5[100] = ~layer_4[526]; 
    wire [1:0] far_5_5201_0;    relay_conn far_5_5201_0_a(.in(layer_4[884]), .out(far_5_5201_0[0]));    relay_conn far_5_5201_0_b(.in(layer_4[973]), .out(far_5_5201_0[1]));
    wire [1:0] far_5_5201_1;    relay_conn far_5_5201_1_a(.in(far_5_5201_0[0]), .out(far_5_5201_1[0]));    relay_conn far_5_5201_1_b(.in(far_5_5201_0[1]), .out(far_5_5201_1[1]));
    assign layer_5[101] = ~far_5_5201_1[0]; 
    assign layer_5[102] = ~layer_4[806] | (layer_4[806] & layer_4[794]); 
    wire [1:0] far_5_5203_0;    relay_conn far_5_5203_0_a(.in(layer_4[588]), .out(far_5_5203_0[0]));    relay_conn far_5_5203_0_b(.in(layer_4[518]), .out(far_5_5203_0[1]));
    wire [1:0] far_5_5203_1;    relay_conn far_5_5203_1_a(.in(far_5_5203_0[0]), .out(far_5_5203_1[0]));    relay_conn far_5_5203_1_b(.in(far_5_5203_0[1]), .out(far_5_5203_1[1]));
    assign layer_5[103] = far_5_5203_1[0] & ~far_5_5203_1[1]; 
    wire [1:0] far_5_5204_0;    relay_conn far_5_5204_0_a(.in(layer_4[412]), .out(far_5_5204_0[0]));    relay_conn far_5_5204_0_b(.in(layer_4[470]), .out(far_5_5204_0[1]));
    assign layer_5[104] = ~far_5_5204_0[0]; 
    wire [1:0] far_5_5205_0;    relay_conn far_5_5205_0_a(.in(layer_4[577]), .out(far_5_5205_0[0]));    relay_conn far_5_5205_0_b(.in(layer_4[666]), .out(far_5_5205_0[1]));
    wire [1:0] far_5_5205_1;    relay_conn far_5_5205_1_a(.in(far_5_5205_0[0]), .out(far_5_5205_1[0]));    relay_conn far_5_5205_1_b(.in(far_5_5205_0[1]), .out(far_5_5205_1[1]));
    assign layer_5[105] = ~far_5_5205_1[0] | (far_5_5205_1[0] & far_5_5205_1[1]); 
    wire [1:0] far_5_5206_0;    relay_conn far_5_5206_0_a(.in(layer_4[66]), .out(far_5_5206_0[0]));    relay_conn far_5_5206_0_b(.in(layer_4[124]), .out(far_5_5206_0[1]));
    assign layer_5[106] = far_5_5206_0[0]; 
    wire [1:0] far_5_5207_0;    relay_conn far_5_5207_0_a(.in(layer_4[1000]), .out(far_5_5207_0[0]));    relay_conn far_5_5207_0_b(.in(layer_4[902]), .out(far_5_5207_0[1]));
    wire [1:0] far_5_5207_1;    relay_conn far_5_5207_1_a(.in(far_5_5207_0[0]), .out(far_5_5207_1[0]));    relay_conn far_5_5207_1_b(.in(far_5_5207_0[1]), .out(far_5_5207_1[1]));
    wire [1:0] far_5_5207_2;    relay_conn far_5_5207_2_a(.in(far_5_5207_1[0]), .out(far_5_5207_2[0]));    relay_conn far_5_5207_2_b(.in(far_5_5207_1[1]), .out(far_5_5207_2[1]));
    assign layer_5[107] = far_5_5207_2[0] ^ far_5_5207_2[1]; 
    wire [1:0] far_5_5208_0;    relay_conn far_5_5208_0_a(.in(layer_4[253]), .out(far_5_5208_0[0]));    relay_conn far_5_5208_0_b(.in(layer_4[322]), .out(far_5_5208_0[1]));
    wire [1:0] far_5_5208_1;    relay_conn far_5_5208_1_a(.in(far_5_5208_0[0]), .out(far_5_5208_1[0]));    relay_conn far_5_5208_1_b(.in(far_5_5208_0[1]), .out(far_5_5208_1[1]));
    assign layer_5[108] = far_5_5208_1[1] & ~far_5_5208_1[0]; 
    wire [1:0] far_5_5209_0;    relay_conn far_5_5209_0_a(.in(layer_4[789]), .out(far_5_5209_0[0]));    relay_conn far_5_5209_0_b(.in(layer_4[858]), .out(far_5_5209_0[1]));
    wire [1:0] far_5_5209_1;    relay_conn far_5_5209_1_a(.in(far_5_5209_0[0]), .out(far_5_5209_1[0]));    relay_conn far_5_5209_1_b(.in(far_5_5209_0[1]), .out(far_5_5209_1[1]));
    assign layer_5[109] = ~far_5_5209_1[1]; 
    wire [1:0] far_5_5210_0;    relay_conn far_5_5210_0_a(.in(layer_4[608]), .out(far_5_5210_0[0]));    relay_conn far_5_5210_0_b(.in(layer_4[656]), .out(far_5_5210_0[1]));
    assign layer_5[110] = ~(far_5_5210_0[0] & far_5_5210_0[1]); 
    wire [1:0] far_5_5211_0;    relay_conn far_5_5211_0_a(.in(layer_4[830]), .out(far_5_5211_0[0]));    relay_conn far_5_5211_0_b(.in(layer_4[893]), .out(far_5_5211_0[1]));
    assign layer_5[111] = ~(far_5_5211_0[0] | far_5_5211_0[1]); 
    assign layer_5[112] = ~layer_4[827]; 
    wire [1:0] far_5_5213_0;    relay_conn far_5_5213_0_a(.in(layer_4[250]), .out(far_5_5213_0[0]));    relay_conn far_5_5213_0_b(.in(layer_4[309]), .out(far_5_5213_0[1]));
    assign layer_5[113] = far_5_5213_0[0] ^ far_5_5213_0[1]; 
    assign layer_5[114] = ~layer_4[831]; 
    wire [1:0] far_5_5215_0;    relay_conn far_5_5215_0_a(.in(layer_4[515]), .out(far_5_5215_0[0]));    relay_conn far_5_5215_0_b(.in(layer_4[554]), .out(far_5_5215_0[1]));
    assign layer_5[115] = far_5_5215_0[0] & far_5_5215_0[1]; 
    assign layer_5[116] = layer_4[62] & ~layer_4[47]; 
    wire [1:0] far_5_5217_0;    relay_conn far_5_5217_0_a(.in(layer_4[719]), .out(far_5_5217_0[0]));    relay_conn far_5_5217_0_b(.in(layer_4[657]), .out(far_5_5217_0[1]));
    assign layer_5[117] = ~far_5_5217_0[0]; 
    wire [1:0] far_5_5218_0;    relay_conn far_5_5218_0_a(.in(layer_4[337]), .out(far_5_5218_0[0]));    relay_conn far_5_5218_0_b(.in(layer_4[210]), .out(far_5_5218_0[1]));
    wire [1:0] far_5_5218_1;    relay_conn far_5_5218_1_a(.in(far_5_5218_0[0]), .out(far_5_5218_1[0]));    relay_conn far_5_5218_1_b(.in(far_5_5218_0[1]), .out(far_5_5218_1[1]));
    wire [1:0] far_5_5218_2;    relay_conn far_5_5218_2_a(.in(far_5_5218_1[0]), .out(far_5_5218_2[0]));    relay_conn far_5_5218_2_b(.in(far_5_5218_1[1]), .out(far_5_5218_2[1]));
    assign layer_5[118] = far_5_5218_2[0] | far_5_5218_2[1]; 
    wire [1:0] far_5_5219_0;    relay_conn far_5_5219_0_a(.in(layer_4[104]), .out(far_5_5219_0[0]));    relay_conn far_5_5219_0_b(.in(layer_4[149]), .out(far_5_5219_0[1]));
    assign layer_5[119] = ~(far_5_5219_0[0] ^ far_5_5219_0[1]); 
    wire [1:0] far_5_5220_0;    relay_conn far_5_5220_0_a(.in(layer_4[42]), .out(far_5_5220_0[0]));    relay_conn far_5_5220_0_b(.in(layer_4[142]), .out(far_5_5220_0[1]));
    wire [1:0] far_5_5220_1;    relay_conn far_5_5220_1_a(.in(far_5_5220_0[0]), .out(far_5_5220_1[0]));    relay_conn far_5_5220_1_b(.in(far_5_5220_0[1]), .out(far_5_5220_1[1]));
    wire [1:0] far_5_5220_2;    relay_conn far_5_5220_2_a(.in(far_5_5220_1[0]), .out(far_5_5220_2[0]));    relay_conn far_5_5220_2_b(.in(far_5_5220_1[1]), .out(far_5_5220_2[1]));
    assign layer_5[120] = far_5_5220_2[0] | far_5_5220_2[1]; 
    wire [1:0] far_5_5221_0;    relay_conn far_5_5221_0_a(.in(layer_4[833]), .out(far_5_5221_0[0]));    relay_conn far_5_5221_0_b(.in(layer_4[958]), .out(far_5_5221_0[1]));
    wire [1:0] far_5_5221_1;    relay_conn far_5_5221_1_a(.in(far_5_5221_0[0]), .out(far_5_5221_1[0]));    relay_conn far_5_5221_1_b(.in(far_5_5221_0[1]), .out(far_5_5221_1[1]));
    wire [1:0] far_5_5221_2;    relay_conn far_5_5221_2_a(.in(far_5_5221_1[0]), .out(far_5_5221_2[0]));    relay_conn far_5_5221_2_b(.in(far_5_5221_1[1]), .out(far_5_5221_2[1]));
    assign layer_5[121] = ~far_5_5221_2[0] | (far_5_5221_2[0] & far_5_5221_2[1]); 
    wire [1:0] far_5_5222_0;    relay_conn far_5_5222_0_a(.in(layer_4[253]), .out(far_5_5222_0[0]));    relay_conn far_5_5222_0_b(.in(layer_4[170]), .out(far_5_5222_0[1]));
    wire [1:0] far_5_5222_1;    relay_conn far_5_5222_1_a(.in(far_5_5222_0[0]), .out(far_5_5222_1[0]));    relay_conn far_5_5222_1_b(.in(far_5_5222_0[1]), .out(far_5_5222_1[1]));
    assign layer_5[122] = far_5_5222_1[0]; 
    wire [1:0] far_5_5223_0;    relay_conn far_5_5223_0_a(.in(layer_4[826]), .out(far_5_5223_0[0]));    relay_conn far_5_5223_0_b(.in(layer_4[922]), .out(far_5_5223_0[1]));
    wire [1:0] far_5_5223_1;    relay_conn far_5_5223_1_a(.in(far_5_5223_0[0]), .out(far_5_5223_1[0]));    relay_conn far_5_5223_1_b(.in(far_5_5223_0[1]), .out(far_5_5223_1[1]));
    wire [1:0] far_5_5223_2;    relay_conn far_5_5223_2_a(.in(far_5_5223_1[0]), .out(far_5_5223_2[0]));    relay_conn far_5_5223_2_b(.in(far_5_5223_1[1]), .out(far_5_5223_2[1]));
    assign layer_5[123] = far_5_5223_2[0] | far_5_5223_2[1]; 
    wire [1:0] far_5_5224_0;    relay_conn far_5_5224_0_a(.in(layer_4[785]), .out(far_5_5224_0[0]));    relay_conn far_5_5224_0_b(.in(layer_4[913]), .out(far_5_5224_0[1]));
    wire [1:0] far_5_5224_1;    relay_conn far_5_5224_1_a(.in(far_5_5224_0[0]), .out(far_5_5224_1[0]));    relay_conn far_5_5224_1_b(.in(far_5_5224_0[1]), .out(far_5_5224_1[1]));
    wire [1:0] far_5_5224_2;    relay_conn far_5_5224_2_a(.in(far_5_5224_1[0]), .out(far_5_5224_2[0]));    relay_conn far_5_5224_2_b(.in(far_5_5224_1[1]), .out(far_5_5224_2[1]));
    wire [1:0] far_5_5224_3;    relay_conn far_5_5224_3_a(.in(far_5_5224_2[0]), .out(far_5_5224_3[0]));    relay_conn far_5_5224_3_b(.in(far_5_5224_2[1]), .out(far_5_5224_3[1]));
    assign layer_5[124] = ~far_5_5224_3[1] | (far_5_5224_3[0] & far_5_5224_3[1]); 
    assign layer_5[125] = ~(layer_4[232] | layer_4[247]); 
    wire [1:0] far_5_5226_0;    relay_conn far_5_5226_0_a(.in(layer_4[725]), .out(far_5_5226_0[0]));    relay_conn far_5_5226_0_b(.in(layer_4[665]), .out(far_5_5226_0[1]));
    assign layer_5[126] = far_5_5226_0[1] & ~far_5_5226_0[0]; 
    assign layer_5[127] = layer_4[947]; 
    wire [1:0] far_5_5228_0;    relay_conn far_5_5228_0_a(.in(layer_4[969]), .out(far_5_5228_0[0]));    relay_conn far_5_5228_0_b(.in(layer_4[921]), .out(far_5_5228_0[1]));
    assign layer_5[128] = far_5_5228_0[0] & far_5_5228_0[1]; 
    wire [1:0] far_5_5229_0;    relay_conn far_5_5229_0_a(.in(layer_4[1019]), .out(far_5_5229_0[0]));    relay_conn far_5_5229_0_b(.in(layer_4[960]), .out(far_5_5229_0[1]));
    assign layer_5[129] = ~far_5_5229_0[1] | (far_5_5229_0[0] & far_5_5229_0[1]); 
    wire [1:0] far_5_5230_0;    relay_conn far_5_5230_0_a(.in(layer_4[84]), .out(far_5_5230_0[0]));    relay_conn far_5_5230_0_b(.in(layer_4[185]), .out(far_5_5230_0[1]));
    wire [1:0] far_5_5230_1;    relay_conn far_5_5230_1_a(.in(far_5_5230_0[0]), .out(far_5_5230_1[0]));    relay_conn far_5_5230_1_b(.in(far_5_5230_0[1]), .out(far_5_5230_1[1]));
    wire [1:0] far_5_5230_2;    relay_conn far_5_5230_2_a(.in(far_5_5230_1[0]), .out(far_5_5230_2[0]));    relay_conn far_5_5230_2_b(.in(far_5_5230_1[1]), .out(far_5_5230_2[1]));
    assign layer_5[130] = ~(far_5_5230_2[0] & far_5_5230_2[1]); 
    wire [1:0] far_5_5231_0;    relay_conn far_5_5231_0_a(.in(layer_4[10]), .out(far_5_5231_0[0]));    relay_conn far_5_5231_0_b(.in(layer_4[134]), .out(far_5_5231_0[1]));
    wire [1:0] far_5_5231_1;    relay_conn far_5_5231_1_a(.in(far_5_5231_0[0]), .out(far_5_5231_1[0]));    relay_conn far_5_5231_1_b(.in(far_5_5231_0[1]), .out(far_5_5231_1[1]));
    wire [1:0] far_5_5231_2;    relay_conn far_5_5231_2_a(.in(far_5_5231_1[0]), .out(far_5_5231_2[0]));    relay_conn far_5_5231_2_b(.in(far_5_5231_1[1]), .out(far_5_5231_2[1]));
    assign layer_5[131] = ~(far_5_5231_2[0] | far_5_5231_2[1]); 
    wire [1:0] far_5_5232_0;    relay_conn far_5_5232_0_a(.in(layer_4[462]), .out(far_5_5232_0[0]));    relay_conn far_5_5232_0_b(.in(layer_4[589]), .out(far_5_5232_0[1]));
    wire [1:0] far_5_5232_1;    relay_conn far_5_5232_1_a(.in(far_5_5232_0[0]), .out(far_5_5232_1[0]));    relay_conn far_5_5232_1_b(.in(far_5_5232_0[1]), .out(far_5_5232_1[1]));
    wire [1:0] far_5_5232_2;    relay_conn far_5_5232_2_a(.in(far_5_5232_1[0]), .out(far_5_5232_2[0]));    relay_conn far_5_5232_2_b(.in(far_5_5232_1[1]), .out(far_5_5232_2[1]));
    assign layer_5[132] = far_5_5232_2[1] & ~far_5_5232_2[0]; 
    wire [1:0] far_5_5233_0;    relay_conn far_5_5233_0_a(.in(layer_4[813]), .out(far_5_5233_0[0]));    relay_conn far_5_5233_0_b(.in(layer_4[690]), .out(far_5_5233_0[1]));
    wire [1:0] far_5_5233_1;    relay_conn far_5_5233_1_a(.in(far_5_5233_0[0]), .out(far_5_5233_1[0]));    relay_conn far_5_5233_1_b(.in(far_5_5233_0[1]), .out(far_5_5233_1[1]));
    wire [1:0] far_5_5233_2;    relay_conn far_5_5233_2_a(.in(far_5_5233_1[0]), .out(far_5_5233_2[0]));    relay_conn far_5_5233_2_b(.in(far_5_5233_1[1]), .out(far_5_5233_2[1]));
    assign layer_5[133] = far_5_5233_2[0] ^ far_5_5233_2[1]; 
    wire [1:0] far_5_5234_0;    relay_conn far_5_5234_0_a(.in(layer_4[636]), .out(far_5_5234_0[0]));    relay_conn far_5_5234_0_b(.in(layer_4[597]), .out(far_5_5234_0[1]));
    assign layer_5[134] = ~far_5_5234_0[0]; 
    assign layer_5[135] = layer_4[29]; 
    wire [1:0] far_5_5236_0;    relay_conn far_5_5236_0_a(.in(layer_4[755]), .out(far_5_5236_0[0]));    relay_conn far_5_5236_0_b(.in(layer_4[839]), .out(far_5_5236_0[1]));
    wire [1:0] far_5_5236_1;    relay_conn far_5_5236_1_a(.in(far_5_5236_0[0]), .out(far_5_5236_1[0]));    relay_conn far_5_5236_1_b(.in(far_5_5236_0[1]), .out(far_5_5236_1[1]));
    assign layer_5[136] = far_5_5236_1[0]; 
    wire [1:0] far_5_5237_0;    relay_conn far_5_5237_0_a(.in(layer_4[867]), .out(far_5_5237_0[0]));    relay_conn far_5_5237_0_b(.in(layer_4[930]), .out(far_5_5237_0[1]));
    assign layer_5[137] = far_5_5237_0[0] & ~far_5_5237_0[1]; 
    assign layer_5[138] = ~layer_4[387]; 
    assign layer_5[139] = layer_4[768] | layer_4[799]; 
    wire [1:0] far_5_5240_0;    relay_conn far_5_5240_0_a(.in(layer_4[962]), .out(far_5_5240_0[0]));    relay_conn far_5_5240_0_b(.in(layer_4[906]), .out(far_5_5240_0[1]));
    assign layer_5[140] = ~(far_5_5240_0[0] & far_5_5240_0[1]); 
    wire [1:0] far_5_5241_0;    relay_conn far_5_5241_0_a(.in(layer_4[9]), .out(far_5_5241_0[0]));    relay_conn far_5_5241_0_b(.in(layer_4[84]), .out(far_5_5241_0[1]));
    wire [1:0] far_5_5241_1;    relay_conn far_5_5241_1_a(.in(far_5_5241_0[0]), .out(far_5_5241_1[0]));    relay_conn far_5_5241_1_b(.in(far_5_5241_0[1]), .out(far_5_5241_1[1]));
    assign layer_5[141] = ~(far_5_5241_1[0] & far_5_5241_1[1]); 
    wire [1:0] far_5_5242_0;    relay_conn far_5_5242_0_a(.in(layer_4[536]), .out(far_5_5242_0[0]));    relay_conn far_5_5242_0_b(.in(layer_4[608]), .out(far_5_5242_0[1]));
    wire [1:0] far_5_5242_1;    relay_conn far_5_5242_1_a(.in(far_5_5242_0[0]), .out(far_5_5242_1[0]));    relay_conn far_5_5242_1_b(.in(far_5_5242_0[1]), .out(far_5_5242_1[1]));
    assign layer_5[142] = ~far_5_5242_1[1]; 
    wire [1:0] far_5_5243_0;    relay_conn far_5_5243_0_a(.in(layer_4[955]), .out(far_5_5243_0[0]));    relay_conn far_5_5243_0_b(.in(layer_4[888]), .out(far_5_5243_0[1]));
    wire [1:0] far_5_5243_1;    relay_conn far_5_5243_1_a(.in(far_5_5243_0[0]), .out(far_5_5243_1[0]));    relay_conn far_5_5243_1_b(.in(far_5_5243_0[1]), .out(far_5_5243_1[1]));
    assign layer_5[143] = far_5_5243_1[0] | far_5_5243_1[1]; 
    wire [1:0] far_5_5244_0;    relay_conn far_5_5244_0_a(.in(layer_4[497]), .out(far_5_5244_0[0]));    relay_conn far_5_5244_0_b(.in(layer_4[559]), .out(far_5_5244_0[1]));
    assign layer_5[144] = ~far_5_5244_0[0]; 
    wire [1:0] far_5_5245_0;    relay_conn far_5_5245_0_a(.in(layer_4[674]), .out(far_5_5245_0[0]));    relay_conn far_5_5245_0_b(.in(layer_4[775]), .out(far_5_5245_0[1]));
    wire [1:0] far_5_5245_1;    relay_conn far_5_5245_1_a(.in(far_5_5245_0[0]), .out(far_5_5245_1[0]));    relay_conn far_5_5245_1_b(.in(far_5_5245_0[1]), .out(far_5_5245_1[1]));
    wire [1:0] far_5_5245_2;    relay_conn far_5_5245_2_a(.in(far_5_5245_1[0]), .out(far_5_5245_2[0]));    relay_conn far_5_5245_2_b(.in(far_5_5245_1[1]), .out(far_5_5245_2[1]));
    assign layer_5[145] = ~far_5_5245_2[0]; 
    assign layer_5[146] = ~layer_4[65] | (layer_4[65] & layer_4[45]); 
    wire [1:0] far_5_5247_0;    relay_conn far_5_5247_0_a(.in(layer_4[437]), .out(far_5_5247_0[0]));    relay_conn far_5_5247_0_b(.in(layer_4[363]), .out(far_5_5247_0[1]));
    wire [1:0] far_5_5247_1;    relay_conn far_5_5247_1_a(.in(far_5_5247_0[0]), .out(far_5_5247_1[0]));    relay_conn far_5_5247_1_b(.in(far_5_5247_0[1]), .out(far_5_5247_1[1]));
    assign layer_5[147] = ~(far_5_5247_1[0] | far_5_5247_1[1]); 
    wire [1:0] far_5_5248_0;    relay_conn far_5_5248_0_a(.in(layer_4[89]), .out(far_5_5248_0[0]));    relay_conn far_5_5248_0_b(.in(layer_4[214]), .out(far_5_5248_0[1]));
    wire [1:0] far_5_5248_1;    relay_conn far_5_5248_1_a(.in(far_5_5248_0[0]), .out(far_5_5248_1[0]));    relay_conn far_5_5248_1_b(.in(far_5_5248_0[1]), .out(far_5_5248_1[1]));
    wire [1:0] far_5_5248_2;    relay_conn far_5_5248_2_a(.in(far_5_5248_1[0]), .out(far_5_5248_2[0]));    relay_conn far_5_5248_2_b(.in(far_5_5248_1[1]), .out(far_5_5248_2[1]));
    assign layer_5[148] = far_5_5248_2[0] & far_5_5248_2[1]; 
    wire [1:0] far_5_5249_0;    relay_conn far_5_5249_0_a(.in(layer_4[307]), .out(far_5_5249_0[0]));    relay_conn far_5_5249_0_b(.in(layer_4[245]), .out(far_5_5249_0[1]));
    assign layer_5[149] = ~(far_5_5249_0[0] & far_5_5249_0[1]); 
    assign layer_5[150] = layer_4[980]; 
    assign layer_5[151] = ~layer_4[980] | (layer_4[980] & layer_4[998]); 
    wire [1:0] far_5_5252_0;    relay_conn far_5_5252_0_a(.in(layer_4[795]), .out(far_5_5252_0[0]));    relay_conn far_5_5252_0_b(.in(layer_4[830]), .out(far_5_5252_0[1]));
    assign layer_5[152] = ~(far_5_5252_0[0] | far_5_5252_0[1]); 
    wire [1:0] far_5_5253_0;    relay_conn far_5_5253_0_a(.in(layer_4[720]), .out(far_5_5253_0[0]));    relay_conn far_5_5253_0_b(.in(layer_4[631]), .out(far_5_5253_0[1]));
    wire [1:0] far_5_5253_1;    relay_conn far_5_5253_1_a(.in(far_5_5253_0[0]), .out(far_5_5253_1[0]));    relay_conn far_5_5253_1_b(.in(far_5_5253_0[1]), .out(far_5_5253_1[1]));
    assign layer_5[153] = far_5_5253_1[1] & ~far_5_5253_1[0]; 
    assign layer_5[154] = layer_4[880] ^ layer_4[900]; 
    wire [1:0] far_5_5255_0;    relay_conn far_5_5255_0_a(.in(layer_4[554]), .out(far_5_5255_0[0]));    relay_conn far_5_5255_0_b(.in(layer_4[443]), .out(far_5_5255_0[1]));
    wire [1:0] far_5_5255_1;    relay_conn far_5_5255_1_a(.in(far_5_5255_0[0]), .out(far_5_5255_1[0]));    relay_conn far_5_5255_1_b(.in(far_5_5255_0[1]), .out(far_5_5255_1[1]));
    wire [1:0] far_5_5255_2;    relay_conn far_5_5255_2_a(.in(far_5_5255_1[0]), .out(far_5_5255_2[0]));    relay_conn far_5_5255_2_b(.in(far_5_5255_1[1]), .out(far_5_5255_2[1]));
    assign layer_5[155] = far_5_5255_2[0] & ~far_5_5255_2[1]; 
    wire [1:0] far_5_5256_0;    relay_conn far_5_5256_0_a(.in(layer_4[89]), .out(far_5_5256_0[0]));    relay_conn far_5_5256_0_b(.in(layer_4[199]), .out(far_5_5256_0[1]));
    wire [1:0] far_5_5256_1;    relay_conn far_5_5256_1_a(.in(far_5_5256_0[0]), .out(far_5_5256_1[0]));    relay_conn far_5_5256_1_b(.in(far_5_5256_0[1]), .out(far_5_5256_1[1]));
    wire [1:0] far_5_5256_2;    relay_conn far_5_5256_2_a(.in(far_5_5256_1[0]), .out(far_5_5256_2[0]));    relay_conn far_5_5256_2_b(.in(far_5_5256_1[1]), .out(far_5_5256_2[1]));
    assign layer_5[156] = ~far_5_5256_2[0]; 
    wire [1:0] far_5_5257_0;    relay_conn far_5_5257_0_a(.in(layer_4[813]), .out(far_5_5257_0[0]));    relay_conn far_5_5257_0_b(.in(layer_4[852]), .out(far_5_5257_0[1]));
    assign layer_5[157] = far_5_5257_0[1] & ~far_5_5257_0[0]; 
    wire [1:0] far_5_5258_0;    relay_conn far_5_5258_0_a(.in(layer_4[945]), .out(far_5_5258_0[0]));    relay_conn far_5_5258_0_b(.in(layer_4[1000]), .out(far_5_5258_0[1]));
    assign layer_5[158] = ~(far_5_5258_0[0] ^ far_5_5258_0[1]); 
    assign layer_5[159] = ~(layer_4[463] | layer_4[442]); 
    assign layer_5[160] = layer_4[381] & layer_4[377]; 
    assign layer_5[161] = ~layer_4[392]; 
    assign layer_5[162] = layer_4[180] ^ layer_4[168]; 
    assign layer_5[163] = layer_4[628]; 
    assign layer_5[164] = ~layer_4[836]; 
    wire [1:0] far_5_5265_0;    relay_conn far_5_5265_0_a(.in(layer_4[709]), .out(far_5_5265_0[0]));    relay_conn far_5_5265_0_b(.in(layer_4[625]), .out(far_5_5265_0[1]));
    wire [1:0] far_5_5265_1;    relay_conn far_5_5265_1_a(.in(far_5_5265_0[0]), .out(far_5_5265_1[0]));    relay_conn far_5_5265_1_b(.in(far_5_5265_0[1]), .out(far_5_5265_1[1]));
    assign layer_5[165] = far_5_5265_1[0] | far_5_5265_1[1]; 
    wire [1:0] far_5_5266_0;    relay_conn far_5_5266_0_a(.in(layer_4[870]), .out(far_5_5266_0[0]));    relay_conn far_5_5266_0_b(.in(layer_4[830]), .out(far_5_5266_0[1]));
    assign layer_5[166] = ~far_5_5266_0[0]; 
    wire [1:0] far_5_5267_0;    relay_conn far_5_5267_0_a(.in(layer_4[368]), .out(far_5_5267_0[0]));    relay_conn far_5_5267_0_b(.in(layer_4[274]), .out(far_5_5267_0[1]));
    wire [1:0] far_5_5267_1;    relay_conn far_5_5267_1_a(.in(far_5_5267_0[0]), .out(far_5_5267_1[0]));    relay_conn far_5_5267_1_b(.in(far_5_5267_0[1]), .out(far_5_5267_1[1]));
    assign layer_5[167] = far_5_5267_1[1] & ~far_5_5267_1[0]; 
    wire [1:0] far_5_5268_0;    relay_conn far_5_5268_0_a(.in(layer_4[526]), .out(far_5_5268_0[0]));    relay_conn far_5_5268_0_b(.in(layer_4[645]), .out(far_5_5268_0[1]));
    wire [1:0] far_5_5268_1;    relay_conn far_5_5268_1_a(.in(far_5_5268_0[0]), .out(far_5_5268_1[0]));    relay_conn far_5_5268_1_b(.in(far_5_5268_0[1]), .out(far_5_5268_1[1]));
    wire [1:0] far_5_5268_2;    relay_conn far_5_5268_2_a(.in(far_5_5268_1[0]), .out(far_5_5268_2[0]));    relay_conn far_5_5268_2_b(.in(far_5_5268_1[1]), .out(far_5_5268_2[1]));
    assign layer_5[168] = ~far_5_5268_2[0]; 
    wire [1:0] far_5_5269_0;    relay_conn far_5_5269_0_a(.in(layer_4[693]), .out(far_5_5269_0[0]));    relay_conn far_5_5269_0_b(.in(layer_4[804]), .out(far_5_5269_0[1]));
    wire [1:0] far_5_5269_1;    relay_conn far_5_5269_1_a(.in(far_5_5269_0[0]), .out(far_5_5269_1[0]));    relay_conn far_5_5269_1_b(.in(far_5_5269_0[1]), .out(far_5_5269_1[1]));
    wire [1:0] far_5_5269_2;    relay_conn far_5_5269_2_a(.in(far_5_5269_1[0]), .out(far_5_5269_2[0]));    relay_conn far_5_5269_2_b(.in(far_5_5269_1[1]), .out(far_5_5269_2[1]));
    assign layer_5[169] = far_5_5269_2[0] | far_5_5269_2[1]; 
    assign layer_5[170] = ~(layer_4[309] | layer_4[325]); 
    wire [1:0] far_5_5271_0;    relay_conn far_5_5271_0_a(.in(layer_4[650]), .out(far_5_5271_0[0]));    relay_conn far_5_5271_0_b(.in(layer_4[599]), .out(far_5_5271_0[1]));
    assign layer_5[171] = far_5_5271_0[0] | far_5_5271_0[1]; 
    wire [1:0] far_5_5272_0;    relay_conn far_5_5272_0_a(.in(layer_4[224]), .out(far_5_5272_0[0]));    relay_conn far_5_5272_0_b(.in(layer_4[149]), .out(far_5_5272_0[1]));
    wire [1:0] far_5_5272_1;    relay_conn far_5_5272_1_a(.in(far_5_5272_0[0]), .out(far_5_5272_1[0]));    relay_conn far_5_5272_1_b(.in(far_5_5272_0[1]), .out(far_5_5272_1[1]));
    assign layer_5[172] = far_5_5272_1[0] | far_5_5272_1[1]; 
    wire [1:0] far_5_5273_0;    relay_conn far_5_5273_0_a(.in(layer_4[474]), .out(far_5_5273_0[0]));    relay_conn far_5_5273_0_b(.in(layer_4[401]), .out(far_5_5273_0[1]));
    wire [1:0] far_5_5273_1;    relay_conn far_5_5273_1_a(.in(far_5_5273_0[0]), .out(far_5_5273_1[0]));    relay_conn far_5_5273_1_b(.in(far_5_5273_0[1]), .out(far_5_5273_1[1]));
    assign layer_5[173] = far_5_5273_1[0] & ~far_5_5273_1[1]; 
    assign layer_5[174] = layer_4[930]; 
    wire [1:0] far_5_5275_0;    relay_conn far_5_5275_0_a(.in(layer_4[401]), .out(far_5_5275_0[0]));    relay_conn far_5_5275_0_b(.in(layer_4[509]), .out(far_5_5275_0[1]));
    wire [1:0] far_5_5275_1;    relay_conn far_5_5275_1_a(.in(far_5_5275_0[0]), .out(far_5_5275_1[0]));    relay_conn far_5_5275_1_b(.in(far_5_5275_0[1]), .out(far_5_5275_1[1]));
    wire [1:0] far_5_5275_2;    relay_conn far_5_5275_2_a(.in(far_5_5275_1[0]), .out(far_5_5275_2[0]));    relay_conn far_5_5275_2_b(.in(far_5_5275_1[1]), .out(far_5_5275_2[1]));
    assign layer_5[175] = ~far_5_5275_2[0]; 
    wire [1:0] far_5_5276_0;    relay_conn far_5_5276_0_a(.in(layer_4[608]), .out(far_5_5276_0[0]));    relay_conn far_5_5276_0_b(.in(layer_4[482]), .out(far_5_5276_0[1]));
    wire [1:0] far_5_5276_1;    relay_conn far_5_5276_1_a(.in(far_5_5276_0[0]), .out(far_5_5276_1[0]));    relay_conn far_5_5276_1_b(.in(far_5_5276_0[1]), .out(far_5_5276_1[1]));
    wire [1:0] far_5_5276_2;    relay_conn far_5_5276_2_a(.in(far_5_5276_1[0]), .out(far_5_5276_2[0]));    relay_conn far_5_5276_2_b(.in(far_5_5276_1[1]), .out(far_5_5276_2[1]));
    assign layer_5[176] = far_5_5276_2[0]; 
    wire [1:0] far_5_5277_0;    relay_conn far_5_5277_0_a(.in(layer_4[109]), .out(far_5_5277_0[0]));    relay_conn far_5_5277_0_b(.in(layer_4[23]), .out(far_5_5277_0[1]));
    wire [1:0] far_5_5277_1;    relay_conn far_5_5277_1_a(.in(far_5_5277_0[0]), .out(far_5_5277_1[0]));    relay_conn far_5_5277_1_b(.in(far_5_5277_0[1]), .out(far_5_5277_1[1]));
    assign layer_5[177] = ~(far_5_5277_1[0] & far_5_5277_1[1]); 
    wire [1:0] far_5_5278_0;    relay_conn far_5_5278_0_a(.in(layer_4[884]), .out(far_5_5278_0[0]));    relay_conn far_5_5278_0_b(.in(layer_4[852]), .out(far_5_5278_0[1]));
    assign layer_5[178] = ~far_5_5278_0[0] | (far_5_5278_0[0] & far_5_5278_0[1]); 
    wire [1:0] far_5_5279_0;    relay_conn far_5_5279_0_a(.in(layer_4[952]), .out(far_5_5279_0[0]));    relay_conn far_5_5279_0_b(.in(layer_4[862]), .out(far_5_5279_0[1]));
    wire [1:0] far_5_5279_1;    relay_conn far_5_5279_1_a(.in(far_5_5279_0[0]), .out(far_5_5279_1[0]));    relay_conn far_5_5279_1_b(.in(far_5_5279_0[1]), .out(far_5_5279_1[1]));
    assign layer_5[179] = far_5_5279_1[1]; 
    wire [1:0] far_5_5280_0;    relay_conn far_5_5280_0_a(.in(layer_4[630]), .out(far_5_5280_0[0]));    relay_conn far_5_5280_0_b(.in(layer_4[516]), .out(far_5_5280_0[1]));
    wire [1:0] far_5_5280_1;    relay_conn far_5_5280_1_a(.in(far_5_5280_0[0]), .out(far_5_5280_1[0]));    relay_conn far_5_5280_1_b(.in(far_5_5280_0[1]), .out(far_5_5280_1[1]));
    wire [1:0] far_5_5280_2;    relay_conn far_5_5280_2_a(.in(far_5_5280_1[0]), .out(far_5_5280_2[0]));    relay_conn far_5_5280_2_b(.in(far_5_5280_1[1]), .out(far_5_5280_2[1]));
    assign layer_5[180] = far_5_5280_2[1]; 
    assign layer_5[181] = layer_4[527] ^ layer_4[534]; 
    wire [1:0] far_5_5282_0;    relay_conn far_5_5282_0_a(.in(layer_4[995]), .out(far_5_5282_0[0]));    relay_conn far_5_5282_0_b(.in(layer_4[899]), .out(far_5_5282_0[1]));
    wire [1:0] far_5_5282_1;    relay_conn far_5_5282_1_a(.in(far_5_5282_0[0]), .out(far_5_5282_1[0]));    relay_conn far_5_5282_1_b(.in(far_5_5282_0[1]), .out(far_5_5282_1[1]));
    wire [1:0] far_5_5282_2;    relay_conn far_5_5282_2_a(.in(far_5_5282_1[0]), .out(far_5_5282_2[0]));    relay_conn far_5_5282_2_b(.in(far_5_5282_1[1]), .out(far_5_5282_2[1]));
    assign layer_5[182] = far_5_5282_2[0]; 
    assign layer_5[183] = ~layer_4[728]; 
    wire [1:0] far_5_5284_0;    relay_conn far_5_5284_0_a(.in(layer_4[536]), .out(far_5_5284_0[0]));    relay_conn far_5_5284_0_b(.in(layer_4[594]), .out(far_5_5284_0[1]));
    assign layer_5[184] = ~far_5_5284_0[0]; 
    wire [1:0] far_5_5285_0;    relay_conn far_5_5285_0_a(.in(layer_4[80]), .out(far_5_5285_0[0]));    relay_conn far_5_5285_0_b(.in(layer_4[45]), .out(far_5_5285_0[1]));
    assign layer_5[185] = ~far_5_5285_0[1] | (far_5_5285_0[0] & far_5_5285_0[1]); 
    wire [1:0] far_5_5286_0;    relay_conn far_5_5286_0_a(.in(layer_4[913]), .out(far_5_5286_0[0]));    relay_conn far_5_5286_0_b(.in(layer_4[997]), .out(far_5_5286_0[1]));
    wire [1:0] far_5_5286_1;    relay_conn far_5_5286_1_a(.in(far_5_5286_0[0]), .out(far_5_5286_1[0]));    relay_conn far_5_5286_1_b(.in(far_5_5286_0[1]), .out(far_5_5286_1[1]));
    assign layer_5[186] = ~far_5_5286_1[0] | (far_5_5286_1[0] & far_5_5286_1[1]); 
    wire [1:0] far_5_5287_0;    relay_conn far_5_5287_0_a(.in(layer_4[542]), .out(far_5_5287_0[0]));    relay_conn far_5_5287_0_b(.in(layer_4[614]), .out(far_5_5287_0[1]));
    wire [1:0] far_5_5287_1;    relay_conn far_5_5287_1_a(.in(far_5_5287_0[0]), .out(far_5_5287_1[0]));    relay_conn far_5_5287_1_b(.in(far_5_5287_0[1]), .out(far_5_5287_1[1]));
    assign layer_5[187] = far_5_5287_1[0] & ~far_5_5287_1[1]; 
    wire [1:0] far_5_5288_0;    relay_conn far_5_5288_0_a(.in(layer_4[502]), .out(far_5_5288_0[0]));    relay_conn far_5_5288_0_b(.in(layer_4[551]), .out(far_5_5288_0[1]));
    assign layer_5[188] = ~(far_5_5288_0[0] ^ far_5_5288_0[1]); 
    wire [1:0] far_5_5289_0;    relay_conn far_5_5289_0_a(.in(layer_4[232]), .out(far_5_5289_0[0]));    relay_conn far_5_5289_0_b(.in(layer_4[172]), .out(far_5_5289_0[1]));
    assign layer_5[189] = ~far_5_5289_0[0] | (far_5_5289_0[0] & far_5_5289_0[1]); 
    wire [1:0] far_5_5290_0;    relay_conn far_5_5290_0_a(.in(layer_4[612]), .out(far_5_5290_0[0]));    relay_conn far_5_5290_0_b(.in(layer_4[720]), .out(far_5_5290_0[1]));
    wire [1:0] far_5_5290_1;    relay_conn far_5_5290_1_a(.in(far_5_5290_0[0]), .out(far_5_5290_1[0]));    relay_conn far_5_5290_1_b(.in(far_5_5290_0[1]), .out(far_5_5290_1[1]));
    wire [1:0] far_5_5290_2;    relay_conn far_5_5290_2_a(.in(far_5_5290_1[0]), .out(far_5_5290_2[0]));    relay_conn far_5_5290_2_b(.in(far_5_5290_1[1]), .out(far_5_5290_2[1]));
    assign layer_5[190] = ~far_5_5290_2[0] | (far_5_5290_2[0] & far_5_5290_2[1]); 
    wire [1:0] far_5_5291_0;    relay_conn far_5_5291_0_a(.in(layer_4[419]), .out(far_5_5291_0[0]));    relay_conn far_5_5291_0_b(.in(layer_4[330]), .out(far_5_5291_0[1]));
    wire [1:0] far_5_5291_1;    relay_conn far_5_5291_1_a(.in(far_5_5291_0[0]), .out(far_5_5291_1[0]));    relay_conn far_5_5291_1_b(.in(far_5_5291_0[1]), .out(far_5_5291_1[1]));
    assign layer_5[191] = ~far_5_5291_1[1]; 
    wire [1:0] far_5_5292_0;    relay_conn far_5_5292_0_a(.in(layer_4[741]), .out(far_5_5292_0[0]));    relay_conn far_5_5292_0_b(.in(layer_4[709]), .out(far_5_5292_0[1]));
    assign layer_5[192] = ~(far_5_5292_0[0] ^ far_5_5292_0[1]); 
    assign layer_5[193] = layer_4[794] ^ layer_4[806]; 
    assign layer_5[194] = ~layer_4[443] | (layer_4[443] & layer_4[424]); 
    wire [1:0] far_5_5295_0;    relay_conn far_5_5295_0_a(.in(layer_4[417]), .out(far_5_5295_0[0]));    relay_conn far_5_5295_0_b(.in(layer_4[385]), .out(far_5_5295_0[1]));
    assign layer_5[195] = far_5_5295_0[0] & ~far_5_5295_0[1]; 
    wire [1:0] far_5_5296_0;    relay_conn far_5_5296_0_a(.in(layer_4[297]), .out(far_5_5296_0[0]));    relay_conn far_5_5296_0_b(.in(layer_4[185]), .out(far_5_5296_0[1]));
    wire [1:0] far_5_5296_1;    relay_conn far_5_5296_1_a(.in(far_5_5296_0[0]), .out(far_5_5296_1[0]));    relay_conn far_5_5296_1_b(.in(far_5_5296_0[1]), .out(far_5_5296_1[1]));
    wire [1:0] far_5_5296_2;    relay_conn far_5_5296_2_a(.in(far_5_5296_1[0]), .out(far_5_5296_2[0]));    relay_conn far_5_5296_2_b(.in(far_5_5296_1[1]), .out(far_5_5296_2[1]));
    assign layer_5[196] = ~(far_5_5296_2[0] & far_5_5296_2[1]); 
    wire [1:0] far_5_5297_0;    relay_conn far_5_5297_0_a(.in(layer_4[508]), .out(far_5_5297_0[0]));    relay_conn far_5_5297_0_b(.in(layer_4[580]), .out(far_5_5297_0[1]));
    wire [1:0] far_5_5297_1;    relay_conn far_5_5297_1_a(.in(far_5_5297_0[0]), .out(far_5_5297_1[0]));    relay_conn far_5_5297_1_b(.in(far_5_5297_0[1]), .out(far_5_5297_1[1]));
    assign layer_5[197] = far_5_5297_1[0] | far_5_5297_1[1]; 
    wire [1:0] far_5_5298_0;    relay_conn far_5_5298_0_a(.in(layer_4[369]), .out(far_5_5298_0[0]));    relay_conn far_5_5298_0_b(.in(layer_4[409]), .out(far_5_5298_0[1]));
    assign layer_5[198] = ~(far_5_5298_0[0] & far_5_5298_0[1]); 
    wire [1:0] far_5_5299_0;    relay_conn far_5_5299_0_a(.in(layer_4[149]), .out(far_5_5299_0[0]));    relay_conn far_5_5299_0_b(.in(layer_4[250]), .out(far_5_5299_0[1]));
    wire [1:0] far_5_5299_1;    relay_conn far_5_5299_1_a(.in(far_5_5299_0[0]), .out(far_5_5299_1[0]));    relay_conn far_5_5299_1_b(.in(far_5_5299_0[1]), .out(far_5_5299_1[1]));
    wire [1:0] far_5_5299_2;    relay_conn far_5_5299_2_a(.in(far_5_5299_1[0]), .out(far_5_5299_2[0]));    relay_conn far_5_5299_2_b(.in(far_5_5299_1[1]), .out(far_5_5299_2[1]));
    assign layer_5[199] = ~(far_5_5299_2[0] & far_5_5299_2[1]); 
    wire [1:0] far_5_5300_0;    relay_conn far_5_5300_0_a(.in(layer_4[1017]), .out(far_5_5300_0[0]));    relay_conn far_5_5300_0_b(.in(layer_4[959]), .out(far_5_5300_0[1]));
    assign layer_5[200] = ~(far_5_5300_0[0] & far_5_5300_0[1]); 
    wire [1:0] far_5_5301_0;    relay_conn far_5_5301_0_a(.in(layer_4[224]), .out(far_5_5301_0[0]));    relay_conn far_5_5301_0_b(.in(layer_4[294]), .out(far_5_5301_0[1]));
    wire [1:0] far_5_5301_1;    relay_conn far_5_5301_1_a(.in(far_5_5301_0[0]), .out(far_5_5301_1[0]));    relay_conn far_5_5301_1_b(.in(far_5_5301_0[1]), .out(far_5_5301_1[1]));
    assign layer_5[201] = far_5_5301_1[0] & far_5_5301_1[1]; 
    wire [1:0] far_5_5302_0;    relay_conn far_5_5302_0_a(.in(layer_4[730]), .out(far_5_5302_0[0]));    relay_conn far_5_5302_0_b(.in(layer_4[602]), .out(far_5_5302_0[1]));
    wire [1:0] far_5_5302_1;    relay_conn far_5_5302_1_a(.in(far_5_5302_0[0]), .out(far_5_5302_1[0]));    relay_conn far_5_5302_1_b(.in(far_5_5302_0[1]), .out(far_5_5302_1[1]));
    wire [1:0] far_5_5302_2;    relay_conn far_5_5302_2_a(.in(far_5_5302_1[0]), .out(far_5_5302_2[0]));    relay_conn far_5_5302_2_b(.in(far_5_5302_1[1]), .out(far_5_5302_2[1]));
    wire [1:0] far_5_5302_3;    relay_conn far_5_5302_3_a(.in(far_5_5302_2[0]), .out(far_5_5302_3[0]));    relay_conn far_5_5302_3_b(.in(far_5_5302_2[1]), .out(far_5_5302_3[1]));
    assign layer_5[202] = ~far_5_5302_3[1] | (far_5_5302_3[0] & far_5_5302_3[1]); 
    wire [1:0] far_5_5303_0;    relay_conn far_5_5303_0_a(.in(layer_4[1019]), .out(far_5_5303_0[0]));    relay_conn far_5_5303_0_b(.in(layer_4[941]), .out(far_5_5303_0[1]));
    wire [1:0] far_5_5303_1;    relay_conn far_5_5303_1_a(.in(far_5_5303_0[0]), .out(far_5_5303_1[0]));    relay_conn far_5_5303_1_b(.in(far_5_5303_0[1]), .out(far_5_5303_1[1]));
    assign layer_5[203] = far_5_5303_1[0] & ~far_5_5303_1[1]; 
    assign layer_5[204] = layer_4[350] | layer_4[324]; 
    wire [1:0] far_5_5305_0;    relay_conn far_5_5305_0_a(.in(layer_4[654]), .out(far_5_5305_0[0]));    relay_conn far_5_5305_0_b(.in(layer_4[716]), .out(far_5_5305_0[1]));
    assign layer_5[205] = ~far_5_5305_0[1]; 
    assign layer_5[206] = layer_4[854] & ~layer_4[882]; 
    wire [1:0] far_5_5307_0;    relay_conn far_5_5307_0_a(.in(layer_4[397]), .out(far_5_5307_0[0]));    relay_conn far_5_5307_0_b(.in(layer_4[277]), .out(far_5_5307_0[1]));
    wire [1:0] far_5_5307_1;    relay_conn far_5_5307_1_a(.in(far_5_5307_0[0]), .out(far_5_5307_1[0]));    relay_conn far_5_5307_1_b(.in(far_5_5307_0[1]), .out(far_5_5307_1[1]));
    wire [1:0] far_5_5307_2;    relay_conn far_5_5307_2_a(.in(far_5_5307_1[0]), .out(far_5_5307_2[0]));    relay_conn far_5_5307_2_b(.in(far_5_5307_1[1]), .out(far_5_5307_2[1]));
    assign layer_5[207] = far_5_5307_2[1] & ~far_5_5307_2[0]; 
    wire [1:0] far_5_5308_0;    relay_conn far_5_5308_0_a(.in(layer_4[186]), .out(far_5_5308_0[0]));    relay_conn far_5_5308_0_b(.in(layer_4[150]), .out(far_5_5308_0[1]));
    assign layer_5[208] = ~far_5_5308_0[1]; 
    assign layer_5[209] = ~(layer_4[773] | layer_4[799]); 
    wire [1:0] far_5_5310_0;    relay_conn far_5_5310_0_a(.in(layer_4[102]), .out(far_5_5310_0[0]));    relay_conn far_5_5310_0_b(.in(layer_4[189]), .out(far_5_5310_0[1]));
    wire [1:0] far_5_5310_1;    relay_conn far_5_5310_1_a(.in(far_5_5310_0[0]), .out(far_5_5310_1[0]));    relay_conn far_5_5310_1_b(.in(far_5_5310_0[1]), .out(far_5_5310_1[1]));
    assign layer_5[210] = ~far_5_5310_1[0]; 
    wire [1:0] far_5_5311_0;    relay_conn far_5_5311_0_a(.in(layer_4[147]), .out(far_5_5311_0[0]));    relay_conn far_5_5311_0_b(.in(layer_4[215]), .out(far_5_5311_0[1]));
    wire [1:0] far_5_5311_1;    relay_conn far_5_5311_1_a(.in(far_5_5311_0[0]), .out(far_5_5311_1[0]));    relay_conn far_5_5311_1_b(.in(far_5_5311_0[1]), .out(far_5_5311_1[1]));
    assign layer_5[211] = ~far_5_5311_1[0]; 
    wire [1:0] far_5_5312_0;    relay_conn far_5_5312_0_a(.in(layer_4[953]), .out(far_5_5312_0[0]));    relay_conn far_5_5312_0_b(.in(layer_4[1013]), .out(far_5_5312_0[1]));
    assign layer_5[212] = ~far_5_5312_0[0]; 
    wire [1:0] far_5_5313_0;    relay_conn far_5_5313_0_a(.in(layer_4[719]), .out(far_5_5313_0[0]));    relay_conn far_5_5313_0_b(.in(layer_4[806]), .out(far_5_5313_0[1]));
    wire [1:0] far_5_5313_1;    relay_conn far_5_5313_1_a(.in(far_5_5313_0[0]), .out(far_5_5313_1[0]));    relay_conn far_5_5313_1_b(.in(far_5_5313_0[1]), .out(far_5_5313_1[1]));
    assign layer_5[213] = ~far_5_5313_1[1]; 
    assign layer_5[214] = layer_4[12] | layer_4[16]; 
    wire [1:0] far_5_5315_0;    relay_conn far_5_5315_0_a(.in(layer_4[955]), .out(far_5_5315_0[0]));    relay_conn far_5_5315_0_b(.in(layer_4[1018]), .out(far_5_5315_0[1]));
    assign layer_5[215] = far_5_5315_0[0] | far_5_5315_0[1]; 
    wire [1:0] far_5_5316_0;    relay_conn far_5_5316_0_a(.in(layer_4[865]), .out(far_5_5316_0[0]));    relay_conn far_5_5316_0_b(.in(layer_4[818]), .out(far_5_5316_0[1]));
    assign layer_5[216] = far_5_5316_0[0]; 
    wire [1:0] far_5_5317_0;    relay_conn far_5_5317_0_a(.in(layer_4[409]), .out(far_5_5317_0[0]));    relay_conn far_5_5317_0_b(.in(layer_4[287]), .out(far_5_5317_0[1]));
    wire [1:0] far_5_5317_1;    relay_conn far_5_5317_1_a(.in(far_5_5317_0[0]), .out(far_5_5317_1[0]));    relay_conn far_5_5317_1_b(.in(far_5_5317_0[1]), .out(far_5_5317_1[1]));
    wire [1:0] far_5_5317_2;    relay_conn far_5_5317_2_a(.in(far_5_5317_1[0]), .out(far_5_5317_2[0]));    relay_conn far_5_5317_2_b(.in(far_5_5317_1[1]), .out(far_5_5317_2[1]));
    assign layer_5[217] = far_5_5317_2[1]; 
    wire [1:0] far_5_5318_0;    relay_conn far_5_5318_0_a(.in(layer_4[964]), .out(far_5_5318_0[0]));    relay_conn far_5_5318_0_b(.in(layer_4[887]), .out(far_5_5318_0[1]));
    wire [1:0] far_5_5318_1;    relay_conn far_5_5318_1_a(.in(far_5_5318_0[0]), .out(far_5_5318_1[0]));    relay_conn far_5_5318_1_b(.in(far_5_5318_0[1]), .out(far_5_5318_1[1]));
    assign layer_5[218] = far_5_5318_1[0]; 
    wire [1:0] far_5_5319_0;    relay_conn far_5_5319_0_a(.in(layer_4[357]), .out(far_5_5319_0[0]));    relay_conn far_5_5319_0_b(.in(layer_4[299]), .out(far_5_5319_0[1]));
    assign layer_5[219] = ~far_5_5319_0[0]; 
    wire [1:0] far_5_5320_0;    relay_conn far_5_5320_0_a(.in(layer_4[819]), .out(far_5_5320_0[0]));    relay_conn far_5_5320_0_b(.in(layer_4[707]), .out(far_5_5320_0[1]));
    wire [1:0] far_5_5320_1;    relay_conn far_5_5320_1_a(.in(far_5_5320_0[0]), .out(far_5_5320_1[0]));    relay_conn far_5_5320_1_b(.in(far_5_5320_0[1]), .out(far_5_5320_1[1]));
    wire [1:0] far_5_5320_2;    relay_conn far_5_5320_2_a(.in(far_5_5320_1[0]), .out(far_5_5320_2[0]));    relay_conn far_5_5320_2_b(.in(far_5_5320_1[1]), .out(far_5_5320_2[1]));
    assign layer_5[220] = far_5_5320_2[0] | far_5_5320_2[1]; 
    assign layer_5[221] = ~layer_4[397] | (layer_4[397] & layer_4[369]); 
    assign layer_5[222] = ~(layer_4[9] | layer_4[20]); 
    assign layer_5[223] = ~(layer_4[795] ^ layer_4[790]); 
    wire [1:0] far_5_5324_0;    relay_conn far_5_5324_0_a(.in(layer_4[597]), .out(far_5_5324_0[0]));    relay_conn far_5_5324_0_b(.in(layer_4[713]), .out(far_5_5324_0[1]));
    wire [1:0] far_5_5324_1;    relay_conn far_5_5324_1_a(.in(far_5_5324_0[0]), .out(far_5_5324_1[0]));    relay_conn far_5_5324_1_b(.in(far_5_5324_0[1]), .out(far_5_5324_1[1]));
    wire [1:0] far_5_5324_2;    relay_conn far_5_5324_2_a(.in(far_5_5324_1[0]), .out(far_5_5324_2[0]));    relay_conn far_5_5324_2_b(.in(far_5_5324_1[1]), .out(far_5_5324_2[1]));
    assign layer_5[224] = far_5_5324_2[0] & far_5_5324_2[1]; 
    wire [1:0] far_5_5325_0;    relay_conn far_5_5325_0_a(.in(layer_4[969]), .out(far_5_5325_0[0]));    relay_conn far_5_5325_0_b(.in(layer_4[1013]), .out(far_5_5325_0[1]));
    assign layer_5[225] = far_5_5325_0[1]; 
    wire [1:0] far_5_5326_0;    relay_conn far_5_5326_0_a(.in(layer_4[785]), .out(far_5_5326_0[0]));    relay_conn far_5_5326_0_b(.in(layer_4[893]), .out(far_5_5326_0[1]));
    wire [1:0] far_5_5326_1;    relay_conn far_5_5326_1_a(.in(far_5_5326_0[0]), .out(far_5_5326_1[0]));    relay_conn far_5_5326_1_b(.in(far_5_5326_0[1]), .out(far_5_5326_1[1]));
    wire [1:0] far_5_5326_2;    relay_conn far_5_5326_2_a(.in(far_5_5326_1[0]), .out(far_5_5326_2[0]));    relay_conn far_5_5326_2_b(.in(far_5_5326_1[1]), .out(far_5_5326_2[1]));
    assign layer_5[226] = ~far_5_5326_2[0]; 
    wire [1:0] far_5_5327_0;    relay_conn far_5_5327_0_a(.in(layer_4[819]), .out(far_5_5327_0[0]));    relay_conn far_5_5327_0_b(.in(layer_4[941]), .out(far_5_5327_0[1]));
    wire [1:0] far_5_5327_1;    relay_conn far_5_5327_1_a(.in(far_5_5327_0[0]), .out(far_5_5327_1[0]));    relay_conn far_5_5327_1_b(.in(far_5_5327_0[1]), .out(far_5_5327_1[1]));
    wire [1:0] far_5_5327_2;    relay_conn far_5_5327_2_a(.in(far_5_5327_1[0]), .out(far_5_5327_2[0]));    relay_conn far_5_5327_2_b(.in(far_5_5327_1[1]), .out(far_5_5327_2[1]));
    assign layer_5[227] = ~far_5_5327_2[1] | (far_5_5327_2[0] & far_5_5327_2[1]); 
    wire [1:0] far_5_5328_0;    relay_conn far_5_5328_0_a(.in(layer_4[636]), .out(far_5_5328_0[0]));    relay_conn far_5_5328_0_b(.in(layer_4[684]), .out(far_5_5328_0[1]));
    assign layer_5[228] = ~far_5_5328_0[1] | (far_5_5328_0[0] & far_5_5328_0[1]); 
    wire [1:0] far_5_5329_0;    relay_conn far_5_5329_0_a(.in(layer_4[355]), .out(far_5_5329_0[0]));    relay_conn far_5_5329_0_b(.in(layer_4[242]), .out(far_5_5329_0[1]));
    wire [1:0] far_5_5329_1;    relay_conn far_5_5329_1_a(.in(far_5_5329_0[0]), .out(far_5_5329_1[0]));    relay_conn far_5_5329_1_b(.in(far_5_5329_0[1]), .out(far_5_5329_1[1]));
    wire [1:0] far_5_5329_2;    relay_conn far_5_5329_2_a(.in(far_5_5329_1[0]), .out(far_5_5329_2[0]));    relay_conn far_5_5329_2_b(.in(far_5_5329_1[1]), .out(far_5_5329_2[1]));
    assign layer_5[229] = far_5_5329_2[0] & ~far_5_5329_2[1]; 
    wire [1:0] far_5_5330_0;    relay_conn far_5_5330_0_a(.in(layer_4[583]), .out(far_5_5330_0[0]));    relay_conn far_5_5330_0_b(.in(layer_4[644]), .out(far_5_5330_0[1]));
    assign layer_5[230] = ~far_5_5330_0[0] | (far_5_5330_0[0] & far_5_5330_0[1]); 
    assign layer_5[231] = ~layer_4[610]; 
    wire [1:0] far_5_5332_0;    relay_conn far_5_5332_0_a(.in(layer_4[662]), .out(far_5_5332_0[0]));    relay_conn far_5_5332_0_b(.in(layer_4[723]), .out(far_5_5332_0[1]));
    assign layer_5[232] = ~far_5_5332_0[1] | (far_5_5332_0[0] & far_5_5332_0[1]); 
    assign layer_5[233] = ~layer_4[228] | (layer_4[228] & layer_4[210]); 
    wire [1:0] far_5_5334_0;    relay_conn far_5_5334_0_a(.in(layer_4[632]), .out(far_5_5334_0[0]));    relay_conn far_5_5334_0_b(.in(layer_4[598]), .out(far_5_5334_0[1]));
    assign layer_5[234] = ~far_5_5334_0[0]; 
    assign layer_5[235] = ~layer_4[299]; 
    wire [1:0] far_5_5336_0;    relay_conn far_5_5336_0_a(.in(layer_4[135]), .out(far_5_5336_0[0]));    relay_conn far_5_5336_0_b(.in(layer_4[232]), .out(far_5_5336_0[1]));
    wire [1:0] far_5_5336_1;    relay_conn far_5_5336_1_a(.in(far_5_5336_0[0]), .out(far_5_5336_1[0]));    relay_conn far_5_5336_1_b(.in(far_5_5336_0[1]), .out(far_5_5336_1[1]));
    wire [1:0] far_5_5336_2;    relay_conn far_5_5336_2_a(.in(far_5_5336_1[0]), .out(far_5_5336_2[0]));    relay_conn far_5_5336_2_b(.in(far_5_5336_1[1]), .out(far_5_5336_2[1]));
    assign layer_5[236] = ~(far_5_5336_2[0] & far_5_5336_2[1]); 
    assign layer_5[237] = ~(layer_4[999] ^ layer_4[983]); 
    wire [1:0] far_5_5338_0;    relay_conn far_5_5338_0_a(.in(layer_4[565]), .out(far_5_5338_0[0]));    relay_conn far_5_5338_0_b(.in(layer_4[474]), .out(far_5_5338_0[1]));
    wire [1:0] far_5_5338_1;    relay_conn far_5_5338_1_a(.in(far_5_5338_0[0]), .out(far_5_5338_1[0]));    relay_conn far_5_5338_1_b(.in(far_5_5338_0[1]), .out(far_5_5338_1[1]));
    assign layer_5[238] = far_5_5338_1[0] & far_5_5338_1[1]; 
    wire [1:0] far_5_5339_0;    relay_conn far_5_5339_0_a(.in(layer_4[104]), .out(far_5_5339_0[0]));    relay_conn far_5_5339_0_b(.in(layer_4[49]), .out(far_5_5339_0[1]));
    assign layer_5[239] = ~(far_5_5339_0[0] & far_5_5339_0[1]); 
    wire [1:0] far_5_5340_0;    relay_conn far_5_5340_0_a(.in(layer_4[364]), .out(far_5_5340_0[0]));    relay_conn far_5_5340_0_b(.in(layer_4[293]), .out(far_5_5340_0[1]));
    wire [1:0] far_5_5340_1;    relay_conn far_5_5340_1_a(.in(far_5_5340_0[0]), .out(far_5_5340_1[0]));    relay_conn far_5_5340_1_b(.in(far_5_5340_0[1]), .out(far_5_5340_1[1]));
    assign layer_5[240] = far_5_5340_1[0] | far_5_5340_1[1]; 
    wire [1:0] far_5_5341_0;    relay_conn far_5_5341_0_a(.in(layer_4[858]), .out(far_5_5341_0[0]));    relay_conn far_5_5341_0_b(.in(layer_4[822]), .out(far_5_5341_0[1]));
    assign layer_5[241] = far_5_5341_0[0] & far_5_5341_0[1]; 
    wire [1:0] far_5_5342_0;    relay_conn far_5_5342_0_a(.in(layer_4[1002]), .out(far_5_5342_0[0]));    relay_conn far_5_5342_0_b(.in(layer_4[922]), .out(far_5_5342_0[1]));
    wire [1:0] far_5_5342_1;    relay_conn far_5_5342_1_a(.in(far_5_5342_0[0]), .out(far_5_5342_1[0]));    relay_conn far_5_5342_1_b(.in(far_5_5342_0[1]), .out(far_5_5342_1[1]));
    assign layer_5[242] = ~(far_5_5342_1[0] & far_5_5342_1[1]); 
    wire [1:0] far_5_5343_0;    relay_conn far_5_5343_0_a(.in(layer_4[287]), .out(far_5_5343_0[0]));    relay_conn far_5_5343_0_b(.in(layer_4[359]), .out(far_5_5343_0[1]));
    wire [1:0] far_5_5343_1;    relay_conn far_5_5343_1_a(.in(far_5_5343_0[0]), .out(far_5_5343_1[0]));    relay_conn far_5_5343_1_b(.in(far_5_5343_0[1]), .out(far_5_5343_1[1]));
    assign layer_5[243] = far_5_5343_1[1]; 
    wire [1:0] far_5_5344_0;    relay_conn far_5_5344_0_a(.in(layer_4[735]), .out(far_5_5344_0[0]));    relay_conn far_5_5344_0_b(.in(layer_4[848]), .out(far_5_5344_0[1]));
    wire [1:0] far_5_5344_1;    relay_conn far_5_5344_1_a(.in(far_5_5344_0[0]), .out(far_5_5344_1[0]));    relay_conn far_5_5344_1_b(.in(far_5_5344_0[1]), .out(far_5_5344_1[1]));
    wire [1:0] far_5_5344_2;    relay_conn far_5_5344_2_a(.in(far_5_5344_1[0]), .out(far_5_5344_2[0]));    relay_conn far_5_5344_2_b(.in(far_5_5344_1[1]), .out(far_5_5344_2[1]));
    assign layer_5[244] = ~far_5_5344_2[1] | (far_5_5344_2[0] & far_5_5344_2[1]); 
    wire [1:0] far_5_5345_0;    relay_conn far_5_5345_0_a(.in(layer_4[678]), .out(far_5_5345_0[0]));    relay_conn far_5_5345_0_b(.in(layer_4[795]), .out(far_5_5345_0[1]));
    wire [1:0] far_5_5345_1;    relay_conn far_5_5345_1_a(.in(far_5_5345_0[0]), .out(far_5_5345_1[0]));    relay_conn far_5_5345_1_b(.in(far_5_5345_0[1]), .out(far_5_5345_1[1]));
    wire [1:0] far_5_5345_2;    relay_conn far_5_5345_2_a(.in(far_5_5345_1[0]), .out(far_5_5345_2[0]));    relay_conn far_5_5345_2_b(.in(far_5_5345_1[1]), .out(far_5_5345_2[1]));
    assign layer_5[245] = ~(far_5_5345_2[0] | far_5_5345_2[1]); 
    wire [1:0] far_5_5346_0;    relay_conn far_5_5346_0_a(.in(layer_4[215]), .out(far_5_5346_0[0]));    relay_conn far_5_5346_0_b(.in(layer_4[171]), .out(far_5_5346_0[1]));
    assign layer_5[246] = ~far_5_5346_0[1] | (far_5_5346_0[0] & far_5_5346_0[1]); 
    wire [1:0] far_5_5347_0;    relay_conn far_5_5347_0_a(.in(layer_4[258]), .out(far_5_5347_0[0]));    relay_conn far_5_5347_0_b(.in(layer_4[307]), .out(far_5_5347_0[1]));
    assign layer_5[247] = far_5_5347_0[0]; 
    wire [1:0] far_5_5348_0;    relay_conn far_5_5348_0_a(.in(layer_4[436]), .out(far_5_5348_0[0]));    relay_conn far_5_5348_0_b(.in(layer_4[511]), .out(far_5_5348_0[1]));
    wire [1:0] far_5_5348_1;    relay_conn far_5_5348_1_a(.in(far_5_5348_0[0]), .out(far_5_5348_1[0]));    relay_conn far_5_5348_1_b(.in(far_5_5348_0[1]), .out(far_5_5348_1[1]));
    assign layer_5[248] = far_5_5348_1[1]; 
    wire [1:0] far_5_5349_0;    relay_conn far_5_5349_0_a(.in(layer_4[287]), .out(far_5_5349_0[0]));    relay_conn far_5_5349_0_b(.in(layer_4[378]), .out(far_5_5349_0[1]));
    wire [1:0] far_5_5349_1;    relay_conn far_5_5349_1_a(.in(far_5_5349_0[0]), .out(far_5_5349_1[0]));    relay_conn far_5_5349_1_b(.in(far_5_5349_0[1]), .out(far_5_5349_1[1]));
    assign layer_5[249] = ~(far_5_5349_1[0] | far_5_5349_1[1]); 
    wire [1:0] far_5_5350_0;    relay_conn far_5_5350_0_a(.in(layer_4[860]), .out(far_5_5350_0[0]));    relay_conn far_5_5350_0_b(.in(layer_4[774]), .out(far_5_5350_0[1]));
    wire [1:0] far_5_5350_1;    relay_conn far_5_5350_1_a(.in(far_5_5350_0[0]), .out(far_5_5350_1[0]));    relay_conn far_5_5350_1_b(.in(far_5_5350_0[1]), .out(far_5_5350_1[1]));
    assign layer_5[250] = ~(far_5_5350_1[0] & far_5_5350_1[1]); 
    wire [1:0] far_5_5351_0;    relay_conn far_5_5351_0_a(.in(layer_4[588]), .out(far_5_5351_0[0]));    relay_conn far_5_5351_0_b(.in(layer_4[650]), .out(far_5_5351_0[1]));
    assign layer_5[251] = far_5_5351_0[0]; 
    assign layer_5[252] = layer_4[455] & ~layer_4[464]; 
    wire [1:0] far_5_5353_0;    relay_conn far_5_5353_0_a(.in(layer_4[505]), .out(far_5_5353_0[0]));    relay_conn far_5_5353_0_b(.in(layer_4[417]), .out(far_5_5353_0[1]));
    wire [1:0] far_5_5353_1;    relay_conn far_5_5353_1_a(.in(far_5_5353_0[0]), .out(far_5_5353_1[0]));    relay_conn far_5_5353_1_b(.in(far_5_5353_0[1]), .out(far_5_5353_1[1]));
    assign layer_5[253] = far_5_5353_1[0] | far_5_5353_1[1]; 
    assign layer_5[254] = layer_4[66]; 
    assign layer_5[255] = ~(layer_4[899] | layer_4[886]); 
    wire [1:0] far_5_5356_0;    relay_conn far_5_5356_0_a(.in(layer_4[600]), .out(far_5_5356_0[0]));    relay_conn far_5_5356_0_b(.in(layer_4[499]), .out(far_5_5356_0[1]));
    wire [1:0] far_5_5356_1;    relay_conn far_5_5356_1_a(.in(far_5_5356_0[0]), .out(far_5_5356_1[0]));    relay_conn far_5_5356_1_b(.in(far_5_5356_0[1]), .out(far_5_5356_1[1]));
    wire [1:0] far_5_5356_2;    relay_conn far_5_5356_2_a(.in(far_5_5356_1[0]), .out(far_5_5356_2[0]));    relay_conn far_5_5356_2_b(.in(far_5_5356_1[1]), .out(far_5_5356_2[1]));
    assign layer_5[256] = far_5_5356_2[0] | far_5_5356_2[1]; 
    wire [1:0] far_5_5357_0;    relay_conn far_5_5357_0_a(.in(layer_4[541]), .out(far_5_5357_0[0]));    relay_conn far_5_5357_0_b(.in(layer_4[586]), .out(far_5_5357_0[1]));
    assign layer_5[257] = far_5_5357_0[0] | far_5_5357_0[1]; 
    wire [1:0] far_5_5358_0;    relay_conn far_5_5358_0_a(.in(layer_4[518]), .out(far_5_5358_0[0]));    relay_conn far_5_5358_0_b(.in(layer_4[408]), .out(far_5_5358_0[1]));
    wire [1:0] far_5_5358_1;    relay_conn far_5_5358_1_a(.in(far_5_5358_0[0]), .out(far_5_5358_1[0]));    relay_conn far_5_5358_1_b(.in(far_5_5358_0[1]), .out(far_5_5358_1[1]));
    wire [1:0] far_5_5358_2;    relay_conn far_5_5358_2_a(.in(far_5_5358_1[0]), .out(far_5_5358_2[0]));    relay_conn far_5_5358_2_b(.in(far_5_5358_1[1]), .out(far_5_5358_2[1]));
    assign layer_5[258] = ~far_5_5358_2[1]; 
    wire [1:0] far_5_5359_0;    relay_conn far_5_5359_0_a(.in(layer_4[692]), .out(far_5_5359_0[0]));    relay_conn far_5_5359_0_b(.in(layer_4[735]), .out(far_5_5359_0[1]));
    assign layer_5[259] = ~far_5_5359_0[1] | (far_5_5359_0[0] & far_5_5359_0[1]); 
    wire [1:0] far_5_5360_0;    relay_conn far_5_5360_0_a(.in(layer_4[967]), .out(far_5_5360_0[0]));    relay_conn far_5_5360_0_b(.in(layer_4[870]), .out(far_5_5360_0[1]));
    wire [1:0] far_5_5360_1;    relay_conn far_5_5360_1_a(.in(far_5_5360_0[0]), .out(far_5_5360_1[0]));    relay_conn far_5_5360_1_b(.in(far_5_5360_0[1]), .out(far_5_5360_1[1]));
    wire [1:0] far_5_5360_2;    relay_conn far_5_5360_2_a(.in(far_5_5360_1[0]), .out(far_5_5360_2[0]));    relay_conn far_5_5360_2_b(.in(far_5_5360_1[1]), .out(far_5_5360_2[1]));
    assign layer_5[260] = far_5_5360_2[0] & ~far_5_5360_2[1]; 
    wire [1:0] far_5_5361_0;    relay_conn far_5_5361_0_a(.in(layer_4[905]), .out(far_5_5361_0[0]));    relay_conn far_5_5361_0_b(.in(layer_4[938]), .out(far_5_5361_0[1]));
    assign layer_5[261] = ~far_5_5361_0[0]; 
    wire [1:0] far_5_5362_0;    relay_conn far_5_5362_0_a(.in(layer_4[423]), .out(far_5_5362_0[0]));    relay_conn far_5_5362_0_b(.in(layer_4[528]), .out(far_5_5362_0[1]));
    wire [1:0] far_5_5362_1;    relay_conn far_5_5362_1_a(.in(far_5_5362_0[0]), .out(far_5_5362_1[0]));    relay_conn far_5_5362_1_b(.in(far_5_5362_0[1]), .out(far_5_5362_1[1]));
    wire [1:0] far_5_5362_2;    relay_conn far_5_5362_2_a(.in(far_5_5362_1[0]), .out(far_5_5362_2[0]));    relay_conn far_5_5362_2_b(.in(far_5_5362_1[1]), .out(far_5_5362_2[1]));
    assign layer_5[262] = ~(far_5_5362_2[0] | far_5_5362_2[1]); 
    wire [1:0] far_5_5363_0;    relay_conn far_5_5363_0_a(.in(layer_4[109]), .out(far_5_5363_0[0]));    relay_conn far_5_5363_0_b(.in(layer_4[215]), .out(far_5_5363_0[1]));
    wire [1:0] far_5_5363_1;    relay_conn far_5_5363_1_a(.in(far_5_5363_0[0]), .out(far_5_5363_1[0]));    relay_conn far_5_5363_1_b(.in(far_5_5363_0[1]), .out(far_5_5363_1[1]));
    wire [1:0] far_5_5363_2;    relay_conn far_5_5363_2_a(.in(far_5_5363_1[0]), .out(far_5_5363_2[0]));    relay_conn far_5_5363_2_b(.in(far_5_5363_1[1]), .out(far_5_5363_2[1]));
    assign layer_5[263] = far_5_5363_2[1]; 
    wire [1:0] far_5_5364_0;    relay_conn far_5_5364_0_a(.in(layer_4[819]), .out(far_5_5364_0[0]));    relay_conn far_5_5364_0_b(.in(layer_4[898]), .out(far_5_5364_0[1]));
    wire [1:0] far_5_5364_1;    relay_conn far_5_5364_1_a(.in(far_5_5364_0[0]), .out(far_5_5364_1[0]));    relay_conn far_5_5364_1_b(.in(far_5_5364_0[1]), .out(far_5_5364_1[1]));
    assign layer_5[264] = ~(far_5_5364_1[0] ^ far_5_5364_1[1]); 
    wire [1:0] far_5_5365_0;    relay_conn far_5_5365_0_a(.in(layer_4[191]), .out(far_5_5365_0[0]));    relay_conn far_5_5365_0_b(.in(layer_4[158]), .out(far_5_5365_0[1]));
    assign layer_5[265] = far_5_5365_0[1] & ~far_5_5365_0[0]; 
    assign layer_5[266] = ~(layer_4[859] | layer_4[850]); 
    assign layer_5[267] = ~layer_4[301] | (layer_4[309] & layer_4[301]); 
    wire [1:0] far_5_5368_0;    relay_conn far_5_5368_0_a(.in(layer_4[277]), .out(far_5_5368_0[0]));    relay_conn far_5_5368_0_b(.in(layer_4[180]), .out(far_5_5368_0[1]));
    wire [1:0] far_5_5368_1;    relay_conn far_5_5368_1_a(.in(far_5_5368_0[0]), .out(far_5_5368_1[0]));    relay_conn far_5_5368_1_b(.in(far_5_5368_0[1]), .out(far_5_5368_1[1]));
    wire [1:0] far_5_5368_2;    relay_conn far_5_5368_2_a(.in(far_5_5368_1[0]), .out(far_5_5368_2[0]));    relay_conn far_5_5368_2_b(.in(far_5_5368_1[1]), .out(far_5_5368_2[1]));
    assign layer_5[268] = ~(far_5_5368_2[0] & far_5_5368_2[1]); 
    assign layer_5[269] = layer_4[654]; 
    wire [1:0] far_5_5370_0;    relay_conn far_5_5370_0_a(.in(layer_4[158]), .out(far_5_5370_0[0]));    relay_conn far_5_5370_0_b(.in(layer_4[210]), .out(far_5_5370_0[1]));
    assign layer_5[270] = ~(far_5_5370_0[0] | far_5_5370_0[1]); 
    wire [1:0] far_5_5371_0;    relay_conn far_5_5371_0_a(.in(layer_4[4]), .out(far_5_5371_0[0]));    relay_conn far_5_5371_0_b(.in(layer_4[99]), .out(far_5_5371_0[1]));
    wire [1:0] far_5_5371_1;    relay_conn far_5_5371_1_a(.in(far_5_5371_0[0]), .out(far_5_5371_1[0]));    relay_conn far_5_5371_1_b(.in(far_5_5371_0[1]), .out(far_5_5371_1[1]));
    assign layer_5[271] = far_5_5371_1[0] & ~far_5_5371_1[1]; 
    wire [1:0] far_5_5372_0;    relay_conn far_5_5372_0_a(.in(layer_4[421]), .out(far_5_5372_0[0]));    relay_conn far_5_5372_0_b(.in(layer_4[302]), .out(far_5_5372_0[1]));
    wire [1:0] far_5_5372_1;    relay_conn far_5_5372_1_a(.in(far_5_5372_0[0]), .out(far_5_5372_1[0]));    relay_conn far_5_5372_1_b(.in(far_5_5372_0[1]), .out(far_5_5372_1[1]));
    wire [1:0] far_5_5372_2;    relay_conn far_5_5372_2_a(.in(far_5_5372_1[0]), .out(far_5_5372_2[0]));    relay_conn far_5_5372_2_b(.in(far_5_5372_1[1]), .out(far_5_5372_2[1]));
    assign layer_5[272] = far_5_5372_2[0] & far_5_5372_2[1]; 
    wire [1:0] far_5_5373_0;    relay_conn far_5_5373_0_a(.in(layer_4[792]), .out(far_5_5373_0[0]));    relay_conn far_5_5373_0_b(.in(layer_4[735]), .out(far_5_5373_0[1]));
    assign layer_5[273] = ~far_5_5373_0[0]; 
    assign layer_5[274] = layer_4[387] & layer_4[379]; 
    wire [1:0] far_5_5375_0;    relay_conn far_5_5375_0_a(.in(layer_4[56]), .out(far_5_5375_0[0]));    relay_conn far_5_5375_0_b(.in(layer_4[167]), .out(far_5_5375_0[1]));
    wire [1:0] far_5_5375_1;    relay_conn far_5_5375_1_a(.in(far_5_5375_0[0]), .out(far_5_5375_1[0]));    relay_conn far_5_5375_1_b(.in(far_5_5375_0[1]), .out(far_5_5375_1[1]));
    wire [1:0] far_5_5375_2;    relay_conn far_5_5375_2_a(.in(far_5_5375_1[0]), .out(far_5_5375_2[0]));    relay_conn far_5_5375_2_b(.in(far_5_5375_1[1]), .out(far_5_5375_2[1]));
    assign layer_5[275] = ~far_5_5375_2[0] | (far_5_5375_2[0] & far_5_5375_2[1]); 
    wire [1:0] far_5_5376_0;    relay_conn far_5_5376_0_a(.in(layer_4[258]), .out(far_5_5376_0[0]));    relay_conn far_5_5376_0_b(.in(layer_4[358]), .out(far_5_5376_0[1]));
    wire [1:0] far_5_5376_1;    relay_conn far_5_5376_1_a(.in(far_5_5376_0[0]), .out(far_5_5376_1[0]));    relay_conn far_5_5376_1_b(.in(far_5_5376_0[1]), .out(far_5_5376_1[1]));
    wire [1:0] far_5_5376_2;    relay_conn far_5_5376_2_a(.in(far_5_5376_1[0]), .out(far_5_5376_2[0]));    relay_conn far_5_5376_2_b(.in(far_5_5376_1[1]), .out(far_5_5376_2[1]));
    assign layer_5[276] = far_5_5376_2[0]; 
    wire [1:0] far_5_5377_0;    relay_conn far_5_5377_0_a(.in(layer_4[773]), .out(far_5_5377_0[0]));    relay_conn far_5_5377_0_b(.in(layer_4[657]), .out(far_5_5377_0[1]));
    wire [1:0] far_5_5377_1;    relay_conn far_5_5377_1_a(.in(far_5_5377_0[0]), .out(far_5_5377_1[0]));    relay_conn far_5_5377_1_b(.in(far_5_5377_0[1]), .out(far_5_5377_1[1]));
    wire [1:0] far_5_5377_2;    relay_conn far_5_5377_2_a(.in(far_5_5377_1[0]), .out(far_5_5377_2[0]));    relay_conn far_5_5377_2_b(.in(far_5_5377_1[1]), .out(far_5_5377_2[1]));
    assign layer_5[277] = ~far_5_5377_2[0] | (far_5_5377_2[0] & far_5_5377_2[1]); 
    wire [1:0] far_5_5378_0;    relay_conn far_5_5378_0_a(.in(layer_4[936]), .out(far_5_5378_0[0]));    relay_conn far_5_5378_0_b(.in(layer_4[999]), .out(far_5_5378_0[1]));
    assign layer_5[278] = ~far_5_5378_0[1] | (far_5_5378_0[0] & far_5_5378_0[1]); 
    assign layer_5[279] = layer_4[99]; 
    wire [1:0] far_5_5380_0;    relay_conn far_5_5380_0_a(.in(layer_4[867]), .out(far_5_5380_0[0]));    relay_conn far_5_5380_0_b(.in(layer_4[796]), .out(far_5_5380_0[1]));
    wire [1:0] far_5_5380_1;    relay_conn far_5_5380_1_a(.in(far_5_5380_0[0]), .out(far_5_5380_1[0]));    relay_conn far_5_5380_1_b(.in(far_5_5380_0[1]), .out(far_5_5380_1[1]));
    assign layer_5[280] = ~far_5_5380_1[1]; 
    assign layer_5[281] = ~layer_4[867] | (layer_4[867] & layer_4[839]); 
    assign layer_5[282] = layer_4[200]; 
    wire [1:0] far_5_5383_0;    relay_conn far_5_5383_0_a(.in(layer_4[296]), .out(far_5_5383_0[0]));    relay_conn far_5_5383_0_b(.in(layer_4[357]), .out(far_5_5383_0[1]));
    assign layer_5[283] = far_5_5383_0[1]; 
    wire [1:0] far_5_5384_0;    relay_conn far_5_5384_0_a(.in(layer_4[767]), .out(far_5_5384_0[0]));    relay_conn far_5_5384_0_b(.in(layer_4[674]), .out(far_5_5384_0[1]));
    wire [1:0] far_5_5384_1;    relay_conn far_5_5384_1_a(.in(far_5_5384_0[0]), .out(far_5_5384_1[0]));    relay_conn far_5_5384_1_b(.in(far_5_5384_0[1]), .out(far_5_5384_1[1]));
    assign layer_5[284] = ~(far_5_5384_1[0] | far_5_5384_1[1]); 
    wire [1:0] far_5_5385_0;    relay_conn far_5_5385_0_a(.in(layer_4[42]), .out(far_5_5385_0[0]));    relay_conn far_5_5385_0_b(.in(layer_4[124]), .out(far_5_5385_0[1]));
    wire [1:0] far_5_5385_1;    relay_conn far_5_5385_1_a(.in(far_5_5385_0[0]), .out(far_5_5385_1[0]));    relay_conn far_5_5385_1_b(.in(far_5_5385_0[1]), .out(far_5_5385_1[1]));
    assign layer_5[285] = ~far_5_5385_1[0]; 
    wire [1:0] far_5_5386_0;    relay_conn far_5_5386_0_a(.in(layer_4[718]), .out(far_5_5386_0[0]));    relay_conn far_5_5386_0_b(.in(layer_4[661]), .out(far_5_5386_0[1]));
    assign layer_5[286] = ~far_5_5386_0[1] | (far_5_5386_0[0] & far_5_5386_0[1]); 
    wire [1:0] far_5_5387_0;    relay_conn far_5_5387_0_a(.in(layer_4[253]), .out(far_5_5387_0[0]));    relay_conn far_5_5387_0_b(.in(layer_4[131]), .out(far_5_5387_0[1]));
    wire [1:0] far_5_5387_1;    relay_conn far_5_5387_1_a(.in(far_5_5387_0[0]), .out(far_5_5387_1[0]));    relay_conn far_5_5387_1_b(.in(far_5_5387_0[1]), .out(far_5_5387_1[1]));
    wire [1:0] far_5_5387_2;    relay_conn far_5_5387_2_a(.in(far_5_5387_1[0]), .out(far_5_5387_2[0]));    relay_conn far_5_5387_2_b(.in(far_5_5387_1[1]), .out(far_5_5387_2[1]));
    assign layer_5[287] = ~(far_5_5387_2[0] & far_5_5387_2[1]); 
    wire [1:0] far_5_5388_0;    relay_conn far_5_5388_0_a(.in(layer_4[974]), .out(far_5_5388_0[0]));    relay_conn far_5_5388_0_b(.in(layer_4[1015]), .out(far_5_5388_0[1]));
    assign layer_5[288] = far_5_5388_0[0] & far_5_5388_0[1]; 
    wire [1:0] far_5_5389_0;    relay_conn far_5_5389_0_a(.in(layer_4[760]), .out(far_5_5389_0[0]));    relay_conn far_5_5389_0_b(.in(layer_4[886]), .out(far_5_5389_0[1]));
    wire [1:0] far_5_5389_1;    relay_conn far_5_5389_1_a(.in(far_5_5389_0[0]), .out(far_5_5389_1[0]));    relay_conn far_5_5389_1_b(.in(far_5_5389_0[1]), .out(far_5_5389_1[1]));
    wire [1:0] far_5_5389_2;    relay_conn far_5_5389_2_a(.in(far_5_5389_1[0]), .out(far_5_5389_2[0]));    relay_conn far_5_5389_2_b(.in(far_5_5389_1[1]), .out(far_5_5389_2[1]));
    assign layer_5[289] = far_5_5389_2[1]; 
    assign layer_5[290] = layer_4[654] & ~layer_4[636]; 
    assign layer_5[291] = layer_4[186]; 
    wire [1:0] far_5_5392_0;    relay_conn far_5_5392_0_a(.in(layer_4[369]), .out(far_5_5392_0[0]));    relay_conn far_5_5392_0_b(.in(layer_4[245]), .out(far_5_5392_0[1]));
    wire [1:0] far_5_5392_1;    relay_conn far_5_5392_1_a(.in(far_5_5392_0[0]), .out(far_5_5392_1[0]));    relay_conn far_5_5392_1_b(.in(far_5_5392_0[1]), .out(far_5_5392_1[1]));
    wire [1:0] far_5_5392_2;    relay_conn far_5_5392_2_a(.in(far_5_5392_1[0]), .out(far_5_5392_2[0]));    relay_conn far_5_5392_2_b(.in(far_5_5392_1[1]), .out(far_5_5392_2[1]));
    assign layer_5[292] = ~(far_5_5392_2[0] | far_5_5392_2[1]); 
    wire [1:0] far_5_5393_0;    relay_conn far_5_5393_0_a(.in(layer_4[115]), .out(far_5_5393_0[0]));    relay_conn far_5_5393_0_b(.in(layer_4[16]), .out(far_5_5393_0[1]));
    wire [1:0] far_5_5393_1;    relay_conn far_5_5393_1_a(.in(far_5_5393_0[0]), .out(far_5_5393_1[0]));    relay_conn far_5_5393_1_b(.in(far_5_5393_0[1]), .out(far_5_5393_1[1]));
    wire [1:0] far_5_5393_2;    relay_conn far_5_5393_2_a(.in(far_5_5393_1[0]), .out(far_5_5393_2[0]));    relay_conn far_5_5393_2_b(.in(far_5_5393_1[1]), .out(far_5_5393_2[1]));
    assign layer_5[293] = ~far_5_5393_2[1] | (far_5_5393_2[0] & far_5_5393_2[1]); 
    wire [1:0] far_5_5394_0;    relay_conn far_5_5394_0_a(.in(layer_4[743]), .out(far_5_5394_0[0]));    relay_conn far_5_5394_0_b(.in(layer_4[707]), .out(far_5_5394_0[1]));
    assign layer_5[294] = far_5_5394_0[1]; 
    wire [1:0] far_5_5395_0;    relay_conn far_5_5395_0_a(.in(layer_4[495]), .out(far_5_5395_0[0]));    relay_conn far_5_5395_0_b(.in(layer_4[538]), .out(far_5_5395_0[1]));
    assign layer_5[295] = far_5_5395_0[1] & ~far_5_5395_0[0]; 
    assign layer_5[296] = layer_4[18] & ~layer_4[20]; 
    wire [1:0] far_5_5397_0;    relay_conn far_5_5397_0_a(.in(layer_4[477]), .out(far_5_5397_0[0]));    relay_conn far_5_5397_0_b(.in(layer_4[548]), .out(far_5_5397_0[1]));
    wire [1:0] far_5_5397_1;    relay_conn far_5_5397_1_a(.in(far_5_5397_0[0]), .out(far_5_5397_1[0]));    relay_conn far_5_5397_1_b(.in(far_5_5397_0[1]), .out(far_5_5397_1[1]));
    assign layer_5[297] = ~far_5_5397_1[0]; 
    assign layer_5[298] = layer_4[574]; 
    wire [1:0] far_5_5399_0;    relay_conn far_5_5399_0_a(.in(layer_4[217]), .out(far_5_5399_0[0]));    relay_conn far_5_5399_0_b(.in(layer_4[294]), .out(far_5_5399_0[1]));
    wire [1:0] far_5_5399_1;    relay_conn far_5_5399_1_a(.in(far_5_5399_0[0]), .out(far_5_5399_1[0]));    relay_conn far_5_5399_1_b(.in(far_5_5399_0[1]), .out(far_5_5399_1[1]));
    assign layer_5[299] = far_5_5399_1[0] ^ far_5_5399_1[1]; 
    wire [1:0] far_5_5400_0;    relay_conn far_5_5400_0_a(.in(layer_4[279]), .out(far_5_5400_0[0]));    relay_conn far_5_5400_0_b(.in(layer_4[210]), .out(far_5_5400_0[1]));
    wire [1:0] far_5_5400_1;    relay_conn far_5_5400_1_a(.in(far_5_5400_0[0]), .out(far_5_5400_1[0]));    relay_conn far_5_5400_1_b(.in(far_5_5400_0[1]), .out(far_5_5400_1[1]));
    assign layer_5[300] = ~far_5_5400_1[1]; 
    assign layer_5[301] = layer_4[898] & layer_4[916]; 
    wire [1:0] far_5_5402_0;    relay_conn far_5_5402_0_a(.in(layer_4[636]), .out(far_5_5402_0[0]));    relay_conn far_5_5402_0_b(.in(layer_4[719]), .out(far_5_5402_0[1]));
    wire [1:0] far_5_5402_1;    relay_conn far_5_5402_1_a(.in(far_5_5402_0[0]), .out(far_5_5402_1[0]));    relay_conn far_5_5402_1_b(.in(far_5_5402_0[1]), .out(far_5_5402_1[1]));
    assign layer_5[302] = far_5_5402_1[1]; 
    wire [1:0] far_5_5403_0;    relay_conn far_5_5403_0_a(.in(layer_4[896]), .out(far_5_5403_0[0]));    relay_conn far_5_5403_0_b(.in(layer_4[1003]), .out(far_5_5403_0[1]));
    wire [1:0] far_5_5403_1;    relay_conn far_5_5403_1_a(.in(far_5_5403_0[0]), .out(far_5_5403_1[0]));    relay_conn far_5_5403_1_b(.in(far_5_5403_0[1]), .out(far_5_5403_1[1]));
    wire [1:0] far_5_5403_2;    relay_conn far_5_5403_2_a(.in(far_5_5403_1[0]), .out(far_5_5403_2[0]));    relay_conn far_5_5403_2_b(.in(far_5_5403_1[1]), .out(far_5_5403_2[1]));
    assign layer_5[303] = far_5_5403_2[0]; 
    assign layer_5[304] = layer_4[426] & ~layer_4[438]; 
    wire [1:0] far_5_5405_0;    relay_conn far_5_5405_0_a(.in(layer_4[736]), .out(far_5_5405_0[0]));    relay_conn far_5_5405_0_b(.in(layer_4[697]), .out(far_5_5405_0[1]));
    assign layer_5[305] = far_5_5405_0[1]; 
    wire [1:0] far_5_5406_0;    relay_conn far_5_5406_0_a(.in(layer_4[974]), .out(far_5_5406_0[0]));    relay_conn far_5_5406_0_b(.in(layer_4[1008]), .out(far_5_5406_0[1]));
    assign layer_5[306] = far_5_5406_0[0] & far_5_5406_0[1]; 
    wire [1:0] far_5_5407_0;    relay_conn far_5_5407_0_a(.in(layer_4[969]), .out(far_5_5407_0[0]));    relay_conn far_5_5407_0_b(.in(layer_4[905]), .out(far_5_5407_0[1]));
    wire [1:0] far_5_5407_1;    relay_conn far_5_5407_1_a(.in(far_5_5407_0[0]), .out(far_5_5407_1[0]));    relay_conn far_5_5407_1_b(.in(far_5_5407_0[1]), .out(far_5_5407_1[1]));
    assign layer_5[307] = ~far_5_5407_1[0]; 
    wire [1:0] far_5_5408_0;    relay_conn far_5_5408_0_a(.in(layer_4[614]), .out(far_5_5408_0[0]));    relay_conn far_5_5408_0_b(.in(layer_4[581]), .out(far_5_5408_0[1]));
    assign layer_5[308] = far_5_5408_0[0] & ~far_5_5408_0[1]; 
    wire [1:0] far_5_5409_0;    relay_conn far_5_5409_0_a(.in(layer_4[13]), .out(far_5_5409_0[0]));    relay_conn far_5_5409_0_b(.in(layer_4[52]), .out(far_5_5409_0[1]));
    assign layer_5[309] = ~(far_5_5409_0[0] ^ far_5_5409_0[1]); 
    wire [1:0] far_5_5410_0;    relay_conn far_5_5410_0_a(.in(layer_4[224]), .out(far_5_5410_0[0]));    relay_conn far_5_5410_0_b(.in(layer_4[258]), .out(far_5_5410_0[1]));
    assign layer_5[310] = ~far_5_5410_0[0]; 
    wire [1:0] far_5_5411_0;    relay_conn far_5_5411_0_a(.in(layer_4[407]), .out(far_5_5411_0[0]));    relay_conn far_5_5411_0_b(.in(layer_4[365]), .out(far_5_5411_0[1]));
    assign layer_5[311] = ~far_5_5411_0[0] | (far_5_5411_0[0] & far_5_5411_0[1]); 
    assign layer_5[312] = ~layer_4[439]; 
    wire [1:0] far_5_5413_0;    relay_conn far_5_5413_0_a(.in(layer_4[813]), .out(far_5_5413_0[0]));    relay_conn far_5_5413_0_b(.in(layer_4[886]), .out(far_5_5413_0[1]));
    wire [1:0] far_5_5413_1;    relay_conn far_5_5413_1_a(.in(far_5_5413_0[0]), .out(far_5_5413_1[0]));    relay_conn far_5_5413_1_b(.in(far_5_5413_0[1]), .out(far_5_5413_1[1]));
    assign layer_5[313] = ~(far_5_5413_1[0] | far_5_5413_1[1]); 
    wire [1:0] far_5_5414_0;    relay_conn far_5_5414_0_a(.in(layer_4[178]), .out(far_5_5414_0[0]));    relay_conn far_5_5414_0_b(.in(layer_4[134]), .out(far_5_5414_0[1]));
    assign layer_5[314] = ~far_5_5414_0[1]; 
    wire [1:0] far_5_5415_0;    relay_conn far_5_5415_0_a(.in(layer_4[16]), .out(far_5_5415_0[0]));    relay_conn far_5_5415_0_b(.in(layer_4[141]), .out(far_5_5415_0[1]));
    wire [1:0] far_5_5415_1;    relay_conn far_5_5415_1_a(.in(far_5_5415_0[0]), .out(far_5_5415_1[0]));    relay_conn far_5_5415_1_b(.in(far_5_5415_0[1]), .out(far_5_5415_1[1]));
    wire [1:0] far_5_5415_2;    relay_conn far_5_5415_2_a(.in(far_5_5415_1[0]), .out(far_5_5415_2[0]));    relay_conn far_5_5415_2_b(.in(far_5_5415_1[1]), .out(far_5_5415_2[1]));
    assign layer_5[315] = ~far_5_5415_2[0] | (far_5_5415_2[0] & far_5_5415_2[1]); 
    wire [1:0] far_5_5416_0;    relay_conn far_5_5416_0_a(.in(layer_4[632]), .out(far_5_5416_0[0]));    relay_conn far_5_5416_0_b(.in(layer_4[666]), .out(far_5_5416_0[1]));
    assign layer_5[316] = ~far_5_5416_0[1]; 
    wire [1:0] far_5_5417_0;    relay_conn far_5_5417_0_a(.in(layer_4[939]), .out(far_5_5417_0[0]));    relay_conn far_5_5417_0_b(.in(layer_4[1015]), .out(far_5_5417_0[1]));
    wire [1:0] far_5_5417_1;    relay_conn far_5_5417_1_a(.in(far_5_5417_0[0]), .out(far_5_5417_1[0]));    relay_conn far_5_5417_1_b(.in(far_5_5417_0[1]), .out(far_5_5417_1[1]));
    assign layer_5[317] = ~(far_5_5417_1[0] | far_5_5417_1[1]); 
    wire [1:0] far_5_5418_0;    relay_conn far_5_5418_0_a(.in(layer_4[254]), .out(far_5_5418_0[0]));    relay_conn far_5_5418_0_b(.in(layer_4[150]), .out(far_5_5418_0[1]));
    wire [1:0] far_5_5418_1;    relay_conn far_5_5418_1_a(.in(far_5_5418_0[0]), .out(far_5_5418_1[0]));    relay_conn far_5_5418_1_b(.in(far_5_5418_0[1]), .out(far_5_5418_1[1]));
    wire [1:0] far_5_5418_2;    relay_conn far_5_5418_2_a(.in(far_5_5418_1[0]), .out(far_5_5418_2[0]));    relay_conn far_5_5418_2_b(.in(far_5_5418_1[1]), .out(far_5_5418_2[1]));
    assign layer_5[318] = far_5_5418_2[1] & ~far_5_5418_2[0]; 
    wire [1:0] far_5_5419_0;    relay_conn far_5_5419_0_a(.in(layer_4[761]), .out(far_5_5419_0[0]));    relay_conn far_5_5419_0_b(.in(layer_4[707]), .out(far_5_5419_0[1]));
    assign layer_5[319] = ~far_5_5419_0[1] | (far_5_5419_0[0] & far_5_5419_0[1]); 
    wire [1:0] far_5_5420_0;    relay_conn far_5_5420_0_a(.in(layer_4[392]), .out(far_5_5420_0[0]));    relay_conn far_5_5420_0_b(.in(layer_4[443]), .out(far_5_5420_0[1]));
    assign layer_5[320] = ~(far_5_5420_0[0] & far_5_5420_0[1]); 
    wire [1:0] far_5_5421_0;    relay_conn far_5_5421_0_a(.in(layer_4[902]), .out(far_5_5421_0[0]));    relay_conn far_5_5421_0_b(.in(layer_4[991]), .out(far_5_5421_0[1]));
    wire [1:0] far_5_5421_1;    relay_conn far_5_5421_1_a(.in(far_5_5421_0[0]), .out(far_5_5421_1[0]));    relay_conn far_5_5421_1_b(.in(far_5_5421_0[1]), .out(far_5_5421_1[1]));
    assign layer_5[321] = ~far_5_5421_1[1] | (far_5_5421_1[0] & far_5_5421_1[1]); 
    wire [1:0] far_5_5422_0;    relay_conn far_5_5422_0_a(.in(layer_4[666]), .out(far_5_5422_0[0]));    relay_conn far_5_5422_0_b(.in(layer_4[712]), .out(far_5_5422_0[1]));
    assign layer_5[322] = ~far_5_5422_0[0]; 
    wire [1:0] far_5_5423_0;    relay_conn far_5_5423_0_a(.in(layer_4[589]), .out(far_5_5423_0[0]));    relay_conn far_5_5423_0_b(.in(layer_4[636]), .out(far_5_5423_0[1]));
    assign layer_5[323] = ~far_5_5423_0[1]; 
    wire [1:0] far_5_5424_0;    relay_conn far_5_5424_0_a(.in(layer_4[1015]), .out(far_5_5424_0[0]));    relay_conn far_5_5424_0_b(.in(layer_4[959]), .out(far_5_5424_0[1]));
    assign layer_5[324] = far_5_5424_0[1] & ~far_5_5424_0[0]; 
    wire [1:0] far_5_5425_0;    relay_conn far_5_5425_0_a(.in(layer_4[654]), .out(far_5_5425_0[0]));    relay_conn far_5_5425_0_b(.in(layer_4[615]), .out(far_5_5425_0[1]));
    assign layer_5[325] = far_5_5425_0[0] & ~far_5_5425_0[1]; 
    wire [1:0] far_5_5426_0;    relay_conn far_5_5426_0_a(.in(layer_4[530]), .out(far_5_5426_0[0]));    relay_conn far_5_5426_0_b(.in(layer_4[408]), .out(far_5_5426_0[1]));
    wire [1:0] far_5_5426_1;    relay_conn far_5_5426_1_a(.in(far_5_5426_0[0]), .out(far_5_5426_1[0]));    relay_conn far_5_5426_1_b(.in(far_5_5426_0[1]), .out(far_5_5426_1[1]));
    wire [1:0] far_5_5426_2;    relay_conn far_5_5426_2_a(.in(far_5_5426_1[0]), .out(far_5_5426_2[0]));    relay_conn far_5_5426_2_b(.in(far_5_5426_1[1]), .out(far_5_5426_2[1]));
    assign layer_5[326] = far_5_5426_2[0] & far_5_5426_2[1]; 
    wire [1:0] far_5_5427_0;    relay_conn far_5_5427_0_a(.in(layer_4[900]), .out(far_5_5427_0[0]));    relay_conn far_5_5427_0_b(.in(layer_4[980]), .out(far_5_5427_0[1]));
    wire [1:0] far_5_5427_1;    relay_conn far_5_5427_1_a(.in(far_5_5427_0[0]), .out(far_5_5427_1[0]));    relay_conn far_5_5427_1_b(.in(far_5_5427_0[1]), .out(far_5_5427_1[1]));
    assign layer_5[327] = far_5_5427_1[0]; 
    assign layer_5[328] = ~layer_4[936]; 
    assign layer_5[329] = layer_4[168] ^ layer_4[141]; 
    wire [1:0] far_5_5430_0;    relay_conn far_5_5430_0_a(.in(layer_4[164]), .out(far_5_5430_0[0]));    relay_conn far_5_5430_0_b(.in(layer_4[266]), .out(far_5_5430_0[1]));
    wire [1:0] far_5_5430_1;    relay_conn far_5_5430_1_a(.in(far_5_5430_0[0]), .out(far_5_5430_1[0]));    relay_conn far_5_5430_1_b(.in(far_5_5430_0[1]), .out(far_5_5430_1[1]));
    wire [1:0] far_5_5430_2;    relay_conn far_5_5430_2_a(.in(far_5_5430_1[0]), .out(far_5_5430_2[0]));    relay_conn far_5_5430_2_b(.in(far_5_5430_1[1]), .out(far_5_5430_2[1]));
    assign layer_5[330] = ~(far_5_5430_2[0] | far_5_5430_2[1]); 
    wire [1:0] far_5_5431_0;    relay_conn far_5_5431_0_a(.in(layer_4[186]), .out(far_5_5431_0[0]));    relay_conn far_5_5431_0_b(.in(layer_4[138]), .out(far_5_5431_0[1]));
    assign layer_5[331] = far_5_5431_0[0] ^ far_5_5431_0[1]; 
    wire [1:0] far_5_5432_0;    relay_conn far_5_5432_0_a(.in(layer_4[10]), .out(far_5_5432_0[0]));    relay_conn far_5_5432_0_b(.in(layer_4[103]), .out(far_5_5432_0[1]));
    wire [1:0] far_5_5432_1;    relay_conn far_5_5432_1_a(.in(far_5_5432_0[0]), .out(far_5_5432_1[0]));    relay_conn far_5_5432_1_b(.in(far_5_5432_0[1]), .out(far_5_5432_1[1]));
    assign layer_5[332] = ~far_5_5432_1[1]; 
    wire [1:0] far_5_5433_0;    relay_conn far_5_5433_0_a(.in(layer_4[994]), .out(far_5_5433_0[0]));    relay_conn far_5_5433_0_b(.in(layer_4[921]), .out(far_5_5433_0[1]));
    wire [1:0] far_5_5433_1;    relay_conn far_5_5433_1_a(.in(far_5_5433_0[0]), .out(far_5_5433_1[0]));    relay_conn far_5_5433_1_b(.in(far_5_5433_0[1]), .out(far_5_5433_1[1]));
    assign layer_5[333] = ~far_5_5433_1[0]; 
    wire [1:0] far_5_5434_0;    relay_conn far_5_5434_0_a(.in(layer_4[395]), .out(far_5_5434_0[0]));    relay_conn far_5_5434_0_b(.in(layer_4[438]), .out(far_5_5434_0[1]));
    assign layer_5[334] = far_5_5434_0[0] | far_5_5434_0[1]; 
    wire [1:0] far_5_5435_0;    relay_conn far_5_5435_0_a(.in(layer_4[690]), .out(far_5_5435_0[0]));    relay_conn far_5_5435_0_b(.in(layer_4[589]), .out(far_5_5435_0[1]));
    wire [1:0] far_5_5435_1;    relay_conn far_5_5435_1_a(.in(far_5_5435_0[0]), .out(far_5_5435_1[0]));    relay_conn far_5_5435_1_b(.in(far_5_5435_0[1]), .out(far_5_5435_1[1]));
    wire [1:0] far_5_5435_2;    relay_conn far_5_5435_2_a(.in(far_5_5435_1[0]), .out(far_5_5435_2[0]));    relay_conn far_5_5435_2_b(.in(far_5_5435_1[1]), .out(far_5_5435_2[1]));
    assign layer_5[335] = ~far_5_5435_2[1]; 
    wire [1:0] far_5_5436_0;    relay_conn far_5_5436_0_a(.in(layer_4[39]), .out(far_5_5436_0[0]));    relay_conn far_5_5436_0_b(.in(layer_4[147]), .out(far_5_5436_0[1]));
    wire [1:0] far_5_5436_1;    relay_conn far_5_5436_1_a(.in(far_5_5436_0[0]), .out(far_5_5436_1[0]));    relay_conn far_5_5436_1_b(.in(far_5_5436_0[1]), .out(far_5_5436_1[1]));
    wire [1:0] far_5_5436_2;    relay_conn far_5_5436_2_a(.in(far_5_5436_1[0]), .out(far_5_5436_2[0]));    relay_conn far_5_5436_2_b(.in(far_5_5436_1[1]), .out(far_5_5436_2[1]));
    assign layer_5[336] = ~(far_5_5436_2[0] & far_5_5436_2[1]); 
    wire [1:0] far_5_5437_0;    relay_conn far_5_5437_0_a(.in(layer_4[261]), .out(far_5_5437_0[0]));    relay_conn far_5_5437_0_b(.in(layer_4[294]), .out(far_5_5437_0[1]));
    assign layer_5[337] = far_5_5437_0[0]; 
    wire [1:0] far_5_5438_0;    relay_conn far_5_5438_0_a(.in(layer_4[366]), .out(far_5_5438_0[0]));    relay_conn far_5_5438_0_b(.in(layer_4[447]), .out(far_5_5438_0[1]));
    wire [1:0] far_5_5438_1;    relay_conn far_5_5438_1_a(.in(far_5_5438_0[0]), .out(far_5_5438_1[0]));    relay_conn far_5_5438_1_b(.in(far_5_5438_0[1]), .out(far_5_5438_1[1]));
    assign layer_5[338] = ~(far_5_5438_1[0] ^ far_5_5438_1[1]); 
    wire [1:0] far_5_5439_0;    relay_conn far_5_5439_0_a(.in(layer_4[559]), .out(far_5_5439_0[0]));    relay_conn far_5_5439_0_b(.in(layer_4[472]), .out(far_5_5439_0[1]));
    wire [1:0] far_5_5439_1;    relay_conn far_5_5439_1_a(.in(far_5_5439_0[0]), .out(far_5_5439_1[0]));    relay_conn far_5_5439_1_b(.in(far_5_5439_0[1]), .out(far_5_5439_1[1]));
    assign layer_5[339] = far_5_5439_1[0] | far_5_5439_1[1]; 
    assign layer_5[340] = ~layer_4[190]; 
    wire [1:0] far_5_5441_0;    relay_conn far_5_5441_0_a(.in(layer_4[154]), .out(far_5_5441_0[0]));    relay_conn far_5_5441_0_b(.in(layer_4[77]), .out(far_5_5441_0[1]));
    wire [1:0] far_5_5441_1;    relay_conn far_5_5441_1_a(.in(far_5_5441_0[0]), .out(far_5_5441_1[0]));    relay_conn far_5_5441_1_b(.in(far_5_5441_0[1]), .out(far_5_5441_1[1]));
    assign layer_5[341] = far_5_5441_1[1]; 
    assign layer_5[342] = ~(layer_4[397] & layer_4[384]); 
    wire [1:0] far_5_5443_0;    relay_conn far_5_5443_0_a(.in(layer_4[576]), .out(far_5_5443_0[0]));    relay_conn far_5_5443_0_b(.in(layer_4[675]), .out(far_5_5443_0[1]));
    wire [1:0] far_5_5443_1;    relay_conn far_5_5443_1_a(.in(far_5_5443_0[0]), .out(far_5_5443_1[0]));    relay_conn far_5_5443_1_b(.in(far_5_5443_0[1]), .out(far_5_5443_1[1]));
    wire [1:0] far_5_5443_2;    relay_conn far_5_5443_2_a(.in(far_5_5443_1[0]), .out(far_5_5443_2[0]));    relay_conn far_5_5443_2_b(.in(far_5_5443_1[1]), .out(far_5_5443_2[1]));
    assign layer_5[343] = far_5_5443_2[0] & far_5_5443_2[1]; 
    wire [1:0] far_5_5444_0;    relay_conn far_5_5444_0_a(.in(layer_4[192]), .out(far_5_5444_0[0]));    relay_conn far_5_5444_0_b(.in(layer_4[266]), .out(far_5_5444_0[1]));
    wire [1:0] far_5_5444_1;    relay_conn far_5_5444_1_a(.in(far_5_5444_0[0]), .out(far_5_5444_1[0]));    relay_conn far_5_5444_1_b(.in(far_5_5444_0[1]), .out(far_5_5444_1[1]));
    assign layer_5[344] = far_5_5444_1[0] | far_5_5444_1[1]; 
    assign layer_5[345] = layer_4[99] | layer_4[107]; 
    wire [1:0] far_5_5446_0;    relay_conn far_5_5446_0_a(.in(layer_4[910]), .out(far_5_5446_0[0]));    relay_conn far_5_5446_0_b(.in(layer_4[850]), .out(far_5_5446_0[1]));
    assign layer_5[346] = ~far_5_5446_0[1]; 
    assign layer_5[347] = layer_4[650] & ~layer_4[658]; 
    wire [1:0] far_5_5448_0;    relay_conn far_5_5448_0_a(.in(layer_4[656]), .out(far_5_5448_0[0]));    relay_conn far_5_5448_0_b(.in(layer_4[616]), .out(far_5_5448_0[1]));
    assign layer_5[348] = ~(far_5_5448_0[0] & far_5_5448_0[1]); 
    wire [1:0] far_5_5449_0;    relay_conn far_5_5449_0_a(.in(layer_4[590]), .out(far_5_5449_0[0]));    relay_conn far_5_5449_0_b(.in(layer_4[544]), .out(far_5_5449_0[1]));
    assign layer_5[349] = ~far_5_5449_0[0] | (far_5_5449_0[0] & far_5_5449_0[1]); 
    wire [1:0] far_5_5450_0;    relay_conn far_5_5450_0_a(.in(layer_4[201]), .out(far_5_5450_0[0]));    relay_conn far_5_5450_0_b(.in(layer_4[140]), .out(far_5_5450_0[1]));
    assign layer_5[350] = ~far_5_5450_0[1]; 
    wire [1:0] far_5_5451_0;    relay_conn far_5_5451_0_a(.in(layer_4[620]), .out(far_5_5451_0[0]));    relay_conn far_5_5451_0_b(.in(layer_4[528]), .out(far_5_5451_0[1]));
    wire [1:0] far_5_5451_1;    relay_conn far_5_5451_1_a(.in(far_5_5451_0[0]), .out(far_5_5451_1[0]));    relay_conn far_5_5451_1_b(.in(far_5_5451_0[1]), .out(far_5_5451_1[1]));
    assign layer_5[351] = ~far_5_5451_1[0] | (far_5_5451_1[0] & far_5_5451_1[1]); 
    assign layer_5[352] = ~layer_4[1001]; 
    assign layer_5[353] = layer_4[220]; 
    wire [1:0] far_5_5454_0;    relay_conn far_5_5454_0_a(.in(layer_4[417]), .out(far_5_5454_0[0]));    relay_conn far_5_5454_0_b(.in(layer_4[453]), .out(far_5_5454_0[1]));
    assign layer_5[354] = ~(far_5_5454_0[0] ^ far_5_5454_0[1]); 
    wire [1:0] far_5_5455_0;    relay_conn far_5_5455_0_a(.in(layer_4[995]), .out(far_5_5455_0[0]));    relay_conn far_5_5455_0_b(.in(layer_4[905]), .out(far_5_5455_0[1]));
    wire [1:0] far_5_5455_1;    relay_conn far_5_5455_1_a(.in(far_5_5455_0[0]), .out(far_5_5455_1[0]));    relay_conn far_5_5455_1_b(.in(far_5_5455_0[1]), .out(far_5_5455_1[1]));
    assign layer_5[355] = ~(far_5_5455_1[0] | far_5_5455_1[1]); 
    wire [1:0] far_5_5456_0;    relay_conn far_5_5456_0_a(.in(layer_4[498]), .out(far_5_5456_0[0]));    relay_conn far_5_5456_0_b(.in(layer_4[604]), .out(far_5_5456_0[1]));
    wire [1:0] far_5_5456_1;    relay_conn far_5_5456_1_a(.in(far_5_5456_0[0]), .out(far_5_5456_1[0]));    relay_conn far_5_5456_1_b(.in(far_5_5456_0[1]), .out(far_5_5456_1[1]));
    wire [1:0] far_5_5456_2;    relay_conn far_5_5456_2_a(.in(far_5_5456_1[0]), .out(far_5_5456_2[0]));    relay_conn far_5_5456_2_b(.in(far_5_5456_1[1]), .out(far_5_5456_2[1]));
    assign layer_5[356] = far_5_5456_2[0] | far_5_5456_2[1]; 
    wire [1:0] far_5_5457_0;    relay_conn far_5_5457_0_a(.in(layer_4[363]), .out(far_5_5457_0[0]));    relay_conn far_5_5457_0_b(.in(layer_4[271]), .out(far_5_5457_0[1]));
    wire [1:0] far_5_5457_1;    relay_conn far_5_5457_1_a(.in(far_5_5457_0[0]), .out(far_5_5457_1[0]));    relay_conn far_5_5457_1_b(.in(far_5_5457_0[1]), .out(far_5_5457_1[1]));
    assign layer_5[357] = ~far_5_5457_1[1]; 
    assign layer_5[358] = layer_4[12] & ~layer_4[43]; 
    assign layer_5[359] = ~layer_4[202] | (layer_4[228] & layer_4[202]); 
    wire [1:0] far_5_5460_0;    relay_conn far_5_5460_0_a(.in(layer_4[692]), .out(far_5_5460_0[0]));    relay_conn far_5_5460_0_b(.in(layer_4[660]), .out(far_5_5460_0[1]));
    assign layer_5[360] = far_5_5460_0[1]; 
    assign layer_5[361] = layer_4[337]; 
    wire [1:0] far_5_5462_0;    relay_conn far_5_5462_0_a(.in(layer_4[813]), .out(far_5_5462_0[0]));    relay_conn far_5_5462_0_b(.in(layer_4[726]), .out(far_5_5462_0[1]));
    wire [1:0] far_5_5462_1;    relay_conn far_5_5462_1_a(.in(far_5_5462_0[0]), .out(far_5_5462_1[0]));    relay_conn far_5_5462_1_b(.in(far_5_5462_0[1]), .out(far_5_5462_1[1]));
    assign layer_5[362] = far_5_5462_1[1] & ~far_5_5462_1[0]; 
    assign layer_5[363] = layer_4[279] & layer_4[300]; 
    wire [1:0] far_5_5464_0;    relay_conn far_5_5464_0_a(.in(layer_4[227]), .out(far_5_5464_0[0]));    relay_conn far_5_5464_0_b(.in(layer_4[141]), .out(far_5_5464_0[1]));
    wire [1:0] far_5_5464_1;    relay_conn far_5_5464_1_a(.in(far_5_5464_0[0]), .out(far_5_5464_1[0]));    relay_conn far_5_5464_1_b(.in(far_5_5464_0[1]), .out(far_5_5464_1[1]));
    assign layer_5[364] = ~far_5_5464_1[0] | (far_5_5464_1[0] & far_5_5464_1[1]); 
    wire [1:0] far_5_5465_0;    relay_conn far_5_5465_0_a(.in(layer_4[640]), .out(far_5_5465_0[0]));    relay_conn far_5_5465_0_b(.in(layer_4[735]), .out(far_5_5465_0[1]));
    wire [1:0] far_5_5465_1;    relay_conn far_5_5465_1_a(.in(far_5_5465_0[0]), .out(far_5_5465_1[0]));    relay_conn far_5_5465_1_b(.in(far_5_5465_0[1]), .out(far_5_5465_1[1]));
    assign layer_5[365] = ~(far_5_5465_1[0] & far_5_5465_1[1]); 
    wire [1:0] far_5_5466_0;    relay_conn far_5_5466_0_a(.in(layer_4[647]), .out(far_5_5466_0[0]));    relay_conn far_5_5466_0_b(.in(layer_4[584]), .out(far_5_5466_0[1]));
    assign layer_5[366] = ~far_5_5466_0[1]; 
    wire [1:0] far_5_5467_0;    relay_conn far_5_5467_0_a(.in(layer_4[134]), .out(far_5_5467_0[0]));    relay_conn far_5_5467_0_b(.in(layer_4[59]), .out(far_5_5467_0[1]));
    wire [1:0] far_5_5467_1;    relay_conn far_5_5467_1_a(.in(far_5_5467_0[0]), .out(far_5_5467_1[0]));    relay_conn far_5_5467_1_b(.in(far_5_5467_0[1]), .out(far_5_5467_1[1]));
    assign layer_5[367] = far_5_5467_1[0] | far_5_5467_1[1]; 
    wire [1:0] far_5_5468_0;    relay_conn far_5_5468_0_a(.in(layer_4[882]), .out(far_5_5468_0[0]));    relay_conn far_5_5468_0_b(.in(layer_4[830]), .out(far_5_5468_0[1]));
    assign layer_5[368] = ~(far_5_5468_0[0] | far_5_5468_0[1]); 
    assign layer_5[369] = layer_4[986]; 
    assign layer_5[370] = layer_4[709] | layer_4[718]; 
    assign layer_5[371] = layer_4[359] | layer_4[386]; 
    wire [1:0] far_5_5472_0;    relay_conn far_5_5472_0_a(.in(layer_4[269]), .out(far_5_5472_0[0]));    relay_conn far_5_5472_0_b(.in(layer_4[386]), .out(far_5_5472_0[1]));
    wire [1:0] far_5_5472_1;    relay_conn far_5_5472_1_a(.in(far_5_5472_0[0]), .out(far_5_5472_1[0]));    relay_conn far_5_5472_1_b(.in(far_5_5472_0[1]), .out(far_5_5472_1[1]));
    wire [1:0] far_5_5472_2;    relay_conn far_5_5472_2_a(.in(far_5_5472_1[0]), .out(far_5_5472_2[0]));    relay_conn far_5_5472_2_b(.in(far_5_5472_1[1]), .out(far_5_5472_2[1]));
    assign layer_5[372] = ~(far_5_5472_2[0] ^ far_5_5472_2[1]); 
    wire [1:0] far_5_5473_0;    relay_conn far_5_5473_0_a(.in(layer_4[748]), .out(far_5_5473_0[0]));    relay_conn far_5_5473_0_b(.in(layer_4[795]), .out(far_5_5473_0[1]));
    assign layer_5[373] = ~(far_5_5473_0[0] | far_5_5473_0[1]); 
    wire [1:0] far_5_5474_0;    relay_conn far_5_5474_0_a(.in(layer_4[81]), .out(far_5_5474_0[0]));    relay_conn far_5_5474_0_b(.in(layer_4[190]), .out(far_5_5474_0[1]));
    wire [1:0] far_5_5474_1;    relay_conn far_5_5474_1_a(.in(far_5_5474_0[0]), .out(far_5_5474_1[0]));    relay_conn far_5_5474_1_b(.in(far_5_5474_0[1]), .out(far_5_5474_1[1]));
    wire [1:0] far_5_5474_2;    relay_conn far_5_5474_2_a(.in(far_5_5474_1[0]), .out(far_5_5474_2[0]));    relay_conn far_5_5474_2_b(.in(far_5_5474_1[1]), .out(far_5_5474_2[1]));
    assign layer_5[374] = ~far_5_5474_2[1]; 
    wire [1:0] far_5_5475_0;    relay_conn far_5_5475_0_a(.in(layer_4[512]), .out(far_5_5475_0[0]));    relay_conn far_5_5475_0_b(.in(layer_4[638]), .out(far_5_5475_0[1]));
    wire [1:0] far_5_5475_1;    relay_conn far_5_5475_1_a(.in(far_5_5475_0[0]), .out(far_5_5475_1[0]));    relay_conn far_5_5475_1_b(.in(far_5_5475_0[1]), .out(far_5_5475_1[1]));
    wire [1:0] far_5_5475_2;    relay_conn far_5_5475_2_a(.in(far_5_5475_1[0]), .out(far_5_5475_2[0]));    relay_conn far_5_5475_2_b(.in(far_5_5475_1[1]), .out(far_5_5475_2[1]));
    assign layer_5[375] = far_5_5475_2[1] & ~far_5_5475_2[0]; 
    wire [1:0] far_5_5476_0;    relay_conn far_5_5476_0_a(.in(layer_4[1016]), .out(far_5_5476_0[0]));    relay_conn far_5_5476_0_b(.in(layer_4[961]), .out(far_5_5476_0[1]));
    assign layer_5[376] = ~far_5_5476_0[0]; 
    wire [1:0] far_5_5477_0;    relay_conn far_5_5477_0_a(.in(layer_4[103]), .out(far_5_5477_0[0]));    relay_conn far_5_5477_0_b(.in(layer_4[208]), .out(far_5_5477_0[1]));
    wire [1:0] far_5_5477_1;    relay_conn far_5_5477_1_a(.in(far_5_5477_0[0]), .out(far_5_5477_1[0]));    relay_conn far_5_5477_1_b(.in(far_5_5477_0[1]), .out(far_5_5477_1[1]));
    wire [1:0] far_5_5477_2;    relay_conn far_5_5477_2_a(.in(far_5_5477_1[0]), .out(far_5_5477_2[0]));    relay_conn far_5_5477_2_b(.in(far_5_5477_1[1]), .out(far_5_5477_2[1]));
    assign layer_5[377] = far_5_5477_2[0] ^ far_5_5477_2[1]; 
    wire [1:0] far_5_5478_0;    relay_conn far_5_5478_0_a(.in(layer_4[300]), .out(far_5_5478_0[0]));    relay_conn far_5_5478_0_b(.in(layer_4[215]), .out(far_5_5478_0[1]));
    wire [1:0] far_5_5478_1;    relay_conn far_5_5478_1_a(.in(far_5_5478_0[0]), .out(far_5_5478_1[0]));    relay_conn far_5_5478_1_b(.in(far_5_5478_0[1]), .out(far_5_5478_1[1]));
    assign layer_5[378] = ~(far_5_5478_1[0] | far_5_5478_1[1]); 
    wire [1:0] far_5_5479_0;    relay_conn far_5_5479_0_a(.in(layer_4[699]), .out(far_5_5479_0[0]));    relay_conn far_5_5479_0_b(.in(layer_4[636]), .out(far_5_5479_0[1]));
    assign layer_5[379] = far_5_5479_0[0] & ~far_5_5479_0[1]; 
    assign layer_5[380] = layer_4[795] | layer_4[813]; 
    wire [1:0] far_5_5481_0;    relay_conn far_5_5481_0_a(.in(layer_4[886]), .out(far_5_5481_0[0]));    relay_conn far_5_5481_0_b(.in(layer_4[806]), .out(far_5_5481_0[1]));
    wire [1:0] far_5_5481_1;    relay_conn far_5_5481_1_a(.in(far_5_5481_0[0]), .out(far_5_5481_1[0]));    relay_conn far_5_5481_1_b(.in(far_5_5481_0[1]), .out(far_5_5481_1[1]));
    assign layer_5[381] = ~far_5_5481_1[0]; 
    assign layer_5[382] = ~layer_4[831] | (layer_4[813] & layer_4[831]); 
    wire [1:0] far_5_5483_0;    relay_conn far_5_5483_0_a(.in(layer_4[921]), .out(far_5_5483_0[0]));    relay_conn far_5_5483_0_b(.in(layer_4[850]), .out(far_5_5483_0[1]));
    wire [1:0] far_5_5483_1;    relay_conn far_5_5483_1_a(.in(far_5_5483_0[0]), .out(far_5_5483_1[0]));    relay_conn far_5_5483_1_b(.in(far_5_5483_0[1]), .out(far_5_5483_1[1]));
    assign layer_5[383] = ~(far_5_5483_1[0] | far_5_5483_1[1]); 
    wire [1:0] far_5_5484_0;    relay_conn far_5_5484_0_a(.in(layer_4[644]), .out(far_5_5484_0[0]));    relay_conn far_5_5484_0_b(.in(layer_4[752]), .out(far_5_5484_0[1]));
    wire [1:0] far_5_5484_1;    relay_conn far_5_5484_1_a(.in(far_5_5484_0[0]), .out(far_5_5484_1[0]));    relay_conn far_5_5484_1_b(.in(far_5_5484_0[1]), .out(far_5_5484_1[1]));
    wire [1:0] far_5_5484_2;    relay_conn far_5_5484_2_a(.in(far_5_5484_1[0]), .out(far_5_5484_2[0]));    relay_conn far_5_5484_2_b(.in(far_5_5484_1[1]), .out(far_5_5484_2[1]));
    assign layer_5[384] = ~far_5_5484_2[1]; 
    wire [1:0] far_5_5485_0;    relay_conn far_5_5485_0_a(.in(layer_4[208]), .out(far_5_5485_0[0]));    relay_conn far_5_5485_0_b(.in(layer_4[287]), .out(far_5_5485_0[1]));
    wire [1:0] far_5_5485_1;    relay_conn far_5_5485_1_a(.in(far_5_5485_0[0]), .out(far_5_5485_1[0]));    relay_conn far_5_5485_1_b(.in(far_5_5485_0[1]), .out(far_5_5485_1[1]));
    assign layer_5[385] = ~far_5_5485_1[1] | (far_5_5485_1[0] & far_5_5485_1[1]); 
    wire [1:0] far_5_5486_0;    relay_conn far_5_5486_0_a(.in(layer_4[410]), .out(far_5_5486_0[0]));    relay_conn far_5_5486_0_b(.in(layer_4[306]), .out(far_5_5486_0[1]));
    wire [1:0] far_5_5486_1;    relay_conn far_5_5486_1_a(.in(far_5_5486_0[0]), .out(far_5_5486_1[0]));    relay_conn far_5_5486_1_b(.in(far_5_5486_0[1]), .out(far_5_5486_1[1]));
    wire [1:0] far_5_5486_2;    relay_conn far_5_5486_2_a(.in(far_5_5486_1[0]), .out(far_5_5486_2[0]));    relay_conn far_5_5486_2_b(.in(far_5_5486_1[1]), .out(far_5_5486_2[1]));
    assign layer_5[386] = ~far_5_5486_2[0] | (far_5_5486_2[0] & far_5_5486_2[1]); 
    assign layer_5[387] = ~(layer_4[495] ^ layer_4[475]); 
    wire [1:0] far_5_5488_0;    relay_conn far_5_5488_0_a(.in(layer_4[131]), .out(far_5_5488_0[0]));    relay_conn far_5_5488_0_b(.in(layer_4[166]), .out(far_5_5488_0[1]));
    assign layer_5[388] = far_5_5488_0[0] & ~far_5_5488_0[1]; 
    wire [1:0] far_5_5489_0;    relay_conn far_5_5489_0_a(.in(layer_4[974]), .out(far_5_5489_0[0]));    relay_conn far_5_5489_0_b(.in(layer_4[871]), .out(far_5_5489_0[1]));
    wire [1:0] far_5_5489_1;    relay_conn far_5_5489_1_a(.in(far_5_5489_0[0]), .out(far_5_5489_1[0]));    relay_conn far_5_5489_1_b(.in(far_5_5489_0[1]), .out(far_5_5489_1[1]));
    wire [1:0] far_5_5489_2;    relay_conn far_5_5489_2_a(.in(far_5_5489_1[0]), .out(far_5_5489_2[0]));    relay_conn far_5_5489_2_b(.in(far_5_5489_1[1]), .out(far_5_5489_2[1]));
    assign layer_5[389] = ~(far_5_5489_2[0] | far_5_5489_2[1]); 
    wire [1:0] far_5_5490_0;    relay_conn far_5_5490_0_a(.in(layer_4[974]), .out(far_5_5490_0[0]));    relay_conn far_5_5490_0_b(.in(layer_4[898]), .out(far_5_5490_0[1]));
    wire [1:0] far_5_5490_1;    relay_conn far_5_5490_1_a(.in(far_5_5490_0[0]), .out(far_5_5490_1[0]));    relay_conn far_5_5490_1_b(.in(far_5_5490_0[1]), .out(far_5_5490_1[1]));
    assign layer_5[390] = ~(far_5_5490_1[0] & far_5_5490_1[1]); 
    assign layer_5[391] = ~(layer_4[2] | layer_4[27]); 
    wire [1:0] far_5_5492_0;    relay_conn far_5_5492_0_a(.in(layer_4[62]), .out(far_5_5492_0[0]));    relay_conn far_5_5492_0_b(.in(layer_4[139]), .out(far_5_5492_0[1]));
    wire [1:0] far_5_5492_1;    relay_conn far_5_5492_1_a(.in(far_5_5492_0[0]), .out(far_5_5492_1[0]));    relay_conn far_5_5492_1_b(.in(far_5_5492_0[1]), .out(far_5_5492_1[1]));
    assign layer_5[392] = ~(far_5_5492_1[0] & far_5_5492_1[1]); 
    assign layer_5[393] = layer_4[813] & ~layer_4[819]; 
    wire [1:0] far_5_5494_0;    relay_conn far_5_5494_0_a(.in(layer_4[497]), .out(far_5_5494_0[0]));    relay_conn far_5_5494_0_b(.in(layer_4[454]), .out(far_5_5494_0[1]));
    assign layer_5[394] = ~far_5_5494_0[0] | (far_5_5494_0[0] & far_5_5494_0[1]); 
    assign layer_5[395] = ~layer_4[357]; 
    wire [1:0] far_5_5496_0;    relay_conn far_5_5496_0_a(.in(layer_4[642]), .out(far_5_5496_0[0]));    relay_conn far_5_5496_0_b(.in(layer_4[589]), .out(far_5_5496_0[1]));
    assign layer_5[396] = ~far_5_5496_0[1]; 
    wire [1:0] far_5_5497_0;    relay_conn far_5_5497_0_a(.in(layer_4[859]), .out(far_5_5497_0[0]));    relay_conn far_5_5497_0_b(.in(layer_4[754]), .out(far_5_5497_0[1]));
    wire [1:0] far_5_5497_1;    relay_conn far_5_5497_1_a(.in(far_5_5497_0[0]), .out(far_5_5497_1[0]));    relay_conn far_5_5497_1_b(.in(far_5_5497_0[1]), .out(far_5_5497_1[1]));
    wire [1:0] far_5_5497_2;    relay_conn far_5_5497_2_a(.in(far_5_5497_1[0]), .out(far_5_5497_2[0]));    relay_conn far_5_5497_2_b(.in(far_5_5497_1[1]), .out(far_5_5497_2[1]));
    assign layer_5[397] = far_5_5497_2[0] | far_5_5497_2[1]; 
    assign layer_5[398] = layer_4[895]; 
    assign layer_5[399] = ~(layer_4[503] & layer_4[502]); 
    wire [1:0] far_5_5500_0;    relay_conn far_5_5500_0_a(.in(layer_4[862]), .out(far_5_5500_0[0]));    relay_conn far_5_5500_0_b(.in(layer_4[902]), .out(far_5_5500_0[1]));
    assign layer_5[400] = far_5_5500_0[0] & ~far_5_5500_0[1]; 
    assign layer_5[401] = ~layer_4[660] | (layer_4[660] & layer_4[676]); 
    assign layer_5[402] = ~layer_4[726] | (layer_4[697] & layer_4[726]); 
    wire [1:0] far_5_5503_0;    relay_conn far_5_5503_0_a(.in(layer_4[589]), .out(far_5_5503_0[0]));    relay_conn far_5_5503_0_b(.in(layer_4[646]), .out(far_5_5503_0[1]));
    assign layer_5[403] = far_5_5503_0[1]; 
    wire [1:0] far_5_5504_0;    relay_conn far_5_5504_0_a(.in(layer_4[716]), .out(far_5_5504_0[0]));    relay_conn far_5_5504_0_b(.in(layer_4[643]), .out(far_5_5504_0[1]));
    wire [1:0] far_5_5504_1;    relay_conn far_5_5504_1_a(.in(far_5_5504_0[0]), .out(far_5_5504_1[0]));    relay_conn far_5_5504_1_b(.in(far_5_5504_0[1]), .out(far_5_5504_1[1]));
    assign layer_5[404] = ~far_5_5504_1[0]; 
    assign layer_5[405] = layer_4[428] & ~layer_4[425]; 
    wire [1:0] far_5_5506_0;    relay_conn far_5_5506_0_a(.in(layer_4[875]), .out(far_5_5506_0[0]));    relay_conn far_5_5506_0_b(.in(layer_4[921]), .out(far_5_5506_0[1]));
    assign layer_5[406] = far_5_5506_0[0]; 
    wire [1:0] far_5_5507_0;    relay_conn far_5_5507_0_a(.in(layer_4[615]), .out(far_5_5507_0[0]));    relay_conn far_5_5507_0_b(.in(layer_4[559]), .out(far_5_5507_0[1]));
    assign layer_5[407] = ~(far_5_5507_0[0] & far_5_5507_0[1]); 
    wire [1:0] far_5_5508_0;    relay_conn far_5_5508_0_a(.in(layer_4[251]), .out(far_5_5508_0[0]));    relay_conn far_5_5508_0_b(.in(layer_4[199]), .out(far_5_5508_0[1]));
    assign layer_5[408] = ~(far_5_5508_0[0] & far_5_5508_0[1]); 
    wire [1:0] far_5_5509_0;    relay_conn far_5_5509_0_a(.in(layer_4[985]), .out(far_5_5509_0[0]));    relay_conn far_5_5509_0_b(.in(layer_4[876]), .out(far_5_5509_0[1]));
    wire [1:0] far_5_5509_1;    relay_conn far_5_5509_1_a(.in(far_5_5509_0[0]), .out(far_5_5509_1[0]));    relay_conn far_5_5509_1_b(.in(far_5_5509_0[1]), .out(far_5_5509_1[1]));
    wire [1:0] far_5_5509_2;    relay_conn far_5_5509_2_a(.in(far_5_5509_1[0]), .out(far_5_5509_2[0]));    relay_conn far_5_5509_2_b(.in(far_5_5509_1[1]), .out(far_5_5509_2[1]));
    assign layer_5[409] = ~(far_5_5509_2[0] | far_5_5509_2[1]); 
    wire [1:0] far_5_5510_0;    relay_conn far_5_5510_0_a(.in(layer_4[670]), .out(far_5_5510_0[0]));    relay_conn far_5_5510_0_b(.in(layer_4[774]), .out(far_5_5510_0[1]));
    wire [1:0] far_5_5510_1;    relay_conn far_5_5510_1_a(.in(far_5_5510_0[0]), .out(far_5_5510_1[0]));    relay_conn far_5_5510_1_b(.in(far_5_5510_0[1]), .out(far_5_5510_1[1]));
    wire [1:0] far_5_5510_2;    relay_conn far_5_5510_2_a(.in(far_5_5510_1[0]), .out(far_5_5510_2[0]));    relay_conn far_5_5510_2_b(.in(far_5_5510_1[1]), .out(far_5_5510_2[1]));
    assign layer_5[410] = ~(far_5_5510_2[0] | far_5_5510_2[1]); 
    assign layer_5[411] = layer_4[675] & layer_4[699]; 
    wire [1:0] far_5_5512_0;    relay_conn far_5_5512_0_a(.in(layer_4[780]), .out(far_5_5512_0[0]));    relay_conn far_5_5512_0_b(.in(layer_4[684]), .out(far_5_5512_0[1]));
    wire [1:0] far_5_5512_1;    relay_conn far_5_5512_1_a(.in(far_5_5512_0[0]), .out(far_5_5512_1[0]));    relay_conn far_5_5512_1_b(.in(far_5_5512_0[1]), .out(far_5_5512_1[1]));
    wire [1:0] far_5_5512_2;    relay_conn far_5_5512_2_a(.in(far_5_5512_1[0]), .out(far_5_5512_2[0]));    relay_conn far_5_5512_2_b(.in(far_5_5512_1[1]), .out(far_5_5512_2[1]));
    assign layer_5[412] = ~far_5_5512_2[0] | (far_5_5512_2[0] & far_5_5512_2[1]); 
    wire [1:0] far_5_5513_0;    relay_conn far_5_5513_0_a(.in(layer_4[428]), .out(far_5_5513_0[0]));    relay_conn far_5_5513_0_b(.in(layer_4[357]), .out(far_5_5513_0[1]));
    wire [1:0] far_5_5513_1;    relay_conn far_5_5513_1_a(.in(far_5_5513_0[0]), .out(far_5_5513_1[0]));    relay_conn far_5_5513_1_b(.in(far_5_5513_0[1]), .out(far_5_5513_1[1]));
    assign layer_5[413] = ~far_5_5513_1[1]; 
    wire [1:0] far_5_5514_0;    relay_conn far_5_5514_0_a(.in(layer_4[511]), .out(far_5_5514_0[0]));    relay_conn far_5_5514_0_b(.in(layer_4[632]), .out(far_5_5514_0[1]));
    wire [1:0] far_5_5514_1;    relay_conn far_5_5514_1_a(.in(far_5_5514_0[0]), .out(far_5_5514_1[0]));    relay_conn far_5_5514_1_b(.in(far_5_5514_0[1]), .out(far_5_5514_1[1]));
    wire [1:0] far_5_5514_2;    relay_conn far_5_5514_2_a(.in(far_5_5514_1[0]), .out(far_5_5514_2[0]));    relay_conn far_5_5514_2_b(.in(far_5_5514_1[1]), .out(far_5_5514_2[1]));
    assign layer_5[414] = ~far_5_5514_2[1]; 
    wire [1:0] far_5_5515_0;    relay_conn far_5_5515_0_a(.in(layer_4[852]), .out(far_5_5515_0[0]));    relay_conn far_5_5515_0_b(.in(layer_4[898]), .out(far_5_5515_0[1]));
    assign layer_5[415] = ~far_5_5515_0[0]; 
    wire [1:0] far_5_5516_0;    relay_conn far_5_5516_0_a(.in(layer_4[520]), .out(far_5_5516_0[0]));    relay_conn far_5_5516_0_b(.in(layer_4[602]), .out(far_5_5516_0[1]));
    wire [1:0] far_5_5516_1;    relay_conn far_5_5516_1_a(.in(far_5_5516_0[0]), .out(far_5_5516_1[0]));    relay_conn far_5_5516_1_b(.in(far_5_5516_0[1]), .out(far_5_5516_1[1]));
    assign layer_5[416] = far_5_5516_1[1] & ~far_5_5516_1[0]; 
    wire [1:0] far_5_5517_0;    relay_conn far_5_5517_0_a(.in(layer_4[333]), .out(far_5_5517_0[0]));    relay_conn far_5_5517_0_b(.in(layer_4[446]), .out(far_5_5517_0[1]));
    wire [1:0] far_5_5517_1;    relay_conn far_5_5517_1_a(.in(far_5_5517_0[0]), .out(far_5_5517_1[0]));    relay_conn far_5_5517_1_b(.in(far_5_5517_0[1]), .out(far_5_5517_1[1]));
    wire [1:0] far_5_5517_2;    relay_conn far_5_5517_2_a(.in(far_5_5517_1[0]), .out(far_5_5517_2[0]));    relay_conn far_5_5517_2_b(.in(far_5_5517_1[1]), .out(far_5_5517_2[1]));
    assign layer_5[417] = ~far_5_5517_2[0] | (far_5_5517_2[0] & far_5_5517_2[1]); 
    wire [1:0] far_5_5518_0;    relay_conn far_5_5518_0_a(.in(layer_4[472]), .out(far_5_5518_0[0]));    relay_conn far_5_5518_0_b(.in(layer_4[552]), .out(far_5_5518_0[1]));
    wire [1:0] far_5_5518_1;    relay_conn far_5_5518_1_a(.in(far_5_5518_0[0]), .out(far_5_5518_1[0]));    relay_conn far_5_5518_1_b(.in(far_5_5518_0[1]), .out(far_5_5518_1[1]));
    assign layer_5[418] = ~far_5_5518_1[0]; 
    wire [1:0] far_5_5519_0;    relay_conn far_5_5519_0_a(.in(layer_4[312]), .out(far_5_5519_0[0]));    relay_conn far_5_5519_0_b(.in(layer_4[274]), .out(far_5_5519_0[1]));
    assign layer_5[419] = far_5_5519_0[0] | far_5_5519_0[1]; 
    wire [1:0] far_5_5520_0;    relay_conn far_5_5520_0_a(.in(layer_4[930]), .out(far_5_5520_0[0]));    relay_conn far_5_5520_0_b(.in(layer_4[867]), .out(far_5_5520_0[1]));
    assign layer_5[420] = far_5_5520_0[1] & ~far_5_5520_0[0]; 
    wire [1:0] far_5_5521_0;    relay_conn far_5_5521_0_a(.in(layer_4[689]), .out(far_5_5521_0[0]));    relay_conn far_5_5521_0_b(.in(layer_4[789]), .out(far_5_5521_0[1]));
    wire [1:0] far_5_5521_1;    relay_conn far_5_5521_1_a(.in(far_5_5521_0[0]), .out(far_5_5521_1[0]));    relay_conn far_5_5521_1_b(.in(far_5_5521_0[1]), .out(far_5_5521_1[1]));
    wire [1:0] far_5_5521_2;    relay_conn far_5_5521_2_a(.in(far_5_5521_1[0]), .out(far_5_5521_2[0]));    relay_conn far_5_5521_2_b(.in(far_5_5521_1[1]), .out(far_5_5521_2[1]));
    assign layer_5[421] = ~far_5_5521_2[1] | (far_5_5521_2[0] & far_5_5521_2[1]); 
    wire [1:0] far_5_5522_0;    relay_conn far_5_5522_0_a(.in(layer_4[666]), .out(far_5_5522_0[0]));    relay_conn far_5_5522_0_b(.in(layer_4[559]), .out(far_5_5522_0[1]));
    wire [1:0] far_5_5522_1;    relay_conn far_5_5522_1_a(.in(far_5_5522_0[0]), .out(far_5_5522_1[0]));    relay_conn far_5_5522_1_b(.in(far_5_5522_0[1]), .out(far_5_5522_1[1]));
    wire [1:0] far_5_5522_2;    relay_conn far_5_5522_2_a(.in(far_5_5522_1[0]), .out(far_5_5522_2[0]));    relay_conn far_5_5522_2_b(.in(far_5_5522_1[1]), .out(far_5_5522_2[1]));
    assign layer_5[422] = ~(far_5_5522_2[0] & far_5_5522_2[1]); 
    wire [1:0] far_5_5523_0;    relay_conn far_5_5523_0_a(.in(layer_4[316]), .out(far_5_5523_0[0]));    relay_conn far_5_5523_0_b(.in(layer_4[232]), .out(far_5_5523_0[1]));
    wire [1:0] far_5_5523_1;    relay_conn far_5_5523_1_a(.in(far_5_5523_0[0]), .out(far_5_5523_1[0]));    relay_conn far_5_5523_1_b(.in(far_5_5523_0[1]), .out(far_5_5523_1[1]));
    assign layer_5[423] = ~far_5_5523_1[0]; 
    assign layer_5[424] = ~(layer_4[409] & layer_4[401]); 
    wire [1:0] far_5_5525_0;    relay_conn far_5_5525_0_a(.in(layer_4[10]), .out(far_5_5525_0[0]));    relay_conn far_5_5525_0_b(.in(layer_4[105]), .out(far_5_5525_0[1]));
    wire [1:0] far_5_5525_1;    relay_conn far_5_5525_1_a(.in(far_5_5525_0[0]), .out(far_5_5525_1[0]));    relay_conn far_5_5525_1_b(.in(far_5_5525_0[1]), .out(far_5_5525_1[1]));
    assign layer_5[425] = ~(far_5_5525_1[0] & far_5_5525_1[1]); 
    assign layer_5[426] = ~layer_4[282]; 
    wire [1:0] far_5_5527_0;    relay_conn far_5_5527_0_a(.in(layer_4[764]), .out(far_5_5527_0[0]));    relay_conn far_5_5527_0_b(.in(layer_4[805]), .out(far_5_5527_0[1]));
    assign layer_5[427] = far_5_5527_0[1]; 
    wire [1:0] far_5_5528_0;    relay_conn far_5_5528_0_a(.in(layer_4[273]), .out(far_5_5528_0[0]));    relay_conn far_5_5528_0_b(.in(layer_4[220]), .out(far_5_5528_0[1]));
    assign layer_5[428] = far_5_5528_0[1] & ~far_5_5528_0[0]; 
    assign layer_5[429] = ~layer_4[675] | (layer_4[675] & layer_4[681]); 
    wire [1:0] far_5_5530_0;    relay_conn far_5_5530_0_a(.in(layer_4[429]), .out(far_5_5530_0[0]));    relay_conn far_5_5530_0_b(.in(layer_4[369]), .out(far_5_5530_0[1]));
    assign layer_5[430] = far_5_5530_0[0] | far_5_5530_0[1]; 
    wire [1:0] far_5_5531_0;    relay_conn far_5_5531_0_a(.in(layer_4[784]), .out(far_5_5531_0[0]));    relay_conn far_5_5531_0_b(.in(layer_4[719]), .out(far_5_5531_0[1]));
    wire [1:0] far_5_5531_1;    relay_conn far_5_5531_1_a(.in(far_5_5531_0[0]), .out(far_5_5531_1[0]));    relay_conn far_5_5531_1_b(.in(far_5_5531_0[1]), .out(far_5_5531_1[1]));
    assign layer_5[431] = far_5_5531_1[0] & ~far_5_5531_1[1]; 
    wire [1:0] far_5_5532_0;    relay_conn far_5_5532_0_a(.in(layer_4[513]), .out(far_5_5532_0[0]));    relay_conn far_5_5532_0_b(.in(layer_4[472]), .out(far_5_5532_0[1]));
    assign layer_5[432] = far_5_5532_0[1]; 
    assign layer_5[433] = layer_4[692] & ~layer_4[661]; 
    assign layer_5[434] = layer_4[174] | layer_4[166]; 
    wire [1:0] far_5_5535_0;    relay_conn far_5_5535_0_a(.in(layer_4[542]), .out(far_5_5535_0[0]));    relay_conn far_5_5535_0_b(.in(layer_4[644]), .out(far_5_5535_0[1]));
    wire [1:0] far_5_5535_1;    relay_conn far_5_5535_1_a(.in(far_5_5535_0[0]), .out(far_5_5535_1[0]));    relay_conn far_5_5535_1_b(.in(far_5_5535_0[1]), .out(far_5_5535_1[1]));
    wire [1:0] far_5_5535_2;    relay_conn far_5_5535_2_a(.in(far_5_5535_1[0]), .out(far_5_5535_2[0]));    relay_conn far_5_5535_2_b(.in(far_5_5535_1[1]), .out(far_5_5535_2[1]));
    assign layer_5[435] = ~far_5_5535_2[0]; 
    wire [1:0] far_5_5536_0;    relay_conn far_5_5536_0_a(.in(layer_4[71]), .out(far_5_5536_0[0]));    relay_conn far_5_5536_0_b(.in(layer_4[135]), .out(far_5_5536_0[1]));
    wire [1:0] far_5_5536_1;    relay_conn far_5_5536_1_a(.in(far_5_5536_0[0]), .out(far_5_5536_1[0]));    relay_conn far_5_5536_1_b(.in(far_5_5536_0[1]), .out(far_5_5536_1[1]));
    assign layer_5[436] = far_5_5536_1[0] ^ far_5_5536_1[1]; 
    wire [1:0] far_5_5537_0;    relay_conn far_5_5537_0_a(.in(layer_4[977]), .out(far_5_5537_0[0]));    relay_conn far_5_5537_0_b(.in(layer_4[875]), .out(far_5_5537_0[1]));
    wire [1:0] far_5_5537_1;    relay_conn far_5_5537_1_a(.in(far_5_5537_0[0]), .out(far_5_5537_1[0]));    relay_conn far_5_5537_1_b(.in(far_5_5537_0[1]), .out(far_5_5537_1[1]));
    wire [1:0] far_5_5537_2;    relay_conn far_5_5537_2_a(.in(far_5_5537_1[0]), .out(far_5_5537_2[0]));    relay_conn far_5_5537_2_b(.in(far_5_5537_1[1]), .out(far_5_5537_2[1]));
    assign layer_5[437] = ~far_5_5537_2[0]; 
    wire [1:0] far_5_5538_0;    relay_conn far_5_5538_0_a(.in(layer_4[644]), .out(far_5_5538_0[0]));    relay_conn far_5_5538_0_b(.in(layer_4[768]), .out(far_5_5538_0[1]));
    wire [1:0] far_5_5538_1;    relay_conn far_5_5538_1_a(.in(far_5_5538_0[0]), .out(far_5_5538_1[0]));    relay_conn far_5_5538_1_b(.in(far_5_5538_0[1]), .out(far_5_5538_1[1]));
    wire [1:0] far_5_5538_2;    relay_conn far_5_5538_2_a(.in(far_5_5538_1[0]), .out(far_5_5538_2[0]));    relay_conn far_5_5538_2_b(.in(far_5_5538_1[1]), .out(far_5_5538_2[1]));
    assign layer_5[438] = ~(far_5_5538_2[0] ^ far_5_5538_2[1]); 
    wire [1:0] far_5_5539_0;    relay_conn far_5_5539_0_a(.in(layer_4[719]), .out(far_5_5539_0[0]));    relay_conn far_5_5539_0_b(.in(layer_4[847]), .out(far_5_5539_0[1]));
    wire [1:0] far_5_5539_1;    relay_conn far_5_5539_1_a(.in(far_5_5539_0[0]), .out(far_5_5539_1[0]));    relay_conn far_5_5539_1_b(.in(far_5_5539_0[1]), .out(far_5_5539_1[1]));
    wire [1:0] far_5_5539_2;    relay_conn far_5_5539_2_a(.in(far_5_5539_1[0]), .out(far_5_5539_2[0]));    relay_conn far_5_5539_2_b(.in(far_5_5539_1[1]), .out(far_5_5539_2[1]));
    wire [1:0] far_5_5539_3;    relay_conn far_5_5539_3_a(.in(far_5_5539_2[0]), .out(far_5_5539_3[0]));    relay_conn far_5_5539_3_b(.in(far_5_5539_2[1]), .out(far_5_5539_3[1]));
    assign layer_5[439] = ~(far_5_5539_3[0] | far_5_5539_3[1]); 
    wire [1:0] far_5_5540_0;    relay_conn far_5_5540_0_a(.in(layer_4[62]), .out(far_5_5540_0[0]));    relay_conn far_5_5540_0_b(.in(layer_4[23]), .out(far_5_5540_0[1]));
    assign layer_5[440] = ~far_5_5540_0[1] | (far_5_5540_0[0] & far_5_5540_0[1]); 
    assign layer_5[441] = ~layer_4[888]; 
    wire [1:0] far_5_5542_0;    relay_conn far_5_5542_0_a(.in(layer_4[31]), .out(far_5_5542_0[0]));    relay_conn far_5_5542_0_b(.in(layer_4[72]), .out(far_5_5542_0[1]));
    assign layer_5[442] = far_5_5542_0[0] ^ far_5_5542_0[1]; 
    wire [1:0] far_5_5543_0;    relay_conn far_5_5543_0_a(.in(layer_4[926]), .out(far_5_5543_0[0]));    relay_conn far_5_5543_0_b(.in(layer_4[888]), .out(far_5_5543_0[1]));
    assign layer_5[443] = far_5_5543_0[0] & far_5_5543_0[1]; 
    wire [1:0] far_5_5544_0;    relay_conn far_5_5544_0_a(.in(layer_4[520]), .out(far_5_5544_0[0]));    relay_conn far_5_5544_0_b(.in(layer_4[477]), .out(far_5_5544_0[1]));
    assign layer_5[444] = ~(far_5_5544_0[0] | far_5_5544_0[1]); 
    assign layer_5[445] = layer_4[632] ^ layer_4[661]; 
    wire [1:0] far_5_5546_0;    relay_conn far_5_5546_0_a(.in(layer_4[624]), .out(far_5_5546_0[0]));    relay_conn far_5_5546_0_b(.in(layer_4[710]), .out(far_5_5546_0[1]));
    wire [1:0] far_5_5546_1;    relay_conn far_5_5546_1_a(.in(far_5_5546_0[0]), .out(far_5_5546_1[0]));    relay_conn far_5_5546_1_b(.in(far_5_5546_0[1]), .out(far_5_5546_1[1]));
    assign layer_5[446] = far_5_5546_1[0] ^ far_5_5546_1[1]; 
    assign layer_5[447] = ~(layer_4[134] ^ layer_4[149]); 
    assign layer_5[448] = layer_4[995] & layer_4[997]; 
    wire [1:0] far_5_5549_0;    relay_conn far_5_5549_0_a(.in(layer_4[218]), .out(far_5_5549_0[0]));    relay_conn far_5_5549_0_b(.in(layer_4[301]), .out(far_5_5549_0[1]));
    wire [1:0] far_5_5549_1;    relay_conn far_5_5549_1_a(.in(far_5_5549_0[0]), .out(far_5_5549_1[0]));    relay_conn far_5_5549_1_b(.in(far_5_5549_0[1]), .out(far_5_5549_1[1]));
    assign layer_5[449] = far_5_5549_1[0] | far_5_5549_1[1]; 
    wire [1:0] far_5_5550_0;    relay_conn far_5_5550_0_a(.in(layer_4[672]), .out(far_5_5550_0[0]));    relay_conn far_5_5550_0_b(.in(layer_4[565]), .out(far_5_5550_0[1]));
    wire [1:0] far_5_5550_1;    relay_conn far_5_5550_1_a(.in(far_5_5550_0[0]), .out(far_5_5550_1[0]));    relay_conn far_5_5550_1_b(.in(far_5_5550_0[1]), .out(far_5_5550_1[1]));
    wire [1:0] far_5_5550_2;    relay_conn far_5_5550_2_a(.in(far_5_5550_1[0]), .out(far_5_5550_2[0]));    relay_conn far_5_5550_2_b(.in(far_5_5550_1[1]), .out(far_5_5550_2[1]));
    assign layer_5[450] = ~(far_5_5550_2[0] | far_5_5550_2[1]); 
    wire [1:0] far_5_5551_0;    relay_conn far_5_5551_0_a(.in(layer_4[378]), .out(far_5_5551_0[0]));    relay_conn far_5_5551_0_b(.in(layer_4[314]), .out(far_5_5551_0[1]));
    wire [1:0] far_5_5551_1;    relay_conn far_5_5551_1_a(.in(far_5_5551_0[0]), .out(far_5_5551_1[0]));    relay_conn far_5_5551_1_b(.in(far_5_5551_0[1]), .out(far_5_5551_1[1]));
    assign layer_5[451] = ~far_5_5551_1[0]; 
    wire [1:0] far_5_5552_0;    relay_conn far_5_5552_0_a(.in(layer_4[656]), .out(far_5_5552_0[0]));    relay_conn far_5_5552_0_b(.in(layer_4[704]), .out(far_5_5552_0[1]));
    assign layer_5[452] = ~far_5_5552_0[1] | (far_5_5552_0[0] & far_5_5552_0[1]); 
    assign layer_5[453] = layer_4[953]; 
    assign layer_5[454] = ~(layer_4[168] & layer_4[176]); 
    wire [1:0] far_5_5555_0;    relay_conn far_5_5555_0_a(.in(layer_4[305]), .out(far_5_5555_0[0]));    relay_conn far_5_5555_0_b(.in(layer_4[232]), .out(far_5_5555_0[1]));
    wire [1:0] far_5_5555_1;    relay_conn far_5_5555_1_a(.in(far_5_5555_0[0]), .out(far_5_5555_1[0]));    relay_conn far_5_5555_1_b(.in(far_5_5555_0[1]), .out(far_5_5555_1[1]));
    assign layer_5[455] = far_5_5555_1[1] & ~far_5_5555_1[0]; 
    wire [1:0] far_5_5556_0;    relay_conn far_5_5556_0_a(.in(layer_4[253]), .out(far_5_5556_0[0]));    relay_conn far_5_5556_0_b(.in(layer_4[381]), .out(far_5_5556_0[1]));
    wire [1:0] far_5_5556_1;    relay_conn far_5_5556_1_a(.in(far_5_5556_0[0]), .out(far_5_5556_1[0]));    relay_conn far_5_5556_1_b(.in(far_5_5556_0[1]), .out(far_5_5556_1[1]));
    wire [1:0] far_5_5556_2;    relay_conn far_5_5556_2_a(.in(far_5_5556_1[0]), .out(far_5_5556_2[0]));    relay_conn far_5_5556_2_b(.in(far_5_5556_1[1]), .out(far_5_5556_2[1]));
    wire [1:0] far_5_5556_3;    relay_conn far_5_5556_3_a(.in(far_5_5556_2[0]), .out(far_5_5556_3[0]));    relay_conn far_5_5556_3_b(.in(far_5_5556_2[1]), .out(far_5_5556_3[1]));
    assign layer_5[456] = far_5_5556_3[1]; 
    wire [1:0] far_5_5557_0;    relay_conn far_5_5557_0_a(.in(layer_4[928]), .out(far_5_5557_0[0]));    relay_conn far_5_5557_0_b(.in(layer_4[861]), .out(far_5_5557_0[1]));
    wire [1:0] far_5_5557_1;    relay_conn far_5_5557_1_a(.in(far_5_5557_0[0]), .out(far_5_5557_1[0]));    relay_conn far_5_5557_1_b(.in(far_5_5557_0[1]), .out(far_5_5557_1[1]));
    assign layer_5[457] = ~(far_5_5557_1[0] | far_5_5557_1[1]); 
    wire [1:0] far_5_5558_0;    relay_conn far_5_5558_0_a(.in(layer_4[333]), .out(far_5_5558_0[0]));    relay_conn far_5_5558_0_b(.in(layer_4[435]), .out(far_5_5558_0[1]));
    wire [1:0] far_5_5558_1;    relay_conn far_5_5558_1_a(.in(far_5_5558_0[0]), .out(far_5_5558_1[0]));    relay_conn far_5_5558_1_b(.in(far_5_5558_0[1]), .out(far_5_5558_1[1]));
    wire [1:0] far_5_5558_2;    relay_conn far_5_5558_2_a(.in(far_5_5558_1[0]), .out(far_5_5558_2[0]));    relay_conn far_5_5558_2_b(.in(far_5_5558_1[1]), .out(far_5_5558_2[1]));
    assign layer_5[458] = far_5_5558_2[1]; 
    wire [1:0] far_5_5559_0;    relay_conn far_5_5559_0_a(.in(layer_4[109]), .out(far_5_5559_0[0]));    relay_conn far_5_5559_0_b(.in(layer_4[144]), .out(far_5_5559_0[1]));
    assign layer_5[459] = ~(far_5_5559_0[0] & far_5_5559_0[1]); 
    wire [1:0] far_5_5560_0;    relay_conn far_5_5560_0_a(.in(layer_4[443]), .out(far_5_5560_0[0]));    relay_conn far_5_5560_0_b(.in(layer_4[495]), .out(far_5_5560_0[1]));
    assign layer_5[460] = far_5_5560_0[0] ^ far_5_5560_0[1]; 
    wire [1:0] far_5_5561_0;    relay_conn far_5_5561_0_a(.in(layer_4[619]), .out(far_5_5561_0[0]));    relay_conn far_5_5561_0_b(.in(layer_4[500]), .out(far_5_5561_0[1]));
    wire [1:0] far_5_5561_1;    relay_conn far_5_5561_1_a(.in(far_5_5561_0[0]), .out(far_5_5561_1[0]));    relay_conn far_5_5561_1_b(.in(far_5_5561_0[1]), .out(far_5_5561_1[1]));
    wire [1:0] far_5_5561_2;    relay_conn far_5_5561_2_a(.in(far_5_5561_1[0]), .out(far_5_5561_2[0]));    relay_conn far_5_5561_2_b(.in(far_5_5561_1[1]), .out(far_5_5561_2[1]));
    assign layer_5[461] = far_5_5561_2[0] & far_5_5561_2[1]; 
    wire [1:0] far_5_5562_0;    relay_conn far_5_5562_0_a(.in(layer_4[415]), .out(far_5_5562_0[0]));    relay_conn far_5_5562_0_b(.in(layer_4[451]), .out(far_5_5562_0[1]));
    assign layer_5[462] = ~(far_5_5562_0[0] | far_5_5562_0[1]); 
    wire [1:0] far_5_5563_0;    relay_conn far_5_5563_0_a(.in(layer_4[170]), .out(far_5_5563_0[0]));    relay_conn far_5_5563_0_b(.in(layer_4[90]), .out(far_5_5563_0[1]));
    wire [1:0] far_5_5563_1;    relay_conn far_5_5563_1_a(.in(far_5_5563_0[0]), .out(far_5_5563_1[0]));    relay_conn far_5_5563_1_b(.in(far_5_5563_0[1]), .out(far_5_5563_1[1]));
    assign layer_5[463] = ~far_5_5563_1[1]; 
    wire [1:0] far_5_5564_0;    relay_conn far_5_5564_0_a(.in(layer_4[718]), .out(far_5_5564_0[0]));    relay_conn far_5_5564_0_b(.in(layer_4[790]), .out(far_5_5564_0[1]));
    wire [1:0] far_5_5564_1;    relay_conn far_5_5564_1_a(.in(far_5_5564_0[0]), .out(far_5_5564_1[0]));    relay_conn far_5_5564_1_b(.in(far_5_5564_0[1]), .out(far_5_5564_1[1]));
    assign layer_5[464] = ~far_5_5564_1[1]; 
    wire [1:0] far_5_5565_0;    relay_conn far_5_5565_0_a(.in(layer_4[835]), .out(far_5_5565_0[0]));    relay_conn far_5_5565_0_b(.in(layer_4[875]), .out(far_5_5565_0[1]));
    assign layer_5[465] = ~(far_5_5565_0[0] ^ far_5_5565_0[1]); 
    assign layer_5[466] = ~(layer_4[10] & layer_4[20]); 
    wire [1:0] far_5_5567_0;    relay_conn far_5_5567_0_a(.in(layer_4[826]), .out(far_5_5567_0[0]));    relay_conn far_5_5567_0_b(.in(layer_4[710]), .out(far_5_5567_0[1]));
    wire [1:0] far_5_5567_1;    relay_conn far_5_5567_1_a(.in(far_5_5567_0[0]), .out(far_5_5567_1[0]));    relay_conn far_5_5567_1_b(.in(far_5_5567_0[1]), .out(far_5_5567_1[1]));
    wire [1:0] far_5_5567_2;    relay_conn far_5_5567_2_a(.in(far_5_5567_1[0]), .out(far_5_5567_2[0]));    relay_conn far_5_5567_2_b(.in(far_5_5567_1[1]), .out(far_5_5567_2[1]));
    assign layer_5[467] = far_5_5567_2[1]; 
    assign layer_5[468] = ~layer_4[225] | (layer_4[202] & layer_4[225]); 
    assign layer_5[469] = layer_4[973]; 
    wire [1:0] far_5_5570_0;    relay_conn far_5_5570_0_a(.in(layer_4[177]), .out(far_5_5570_0[0]));    relay_conn far_5_5570_0_b(.in(layer_4[258]), .out(far_5_5570_0[1]));
    wire [1:0] far_5_5570_1;    relay_conn far_5_5570_1_a(.in(far_5_5570_0[0]), .out(far_5_5570_1[0]));    relay_conn far_5_5570_1_b(.in(far_5_5570_0[1]), .out(far_5_5570_1[1]));
    assign layer_5[470] = ~far_5_5570_1[1]; 
    wire [1:0] far_5_5571_0;    relay_conn far_5_5571_0_a(.in(layer_4[650]), .out(far_5_5571_0[0]));    relay_conn far_5_5571_0_b(.in(layer_4[716]), .out(far_5_5571_0[1]));
    wire [1:0] far_5_5571_1;    relay_conn far_5_5571_1_a(.in(far_5_5571_0[0]), .out(far_5_5571_1[0]));    relay_conn far_5_5571_1_b(.in(far_5_5571_0[1]), .out(far_5_5571_1[1]));
    assign layer_5[471] = ~far_5_5571_1[0] | (far_5_5571_1[0] & far_5_5571_1[1]); 
    wire [1:0] far_5_5572_0;    relay_conn far_5_5572_0_a(.in(layer_4[619]), .out(far_5_5572_0[0]));    relay_conn far_5_5572_0_b(.in(layer_4[721]), .out(far_5_5572_0[1]));
    wire [1:0] far_5_5572_1;    relay_conn far_5_5572_1_a(.in(far_5_5572_0[0]), .out(far_5_5572_1[0]));    relay_conn far_5_5572_1_b(.in(far_5_5572_0[1]), .out(far_5_5572_1[1]));
    wire [1:0] far_5_5572_2;    relay_conn far_5_5572_2_a(.in(far_5_5572_1[0]), .out(far_5_5572_2[0]));    relay_conn far_5_5572_2_b(.in(far_5_5572_1[1]), .out(far_5_5572_2[1]));
    assign layer_5[472] = far_5_5572_2[1]; 
    wire [1:0] far_5_5573_0;    relay_conn far_5_5573_0_a(.in(layer_4[832]), .out(far_5_5573_0[0]));    relay_conn far_5_5573_0_b(.in(layer_4[902]), .out(far_5_5573_0[1]));
    wire [1:0] far_5_5573_1;    relay_conn far_5_5573_1_a(.in(far_5_5573_0[0]), .out(far_5_5573_1[0]));    relay_conn far_5_5573_1_b(.in(far_5_5573_0[1]), .out(far_5_5573_1[1]));
    assign layer_5[473] = far_5_5573_1[1] & ~far_5_5573_1[0]; 
    wire [1:0] far_5_5574_0;    relay_conn far_5_5574_0_a(.in(layer_4[1012]), .out(far_5_5574_0[0]));    relay_conn far_5_5574_0_b(.in(layer_4[914]), .out(far_5_5574_0[1]));
    wire [1:0] far_5_5574_1;    relay_conn far_5_5574_1_a(.in(far_5_5574_0[0]), .out(far_5_5574_1[0]));    relay_conn far_5_5574_1_b(.in(far_5_5574_0[1]), .out(far_5_5574_1[1]));
    wire [1:0] far_5_5574_2;    relay_conn far_5_5574_2_a(.in(far_5_5574_1[0]), .out(far_5_5574_2[0]));    relay_conn far_5_5574_2_b(.in(far_5_5574_1[1]), .out(far_5_5574_2[1]));
    assign layer_5[474] = ~(far_5_5574_2[0] & far_5_5574_2[1]); 
    wire [1:0] far_5_5575_0;    relay_conn far_5_5575_0_a(.in(layer_4[523]), .out(far_5_5575_0[0]));    relay_conn far_5_5575_0_b(.in(layer_4[597]), .out(far_5_5575_0[1]));
    wire [1:0] far_5_5575_1;    relay_conn far_5_5575_1_a(.in(far_5_5575_0[0]), .out(far_5_5575_1[0]));    relay_conn far_5_5575_1_b(.in(far_5_5575_0[1]), .out(far_5_5575_1[1]));
    assign layer_5[475] = far_5_5575_1[0] | far_5_5575_1[1]; 
    wire [1:0] far_5_5576_0;    relay_conn far_5_5576_0_a(.in(layer_4[387]), .out(far_5_5576_0[0]));    relay_conn far_5_5576_0_b(.in(layer_4[464]), .out(far_5_5576_0[1]));
    wire [1:0] far_5_5576_1;    relay_conn far_5_5576_1_a(.in(far_5_5576_0[0]), .out(far_5_5576_1[0]));    relay_conn far_5_5576_1_b(.in(far_5_5576_0[1]), .out(far_5_5576_1[1]));
    assign layer_5[476] = ~far_5_5576_1[1] | (far_5_5576_1[0] & far_5_5576_1[1]); 
    wire [1:0] far_5_5577_0;    relay_conn far_5_5577_0_a(.in(layer_4[939]), .out(far_5_5577_0[0]));    relay_conn far_5_5577_0_b(.in(layer_4[860]), .out(far_5_5577_0[1]));
    wire [1:0] far_5_5577_1;    relay_conn far_5_5577_1_a(.in(far_5_5577_0[0]), .out(far_5_5577_1[0]));    relay_conn far_5_5577_1_b(.in(far_5_5577_0[1]), .out(far_5_5577_1[1]));
    assign layer_5[477] = ~(far_5_5577_1[0] | far_5_5577_1[1]); 
    wire [1:0] far_5_5578_0;    relay_conn far_5_5578_0_a(.in(layer_4[100]), .out(far_5_5578_0[0]));    relay_conn far_5_5578_0_b(.in(layer_4[134]), .out(far_5_5578_0[1]));
    assign layer_5[478] = ~(far_5_5578_0[0] | far_5_5578_0[1]); 
    assign layer_5[479] = layer_4[1013] & layer_4[991]; 
    wire [1:0] far_5_5580_0;    relay_conn far_5_5580_0_a(.in(layer_4[149]), .out(far_5_5580_0[0]));    relay_conn far_5_5580_0_b(.in(layer_4[96]), .out(far_5_5580_0[1]));
    assign layer_5[480] = ~(far_5_5580_0[0] & far_5_5580_0[1]); 
    wire [1:0] far_5_5581_0;    relay_conn far_5_5581_0_a(.in(layer_4[122]), .out(far_5_5581_0[0]));    relay_conn far_5_5581_0_b(.in(layer_4[4]), .out(far_5_5581_0[1]));
    wire [1:0] far_5_5581_1;    relay_conn far_5_5581_1_a(.in(far_5_5581_0[0]), .out(far_5_5581_1[0]));    relay_conn far_5_5581_1_b(.in(far_5_5581_0[1]), .out(far_5_5581_1[1]));
    wire [1:0] far_5_5581_2;    relay_conn far_5_5581_2_a(.in(far_5_5581_1[0]), .out(far_5_5581_2[0]));    relay_conn far_5_5581_2_b(.in(far_5_5581_1[1]), .out(far_5_5581_2[1]));
    assign layer_5[481] = far_5_5581_2[1]; 
    wire [1:0] far_5_5582_0;    relay_conn far_5_5582_0_a(.in(layer_4[812]), .out(far_5_5582_0[0]));    relay_conn far_5_5582_0_b(.in(layer_4[875]), .out(far_5_5582_0[1]));
    assign layer_5[482] = far_5_5582_0[1] & ~far_5_5582_0[0]; 
    wire [1:0] far_5_5583_0;    relay_conn far_5_5583_0_a(.in(layer_4[495]), .out(far_5_5583_0[0]));    relay_conn far_5_5583_0_b(.in(layer_4[452]), .out(far_5_5583_0[1]));
    assign layer_5[483] = ~(far_5_5583_0[0] & far_5_5583_0[1]); 
    wire [1:0] far_5_5584_0;    relay_conn far_5_5584_0_a(.in(layer_4[952]), .out(far_5_5584_0[0]));    relay_conn far_5_5584_0_b(.in(layer_4[879]), .out(far_5_5584_0[1]));
    wire [1:0] far_5_5584_1;    relay_conn far_5_5584_1_a(.in(far_5_5584_0[0]), .out(far_5_5584_1[0]));    relay_conn far_5_5584_1_b(.in(far_5_5584_0[1]), .out(far_5_5584_1[1]));
    assign layer_5[484] = far_5_5584_1[0] & far_5_5584_1[1]; 
    wire [1:0] far_5_5585_0;    relay_conn far_5_5585_0_a(.in(layer_4[661]), .out(far_5_5585_0[0]));    relay_conn far_5_5585_0_b(.in(layer_4[555]), .out(far_5_5585_0[1]));
    wire [1:0] far_5_5585_1;    relay_conn far_5_5585_1_a(.in(far_5_5585_0[0]), .out(far_5_5585_1[0]));    relay_conn far_5_5585_1_b(.in(far_5_5585_0[1]), .out(far_5_5585_1[1]));
    wire [1:0] far_5_5585_2;    relay_conn far_5_5585_2_a(.in(far_5_5585_1[0]), .out(far_5_5585_2[0]));    relay_conn far_5_5585_2_b(.in(far_5_5585_1[1]), .out(far_5_5585_2[1]));
    assign layer_5[485] = far_5_5585_2[1] & ~far_5_5585_2[0]; 
    wire [1:0] far_5_5586_0;    relay_conn far_5_5586_0_a(.in(layer_4[535]), .out(far_5_5586_0[0]));    relay_conn far_5_5586_0_b(.in(layer_4[424]), .out(far_5_5586_0[1]));
    wire [1:0] far_5_5586_1;    relay_conn far_5_5586_1_a(.in(far_5_5586_0[0]), .out(far_5_5586_1[0]));    relay_conn far_5_5586_1_b(.in(far_5_5586_0[1]), .out(far_5_5586_1[1]));
    wire [1:0] far_5_5586_2;    relay_conn far_5_5586_2_a(.in(far_5_5586_1[0]), .out(far_5_5586_2[0]));    relay_conn far_5_5586_2_b(.in(far_5_5586_1[1]), .out(far_5_5586_2[1]));
    assign layer_5[486] = ~far_5_5586_2[1] | (far_5_5586_2[0] & far_5_5586_2[1]); 
    assign layer_5[487] = layer_4[357]; 
    wire [1:0] far_5_5588_0;    relay_conn far_5_5588_0_a(.in(layer_4[920]), .out(far_5_5588_0[0]));    relay_conn far_5_5588_0_b(.in(layer_4[961]), .out(far_5_5588_0[1]));
    assign layer_5[488] = far_5_5588_0[1] & ~far_5_5588_0[0]; 
    wire [1:0] far_5_5589_0;    relay_conn far_5_5589_0_a(.in(layer_4[683]), .out(far_5_5589_0[0]));    relay_conn far_5_5589_0_b(.in(layer_4[780]), .out(far_5_5589_0[1]));
    wire [1:0] far_5_5589_1;    relay_conn far_5_5589_1_a(.in(far_5_5589_0[0]), .out(far_5_5589_1[0]));    relay_conn far_5_5589_1_b(.in(far_5_5589_0[1]), .out(far_5_5589_1[1]));
    wire [1:0] far_5_5589_2;    relay_conn far_5_5589_2_a(.in(far_5_5589_1[0]), .out(far_5_5589_2[0]));    relay_conn far_5_5589_2_b(.in(far_5_5589_1[1]), .out(far_5_5589_2[1]));
    assign layer_5[489] = far_5_5589_2[0] & ~far_5_5589_2[1]; 
    wire [1:0] far_5_5590_0;    relay_conn far_5_5590_0_a(.in(layer_4[243]), .out(far_5_5590_0[0]));    relay_conn far_5_5590_0_b(.in(layer_4[124]), .out(far_5_5590_0[1]));
    wire [1:0] far_5_5590_1;    relay_conn far_5_5590_1_a(.in(far_5_5590_0[0]), .out(far_5_5590_1[0]));    relay_conn far_5_5590_1_b(.in(far_5_5590_0[1]), .out(far_5_5590_1[1]));
    wire [1:0] far_5_5590_2;    relay_conn far_5_5590_2_a(.in(far_5_5590_1[0]), .out(far_5_5590_2[0]));    relay_conn far_5_5590_2_b(.in(far_5_5590_1[1]), .out(far_5_5590_2[1]));
    assign layer_5[490] = ~far_5_5590_2[0] | (far_5_5590_2[0] & far_5_5590_2[1]); 
    wire [1:0] far_5_5591_0;    relay_conn far_5_5591_0_a(.in(layer_4[823]), .out(far_5_5591_0[0]));    relay_conn far_5_5591_0_b(.in(layer_4[735]), .out(far_5_5591_0[1]));
    wire [1:0] far_5_5591_1;    relay_conn far_5_5591_1_a(.in(far_5_5591_0[0]), .out(far_5_5591_1[0]));    relay_conn far_5_5591_1_b(.in(far_5_5591_0[1]), .out(far_5_5591_1[1]));
    assign layer_5[491] = far_5_5591_1[0]; 
    wire [1:0] far_5_5592_0;    relay_conn far_5_5592_0_a(.in(layer_4[22]), .out(far_5_5592_0[0]));    relay_conn far_5_5592_0_b(.in(layer_4[134]), .out(far_5_5592_0[1]));
    wire [1:0] far_5_5592_1;    relay_conn far_5_5592_1_a(.in(far_5_5592_0[0]), .out(far_5_5592_1[0]));    relay_conn far_5_5592_1_b(.in(far_5_5592_0[1]), .out(far_5_5592_1[1]));
    wire [1:0] far_5_5592_2;    relay_conn far_5_5592_2_a(.in(far_5_5592_1[0]), .out(far_5_5592_2[0]));    relay_conn far_5_5592_2_b(.in(far_5_5592_1[1]), .out(far_5_5592_2[1]));
    assign layer_5[492] = far_5_5592_2[1]; 
    assign layer_5[493] = layer_4[401] & ~layer_4[380]; 
    wire [1:0] far_5_5594_0;    relay_conn far_5_5594_0_a(.in(layer_4[790]), .out(far_5_5594_0[0]));    relay_conn far_5_5594_0_b(.in(layer_4[826]), .out(far_5_5594_0[1]));
    assign layer_5[494] = far_5_5594_0[1] & ~far_5_5594_0[0]; 
    wire [1:0] far_5_5595_0;    relay_conn far_5_5595_0_a(.in(layer_4[624]), .out(far_5_5595_0[0]));    relay_conn far_5_5595_0_b(.in(layer_4[745]), .out(far_5_5595_0[1]));
    wire [1:0] far_5_5595_1;    relay_conn far_5_5595_1_a(.in(far_5_5595_0[0]), .out(far_5_5595_1[0]));    relay_conn far_5_5595_1_b(.in(far_5_5595_0[1]), .out(far_5_5595_1[1]));
    wire [1:0] far_5_5595_2;    relay_conn far_5_5595_2_a(.in(far_5_5595_1[0]), .out(far_5_5595_2[0]));    relay_conn far_5_5595_2_b(.in(far_5_5595_1[1]), .out(far_5_5595_2[1]));
    assign layer_5[495] = far_5_5595_2[1] & ~far_5_5595_2[0]; 
    wire [1:0] far_5_5596_0;    relay_conn far_5_5596_0_a(.in(layer_4[931]), .out(far_5_5596_0[0]));    relay_conn far_5_5596_0_b(.in(layer_4[806]), .out(far_5_5596_0[1]));
    wire [1:0] far_5_5596_1;    relay_conn far_5_5596_1_a(.in(far_5_5596_0[0]), .out(far_5_5596_1[0]));    relay_conn far_5_5596_1_b(.in(far_5_5596_0[1]), .out(far_5_5596_1[1]));
    wire [1:0] far_5_5596_2;    relay_conn far_5_5596_2_a(.in(far_5_5596_1[0]), .out(far_5_5596_2[0]));    relay_conn far_5_5596_2_b(.in(far_5_5596_1[1]), .out(far_5_5596_2[1]));
    assign layer_5[496] = far_5_5596_2[1]; 
    assign layer_5[497] = ~layer_4[983] | (layer_4[997] & layer_4[983]); 
    wire [1:0] far_5_5598_0;    relay_conn far_5_5598_0_a(.in(layer_4[447]), .out(far_5_5598_0[0]));    relay_conn far_5_5598_0_b(.in(layer_4[363]), .out(far_5_5598_0[1]));
    wire [1:0] far_5_5598_1;    relay_conn far_5_5598_1_a(.in(far_5_5598_0[0]), .out(far_5_5598_1[0]));    relay_conn far_5_5598_1_b(.in(far_5_5598_0[1]), .out(far_5_5598_1[1]));
    assign layer_5[498] = far_5_5598_1[1]; 
    assign layer_5[499] = layer_4[208] & layer_4[191]; 
    wire [1:0] far_5_5600_0;    relay_conn far_5_5600_0_a(.in(layer_4[384]), .out(far_5_5600_0[0]));    relay_conn far_5_5600_0_b(.in(layer_4[454]), .out(far_5_5600_0[1]));
    wire [1:0] far_5_5600_1;    relay_conn far_5_5600_1_a(.in(far_5_5600_0[0]), .out(far_5_5600_1[0]));    relay_conn far_5_5600_1_b(.in(far_5_5600_0[1]), .out(far_5_5600_1[1]));
    assign layer_5[500] = ~far_5_5600_1[1]; 
    wire [1:0] far_5_5601_0;    relay_conn far_5_5601_0_a(.in(layer_4[293]), .out(far_5_5601_0[0]));    relay_conn far_5_5601_0_b(.in(layer_4[255]), .out(far_5_5601_0[1]));
    assign layer_5[501] = far_5_5601_0[0] & ~far_5_5601_0[1]; 
    assign layer_5[502] = layer_4[84]; 
    wire [1:0] far_5_5603_0;    relay_conn far_5_5603_0_a(.in(layer_4[614]), .out(far_5_5603_0[0]));    relay_conn far_5_5603_0_b(.in(layer_4[674]), .out(far_5_5603_0[1]));
    assign layer_5[503] = far_5_5603_0[0]; 
    wire [1:0] far_5_5604_0;    relay_conn far_5_5604_0_a(.in(layer_4[309]), .out(far_5_5604_0[0]));    relay_conn far_5_5604_0_b(.in(layer_4[192]), .out(far_5_5604_0[1]));
    wire [1:0] far_5_5604_1;    relay_conn far_5_5604_1_a(.in(far_5_5604_0[0]), .out(far_5_5604_1[0]));    relay_conn far_5_5604_1_b(.in(far_5_5604_0[1]), .out(far_5_5604_1[1]));
    wire [1:0] far_5_5604_2;    relay_conn far_5_5604_2_a(.in(far_5_5604_1[0]), .out(far_5_5604_2[0]));    relay_conn far_5_5604_2_b(.in(far_5_5604_1[1]), .out(far_5_5604_2[1]));
    assign layer_5[504] = far_5_5604_2[0] | far_5_5604_2[1]; 
    wire [1:0] far_5_5605_0;    relay_conn far_5_5605_0_a(.in(layer_4[559]), .out(far_5_5605_0[0]));    relay_conn far_5_5605_0_b(.in(layer_4[665]), .out(far_5_5605_0[1]));
    wire [1:0] far_5_5605_1;    relay_conn far_5_5605_1_a(.in(far_5_5605_0[0]), .out(far_5_5605_1[0]));    relay_conn far_5_5605_1_b(.in(far_5_5605_0[1]), .out(far_5_5605_1[1]));
    wire [1:0] far_5_5605_2;    relay_conn far_5_5605_2_a(.in(far_5_5605_1[0]), .out(far_5_5605_2[0]));    relay_conn far_5_5605_2_b(.in(far_5_5605_1[1]), .out(far_5_5605_2[1]));
    assign layer_5[505] = ~far_5_5605_2[1]; 
    wire [1:0] far_5_5606_0;    relay_conn far_5_5606_0_a(.in(layer_4[133]), .out(far_5_5606_0[0]));    relay_conn far_5_5606_0_b(.in(layer_4[28]), .out(far_5_5606_0[1]));
    wire [1:0] far_5_5606_1;    relay_conn far_5_5606_1_a(.in(far_5_5606_0[0]), .out(far_5_5606_1[0]));    relay_conn far_5_5606_1_b(.in(far_5_5606_0[1]), .out(far_5_5606_1[1]));
    wire [1:0] far_5_5606_2;    relay_conn far_5_5606_2_a(.in(far_5_5606_1[0]), .out(far_5_5606_2[0]));    relay_conn far_5_5606_2_b(.in(far_5_5606_1[1]), .out(far_5_5606_2[1]));
    assign layer_5[506] = far_5_5606_2[1]; 
    assign layer_5[507] = layer_4[692] & ~layer_4[684]; 
    wire [1:0] far_5_5608_0;    relay_conn far_5_5608_0_a(.in(layer_4[573]), .out(far_5_5608_0[0]));    relay_conn far_5_5608_0_b(.in(layer_4[674]), .out(far_5_5608_0[1]));
    wire [1:0] far_5_5608_1;    relay_conn far_5_5608_1_a(.in(far_5_5608_0[0]), .out(far_5_5608_1[0]));    relay_conn far_5_5608_1_b(.in(far_5_5608_0[1]), .out(far_5_5608_1[1]));
    wire [1:0] far_5_5608_2;    relay_conn far_5_5608_2_a(.in(far_5_5608_1[0]), .out(far_5_5608_2[0]));    relay_conn far_5_5608_2_b(.in(far_5_5608_1[1]), .out(far_5_5608_2[1]));
    assign layer_5[508] = far_5_5608_2[0]; 
    wire [1:0] far_5_5609_0;    relay_conn far_5_5609_0_a(.in(layer_4[740]), .out(far_5_5609_0[0]));    relay_conn far_5_5609_0_b(.in(layer_4[650]), .out(far_5_5609_0[1]));
    wire [1:0] far_5_5609_1;    relay_conn far_5_5609_1_a(.in(far_5_5609_0[0]), .out(far_5_5609_1[0]));    relay_conn far_5_5609_1_b(.in(far_5_5609_0[1]), .out(far_5_5609_1[1]));
    assign layer_5[509] = far_5_5609_1[0] | far_5_5609_1[1]; 
    wire [1:0] far_5_5610_0;    relay_conn far_5_5610_0_a(.in(layer_4[1013]), .out(far_5_5610_0[0]));    relay_conn far_5_5610_0_b(.in(layer_4[898]), .out(far_5_5610_0[1]));
    wire [1:0] far_5_5610_1;    relay_conn far_5_5610_1_a(.in(far_5_5610_0[0]), .out(far_5_5610_1[0]));    relay_conn far_5_5610_1_b(.in(far_5_5610_0[1]), .out(far_5_5610_1[1]));
    wire [1:0] far_5_5610_2;    relay_conn far_5_5610_2_a(.in(far_5_5610_1[0]), .out(far_5_5610_2[0]));    relay_conn far_5_5610_2_b(.in(far_5_5610_1[1]), .out(far_5_5610_2[1]));
    assign layer_5[510] = far_5_5610_2[1] & ~far_5_5610_2[0]; 
    assign layer_5[511] = ~layer_4[69]; 
    assign layer_5[512] = layer_4[318] | layer_4[293]; 
    wire [1:0] far_5_5613_0;    relay_conn far_5_5613_0_a(.in(layer_4[880]), .out(far_5_5613_0[0]));    relay_conn far_5_5613_0_b(.in(layer_4[959]), .out(far_5_5613_0[1]));
    wire [1:0] far_5_5613_1;    relay_conn far_5_5613_1_a(.in(far_5_5613_0[0]), .out(far_5_5613_1[0]));    relay_conn far_5_5613_1_b(.in(far_5_5613_0[1]), .out(far_5_5613_1[1]));
    assign layer_5[513] = far_5_5613_1[1]; 
    assign layer_5[514] = layer_4[627] & ~layer_4[645]; 
    wire [1:0] far_5_5615_0;    relay_conn far_5_5615_0_a(.in(layer_4[134]), .out(far_5_5615_0[0]));    relay_conn far_5_5615_0_b(.in(layer_4[102]), .out(far_5_5615_0[1]));
    assign layer_5[515] = ~far_5_5615_0[1] | (far_5_5615_0[0] & far_5_5615_0[1]); 
    wire [1:0] far_5_5616_0;    relay_conn far_5_5616_0_a(.in(layer_4[325]), .out(far_5_5616_0[0]));    relay_conn far_5_5616_0_b(.in(layer_4[443]), .out(far_5_5616_0[1]));
    wire [1:0] far_5_5616_1;    relay_conn far_5_5616_1_a(.in(far_5_5616_0[0]), .out(far_5_5616_1[0]));    relay_conn far_5_5616_1_b(.in(far_5_5616_0[1]), .out(far_5_5616_1[1]));
    wire [1:0] far_5_5616_2;    relay_conn far_5_5616_2_a(.in(far_5_5616_1[0]), .out(far_5_5616_2[0]));    relay_conn far_5_5616_2_b(.in(far_5_5616_1[1]), .out(far_5_5616_2[1]));
    assign layer_5[516] = ~far_5_5616_2[1]; 
    wire [1:0] far_5_5617_0;    relay_conn far_5_5617_0_a(.in(layer_4[500]), .out(far_5_5617_0[0]));    relay_conn far_5_5617_0_b(.in(layer_4[553]), .out(far_5_5617_0[1]));
    assign layer_5[517] = ~(far_5_5617_0[0] & far_5_5617_0[1]); 
    wire [1:0] far_5_5618_0;    relay_conn far_5_5618_0_a(.in(layer_4[526]), .out(far_5_5618_0[0]));    relay_conn far_5_5618_0_b(.in(layer_4[651]), .out(far_5_5618_0[1]));
    wire [1:0] far_5_5618_1;    relay_conn far_5_5618_1_a(.in(far_5_5618_0[0]), .out(far_5_5618_1[0]));    relay_conn far_5_5618_1_b(.in(far_5_5618_0[1]), .out(far_5_5618_1[1]));
    wire [1:0] far_5_5618_2;    relay_conn far_5_5618_2_a(.in(far_5_5618_1[0]), .out(far_5_5618_2[0]));    relay_conn far_5_5618_2_b(.in(far_5_5618_1[1]), .out(far_5_5618_2[1]));
    assign layer_5[518] = far_5_5618_2[1] & ~far_5_5618_2[0]; 
    wire [1:0] far_5_5619_0;    relay_conn far_5_5619_0_a(.in(layer_4[482]), .out(far_5_5619_0[0]));    relay_conn far_5_5619_0_b(.in(layer_4[545]), .out(far_5_5619_0[1]));
    assign layer_5[519] = ~(far_5_5619_0[0] & far_5_5619_0[1]); 
    wire [1:0] far_5_5620_0;    relay_conn far_5_5620_0_a(.in(layer_4[19]), .out(far_5_5620_0[0]));    relay_conn far_5_5620_0_b(.in(layer_4[131]), .out(far_5_5620_0[1]));
    wire [1:0] far_5_5620_1;    relay_conn far_5_5620_1_a(.in(far_5_5620_0[0]), .out(far_5_5620_1[0]));    relay_conn far_5_5620_1_b(.in(far_5_5620_0[1]), .out(far_5_5620_1[1]));
    wire [1:0] far_5_5620_2;    relay_conn far_5_5620_2_a(.in(far_5_5620_1[0]), .out(far_5_5620_2[0]));    relay_conn far_5_5620_2_b(.in(far_5_5620_1[1]), .out(far_5_5620_2[1]));
    assign layer_5[520] = far_5_5620_2[0] | far_5_5620_2[1]; 
    assign layer_5[521] = layer_4[88]; 
    wire [1:0] far_5_5622_0;    relay_conn far_5_5622_0_a(.in(layer_4[409]), .out(far_5_5622_0[0]));    relay_conn far_5_5622_0_b(.in(layer_4[294]), .out(far_5_5622_0[1]));
    wire [1:0] far_5_5622_1;    relay_conn far_5_5622_1_a(.in(far_5_5622_0[0]), .out(far_5_5622_1[0]));    relay_conn far_5_5622_1_b(.in(far_5_5622_0[1]), .out(far_5_5622_1[1]));
    wire [1:0] far_5_5622_2;    relay_conn far_5_5622_2_a(.in(far_5_5622_1[0]), .out(far_5_5622_2[0]));    relay_conn far_5_5622_2_b(.in(far_5_5622_1[1]), .out(far_5_5622_2[1]));
    assign layer_5[522] = ~far_5_5622_2[1]; 
    wire [1:0] far_5_5623_0;    relay_conn far_5_5623_0_a(.in(layer_4[277]), .out(far_5_5623_0[0]));    relay_conn far_5_5623_0_b(.in(layer_4[166]), .out(far_5_5623_0[1]));
    wire [1:0] far_5_5623_1;    relay_conn far_5_5623_1_a(.in(far_5_5623_0[0]), .out(far_5_5623_1[0]));    relay_conn far_5_5623_1_b(.in(far_5_5623_0[1]), .out(far_5_5623_1[1]));
    wire [1:0] far_5_5623_2;    relay_conn far_5_5623_2_a(.in(far_5_5623_1[0]), .out(far_5_5623_2[0]));    relay_conn far_5_5623_2_b(.in(far_5_5623_1[1]), .out(far_5_5623_2[1]));
    assign layer_5[523] = ~far_5_5623_2[0] | (far_5_5623_2[0] & far_5_5623_2[1]); 
    wire [1:0] far_5_5624_0;    relay_conn far_5_5624_0_a(.in(layer_4[656]), .out(far_5_5624_0[0]));    relay_conn far_5_5624_0_b(.in(layer_4[590]), .out(far_5_5624_0[1]));
    wire [1:0] far_5_5624_1;    relay_conn far_5_5624_1_a(.in(far_5_5624_0[0]), .out(far_5_5624_1[0]));    relay_conn far_5_5624_1_b(.in(far_5_5624_0[1]), .out(far_5_5624_1[1]));
    assign layer_5[524] = ~far_5_5624_1[1] | (far_5_5624_1[0] & far_5_5624_1[1]); 
    wire [1:0] far_5_5625_0;    relay_conn far_5_5625_0_a(.in(layer_4[850]), .out(far_5_5625_0[0]));    relay_conn far_5_5625_0_b(.in(layer_4[969]), .out(far_5_5625_0[1]));
    wire [1:0] far_5_5625_1;    relay_conn far_5_5625_1_a(.in(far_5_5625_0[0]), .out(far_5_5625_1[0]));    relay_conn far_5_5625_1_b(.in(far_5_5625_0[1]), .out(far_5_5625_1[1]));
    wire [1:0] far_5_5625_2;    relay_conn far_5_5625_2_a(.in(far_5_5625_1[0]), .out(far_5_5625_2[0]));    relay_conn far_5_5625_2_b(.in(far_5_5625_1[1]), .out(far_5_5625_2[1]));
    assign layer_5[525] = far_5_5625_2[1] & ~far_5_5625_2[0]; 
    wire [1:0] far_5_5626_0;    relay_conn far_5_5626_0_a(.in(layer_4[597]), .out(far_5_5626_0[0]));    relay_conn far_5_5626_0_b(.in(layer_4[485]), .out(far_5_5626_0[1]));
    wire [1:0] far_5_5626_1;    relay_conn far_5_5626_1_a(.in(far_5_5626_0[0]), .out(far_5_5626_1[0]));    relay_conn far_5_5626_1_b(.in(far_5_5626_0[1]), .out(far_5_5626_1[1]));
    wire [1:0] far_5_5626_2;    relay_conn far_5_5626_2_a(.in(far_5_5626_1[0]), .out(far_5_5626_2[0]));    relay_conn far_5_5626_2_b(.in(far_5_5626_1[1]), .out(far_5_5626_2[1]));
    assign layer_5[526] = ~(far_5_5626_2[0] | far_5_5626_2[1]); 
    assign layer_5[527] = ~(layer_4[884] | layer_4[885]); 
    wire [1:0] far_5_5628_0;    relay_conn far_5_5628_0_a(.in(layer_4[964]), .out(far_5_5628_0[0]));    relay_conn far_5_5628_0_b(.in(layer_4[894]), .out(far_5_5628_0[1]));
    wire [1:0] far_5_5628_1;    relay_conn far_5_5628_1_a(.in(far_5_5628_0[0]), .out(far_5_5628_1[0]));    relay_conn far_5_5628_1_b(.in(far_5_5628_0[1]), .out(far_5_5628_1[1]));
    assign layer_5[528] = ~far_5_5628_1[0]; 
    wire [1:0] far_5_5629_0;    relay_conn far_5_5629_0_a(.in(layer_4[718]), .out(far_5_5629_0[0]));    relay_conn far_5_5629_0_b(.in(layer_4[602]), .out(far_5_5629_0[1]));
    wire [1:0] far_5_5629_1;    relay_conn far_5_5629_1_a(.in(far_5_5629_0[0]), .out(far_5_5629_1[0]));    relay_conn far_5_5629_1_b(.in(far_5_5629_0[1]), .out(far_5_5629_1[1]));
    wire [1:0] far_5_5629_2;    relay_conn far_5_5629_2_a(.in(far_5_5629_1[0]), .out(far_5_5629_2[0]));    relay_conn far_5_5629_2_b(.in(far_5_5629_1[1]), .out(far_5_5629_2[1]));
    assign layer_5[529] = ~far_5_5629_2[0] | (far_5_5629_2[0] & far_5_5629_2[1]); 
    wire [1:0] far_5_5630_0;    relay_conn far_5_5630_0_a(.in(layer_4[754]), .out(far_5_5630_0[0]));    relay_conn far_5_5630_0_b(.in(layer_4[697]), .out(far_5_5630_0[1]));
    assign layer_5[530] = ~far_5_5630_0[1] | (far_5_5630_0[0] & far_5_5630_0[1]); 
    assign layer_5[531] = layer_4[773] ^ layer_4[751]; 
    wire [1:0] far_5_5632_0;    relay_conn far_5_5632_0_a(.in(layer_4[100]), .out(far_5_5632_0[0]));    relay_conn far_5_5632_0_b(.in(layer_4[43]), .out(far_5_5632_0[1]));
    assign layer_5[532] = far_5_5632_0[0] ^ far_5_5632_0[1]; 
    assign layer_5[533] = layer_4[895]; 
    wire [1:0] far_5_5634_0;    relay_conn far_5_5634_0_a(.in(layer_4[149]), .out(far_5_5634_0[0]));    relay_conn far_5_5634_0_b(.in(layer_4[117]), .out(far_5_5634_0[1]));
    assign layer_5[534] = far_5_5634_0[0] & far_5_5634_0[1]; 
    wire [1:0] far_5_5635_0;    relay_conn far_5_5635_0_a(.in(layer_4[89]), .out(far_5_5635_0[0]));    relay_conn far_5_5635_0_b(.in(layer_4[149]), .out(far_5_5635_0[1]));
    assign layer_5[535] = ~far_5_5635_0[0]; 
    wire [1:0] far_5_5636_0;    relay_conn far_5_5636_0_a(.in(layer_4[718]), .out(far_5_5636_0[0]));    relay_conn far_5_5636_0_b(.in(layer_4[608]), .out(far_5_5636_0[1]));
    wire [1:0] far_5_5636_1;    relay_conn far_5_5636_1_a(.in(far_5_5636_0[0]), .out(far_5_5636_1[0]));    relay_conn far_5_5636_1_b(.in(far_5_5636_0[1]), .out(far_5_5636_1[1]));
    wire [1:0] far_5_5636_2;    relay_conn far_5_5636_2_a(.in(far_5_5636_1[0]), .out(far_5_5636_2[0]));    relay_conn far_5_5636_2_b(.in(far_5_5636_1[1]), .out(far_5_5636_2[1]));
    assign layer_5[536] = far_5_5636_2[1]; 
    wire [1:0] far_5_5637_0;    relay_conn far_5_5637_0_a(.in(layer_4[333]), .out(far_5_5637_0[0]));    relay_conn far_5_5637_0_b(.in(layer_4[249]), .out(far_5_5637_0[1]));
    wire [1:0] far_5_5637_1;    relay_conn far_5_5637_1_a(.in(far_5_5637_0[0]), .out(far_5_5637_1[0]));    relay_conn far_5_5637_1_b(.in(far_5_5637_0[1]), .out(far_5_5637_1[1]));
    assign layer_5[537] = far_5_5637_1[1]; 
    wire [1:0] far_5_5638_0;    relay_conn far_5_5638_0_a(.in(layer_4[443]), .out(far_5_5638_0[0]));    relay_conn far_5_5638_0_b(.in(layer_4[349]), .out(far_5_5638_0[1]));
    wire [1:0] far_5_5638_1;    relay_conn far_5_5638_1_a(.in(far_5_5638_0[0]), .out(far_5_5638_1[0]));    relay_conn far_5_5638_1_b(.in(far_5_5638_0[1]), .out(far_5_5638_1[1]));
    assign layer_5[538] = far_5_5638_1[1] & ~far_5_5638_1[0]; 
    wire [1:0] far_5_5639_0;    relay_conn far_5_5639_0_a(.in(layer_4[574]), .out(far_5_5639_0[0]));    relay_conn far_5_5639_0_b(.in(layer_4[468]), .out(far_5_5639_0[1]));
    wire [1:0] far_5_5639_1;    relay_conn far_5_5639_1_a(.in(far_5_5639_0[0]), .out(far_5_5639_1[0]));    relay_conn far_5_5639_1_b(.in(far_5_5639_0[1]), .out(far_5_5639_1[1]));
    wire [1:0] far_5_5639_2;    relay_conn far_5_5639_2_a(.in(far_5_5639_1[0]), .out(far_5_5639_2[0]));    relay_conn far_5_5639_2_b(.in(far_5_5639_1[1]), .out(far_5_5639_2[1]));
    assign layer_5[539] = ~far_5_5639_2[0]; 
    wire [1:0] far_5_5640_0;    relay_conn far_5_5640_0_a(.in(layer_4[59]), .out(far_5_5640_0[0]));    relay_conn far_5_5640_0_b(.in(layer_4[129]), .out(far_5_5640_0[1]));
    wire [1:0] far_5_5640_1;    relay_conn far_5_5640_1_a(.in(far_5_5640_0[0]), .out(far_5_5640_1[0]));    relay_conn far_5_5640_1_b(.in(far_5_5640_0[1]), .out(far_5_5640_1[1]));
    assign layer_5[540] = far_5_5640_1[1] & ~far_5_5640_1[0]; 
    wire [1:0] far_5_5641_0;    relay_conn far_5_5641_0_a(.in(layer_4[642]), .out(far_5_5641_0[0]));    relay_conn far_5_5641_0_b(.in(layer_4[523]), .out(far_5_5641_0[1]));
    wire [1:0] far_5_5641_1;    relay_conn far_5_5641_1_a(.in(far_5_5641_0[0]), .out(far_5_5641_1[0]));    relay_conn far_5_5641_1_b(.in(far_5_5641_0[1]), .out(far_5_5641_1[1]));
    wire [1:0] far_5_5641_2;    relay_conn far_5_5641_2_a(.in(far_5_5641_1[0]), .out(far_5_5641_2[0]));    relay_conn far_5_5641_2_b(.in(far_5_5641_1[1]), .out(far_5_5641_2[1]));
    assign layer_5[541] = ~(far_5_5641_2[0] ^ far_5_5641_2[1]); 
    wire [1:0] far_5_5642_0;    relay_conn far_5_5642_0_a(.in(layer_4[200]), .out(far_5_5642_0[0]));    relay_conn far_5_5642_0_b(.in(layer_4[142]), .out(far_5_5642_0[1]));
    assign layer_5[542] = far_5_5642_0[0]; 
    wire [1:0] far_5_5643_0;    relay_conn far_5_5643_0_a(.in(layer_4[725]), .out(far_5_5643_0[0]));    relay_conn far_5_5643_0_b(.in(layer_4[617]), .out(far_5_5643_0[1]));
    wire [1:0] far_5_5643_1;    relay_conn far_5_5643_1_a(.in(far_5_5643_0[0]), .out(far_5_5643_1[0]));    relay_conn far_5_5643_1_b(.in(far_5_5643_0[1]), .out(far_5_5643_1[1]));
    wire [1:0] far_5_5643_2;    relay_conn far_5_5643_2_a(.in(far_5_5643_1[0]), .out(far_5_5643_2[0]));    relay_conn far_5_5643_2_b(.in(far_5_5643_1[1]), .out(far_5_5643_2[1]));
    assign layer_5[543] = far_5_5643_2[0]; 
    wire [1:0] far_5_5644_0;    relay_conn far_5_5644_0_a(.in(layer_4[646]), .out(far_5_5644_0[0]));    relay_conn far_5_5644_0_b(.in(layer_4[748]), .out(far_5_5644_0[1]));
    wire [1:0] far_5_5644_1;    relay_conn far_5_5644_1_a(.in(far_5_5644_0[0]), .out(far_5_5644_1[0]));    relay_conn far_5_5644_1_b(.in(far_5_5644_0[1]), .out(far_5_5644_1[1]));
    wire [1:0] far_5_5644_2;    relay_conn far_5_5644_2_a(.in(far_5_5644_1[0]), .out(far_5_5644_2[0]));    relay_conn far_5_5644_2_b(.in(far_5_5644_1[1]), .out(far_5_5644_2[1]));
    assign layer_5[544] = far_5_5644_2[1]; 
    wire [1:0] far_5_5645_0;    relay_conn far_5_5645_0_a(.in(layer_4[377]), .out(far_5_5645_0[0]));    relay_conn far_5_5645_0_b(.in(layer_4[423]), .out(far_5_5645_0[1]));
    assign layer_5[545] = far_5_5645_0[0]; 
    assign layer_5[546] = ~layer_4[282]; 
    wire [1:0] far_5_5647_0;    relay_conn far_5_5647_0_a(.in(layer_4[1006]), .out(far_5_5647_0[0]));    relay_conn far_5_5647_0_b(.in(layer_4[928]), .out(far_5_5647_0[1]));
    wire [1:0] far_5_5647_1;    relay_conn far_5_5647_1_a(.in(far_5_5647_0[0]), .out(far_5_5647_1[0]));    relay_conn far_5_5647_1_b(.in(far_5_5647_0[1]), .out(far_5_5647_1[1]));
    assign layer_5[547] = ~far_5_5647_1[0] | (far_5_5647_1[0] & far_5_5647_1[1]); 
    assign layer_5[548] = ~(layer_4[94] | layer_4[78]); 
    wire [1:0] far_5_5649_0;    relay_conn far_5_5649_0_a(.in(layer_4[870]), .out(far_5_5649_0[0]));    relay_conn far_5_5649_0_b(.in(layer_4[806]), .out(far_5_5649_0[1]));
    wire [1:0] far_5_5649_1;    relay_conn far_5_5649_1_a(.in(far_5_5649_0[0]), .out(far_5_5649_1[0]));    relay_conn far_5_5649_1_b(.in(far_5_5649_0[1]), .out(far_5_5649_1[1]));
    assign layer_5[549] = ~far_5_5649_1[0]; 
    wire [1:0] far_5_5650_0;    relay_conn far_5_5650_0_a(.in(layer_4[935]), .out(far_5_5650_0[0]));    relay_conn far_5_5650_0_b(.in(layer_4[902]), .out(far_5_5650_0[1]));
    assign layer_5[550] = far_5_5650_0[1] & ~far_5_5650_0[0]; 
    wire [1:0] far_5_5651_0;    relay_conn far_5_5651_0_a(.in(layer_4[545]), .out(far_5_5651_0[0]));    relay_conn far_5_5651_0_b(.in(layer_4[487]), .out(far_5_5651_0[1]));
    assign layer_5[551] = far_5_5651_0[0]; 
    wire [1:0] far_5_5652_0;    relay_conn far_5_5652_0_a(.in(layer_4[636]), .out(far_5_5652_0[0]));    relay_conn far_5_5652_0_b(.in(layer_4[571]), .out(far_5_5652_0[1]));
    wire [1:0] far_5_5652_1;    relay_conn far_5_5652_1_a(.in(far_5_5652_0[0]), .out(far_5_5652_1[0]));    relay_conn far_5_5652_1_b(.in(far_5_5652_0[1]), .out(far_5_5652_1[1]));
    assign layer_5[552] = ~(far_5_5652_1[0] | far_5_5652_1[1]); 
    wire [1:0] far_5_5653_0;    relay_conn far_5_5653_0_a(.in(layer_4[485]), .out(far_5_5653_0[0]));    relay_conn far_5_5653_0_b(.in(layer_4[554]), .out(far_5_5653_0[1]));
    wire [1:0] far_5_5653_1;    relay_conn far_5_5653_1_a(.in(far_5_5653_0[0]), .out(far_5_5653_1[0]));    relay_conn far_5_5653_1_b(.in(far_5_5653_0[1]), .out(far_5_5653_1[1]));
    assign layer_5[553] = ~far_5_5653_1[0]; 
    wire [1:0] far_5_5654_0;    relay_conn far_5_5654_0_a(.in(layer_4[754]), .out(far_5_5654_0[0]));    relay_conn far_5_5654_0_b(.in(layer_4[689]), .out(far_5_5654_0[1]));
    wire [1:0] far_5_5654_1;    relay_conn far_5_5654_1_a(.in(far_5_5654_0[0]), .out(far_5_5654_1[0]));    relay_conn far_5_5654_1_b(.in(far_5_5654_0[1]), .out(far_5_5654_1[1]));
    assign layer_5[554] = ~far_5_5654_1[1]; 
    wire [1:0] far_5_5655_0;    relay_conn far_5_5655_0_a(.in(layer_4[895]), .out(far_5_5655_0[0]));    relay_conn far_5_5655_0_b(.in(layer_4[1006]), .out(far_5_5655_0[1]));
    wire [1:0] far_5_5655_1;    relay_conn far_5_5655_1_a(.in(far_5_5655_0[0]), .out(far_5_5655_1[0]));    relay_conn far_5_5655_1_b(.in(far_5_5655_0[1]), .out(far_5_5655_1[1]));
    wire [1:0] far_5_5655_2;    relay_conn far_5_5655_2_a(.in(far_5_5655_1[0]), .out(far_5_5655_2[0]));    relay_conn far_5_5655_2_b(.in(far_5_5655_1[1]), .out(far_5_5655_2[1]));
    assign layer_5[555] = far_5_5655_2[0]; 
    wire [1:0] far_5_5656_0;    relay_conn far_5_5656_0_a(.in(layer_4[800]), .out(far_5_5656_0[0]));    relay_conn far_5_5656_0_b(.in(layer_4[675]), .out(far_5_5656_0[1]));
    wire [1:0] far_5_5656_1;    relay_conn far_5_5656_1_a(.in(far_5_5656_0[0]), .out(far_5_5656_1[0]));    relay_conn far_5_5656_1_b(.in(far_5_5656_0[1]), .out(far_5_5656_1[1]));
    wire [1:0] far_5_5656_2;    relay_conn far_5_5656_2_a(.in(far_5_5656_1[0]), .out(far_5_5656_2[0]));    relay_conn far_5_5656_2_b(.in(far_5_5656_1[1]), .out(far_5_5656_2[1]));
    assign layer_5[556] = far_5_5656_2[0]; 
    wire [1:0] far_5_5657_0;    relay_conn far_5_5657_0_a(.in(layer_4[79]), .out(far_5_5657_0[0]));    relay_conn far_5_5657_0_b(.in(layer_4[42]), .out(far_5_5657_0[1]));
    assign layer_5[557] = ~(far_5_5657_0[0] ^ far_5_5657_0[1]); 
    assign layer_5[558] = ~(layer_4[443] & layer_4[428]); 
    wire [1:0] far_5_5659_0;    relay_conn far_5_5659_0_a(.in(layer_4[875]), .out(far_5_5659_0[0]));    relay_conn far_5_5659_0_b(.in(layer_4[759]), .out(far_5_5659_0[1]));
    wire [1:0] far_5_5659_1;    relay_conn far_5_5659_1_a(.in(far_5_5659_0[0]), .out(far_5_5659_1[0]));    relay_conn far_5_5659_1_b(.in(far_5_5659_0[1]), .out(far_5_5659_1[1]));
    wire [1:0] far_5_5659_2;    relay_conn far_5_5659_2_a(.in(far_5_5659_1[0]), .out(far_5_5659_2[0]));    relay_conn far_5_5659_2_b(.in(far_5_5659_1[1]), .out(far_5_5659_2[1]));
    assign layer_5[559] = far_5_5659_2[0]; 
    assign layer_5[560] = layer_4[838] | layer_4[861]; 
    assign layer_5[561] = ~layer_4[102]; 
    wire [1:0] far_5_5662_0;    relay_conn far_5_5662_0_a(.in(layer_4[261]), .out(far_5_5662_0[0]));    relay_conn far_5_5662_0_b(.in(layer_4[369]), .out(far_5_5662_0[1]));
    wire [1:0] far_5_5662_1;    relay_conn far_5_5662_1_a(.in(far_5_5662_0[0]), .out(far_5_5662_1[0]));    relay_conn far_5_5662_1_b(.in(far_5_5662_0[1]), .out(far_5_5662_1[1]));
    wire [1:0] far_5_5662_2;    relay_conn far_5_5662_2_a(.in(far_5_5662_1[0]), .out(far_5_5662_2[0]));    relay_conn far_5_5662_2_b(.in(far_5_5662_1[1]), .out(far_5_5662_2[1]));
    assign layer_5[562] = ~far_5_5662_2[1] | (far_5_5662_2[0] & far_5_5662_2[1]); 
    wire [1:0] far_5_5663_0;    relay_conn far_5_5663_0_a(.in(layer_4[761]), .out(far_5_5663_0[0]));    relay_conn far_5_5663_0_b(.in(layer_4[886]), .out(far_5_5663_0[1]));
    wire [1:0] far_5_5663_1;    relay_conn far_5_5663_1_a(.in(far_5_5663_0[0]), .out(far_5_5663_1[0]));    relay_conn far_5_5663_1_b(.in(far_5_5663_0[1]), .out(far_5_5663_1[1]));
    wire [1:0] far_5_5663_2;    relay_conn far_5_5663_2_a(.in(far_5_5663_1[0]), .out(far_5_5663_2[0]));    relay_conn far_5_5663_2_b(.in(far_5_5663_1[1]), .out(far_5_5663_2[1]));
    assign layer_5[563] = ~far_5_5663_2[0] | (far_5_5663_2[0] & far_5_5663_2[1]); 
    assign layer_5[564] = layer_4[6] & ~layer_4[13]; 
    wire [1:0] far_5_5665_0;    relay_conn far_5_5665_0_a(.in(layer_4[71]), .out(far_5_5665_0[0]));    relay_conn far_5_5665_0_b(.in(layer_4[16]), .out(far_5_5665_0[1]));
    assign layer_5[565] = ~far_5_5665_0[1] | (far_5_5665_0[0] & far_5_5665_0[1]); 
    assign layer_5[566] = layer_4[444] & ~layer_4[443]; 
    assign layer_5[567] = ~(layer_4[517] & layer_4[538]); 
    wire [1:0] far_5_5668_0;    relay_conn far_5_5668_0_a(.in(layer_4[141]), .out(far_5_5668_0[0]));    relay_conn far_5_5668_0_b(.in(layer_4[18]), .out(far_5_5668_0[1]));
    wire [1:0] far_5_5668_1;    relay_conn far_5_5668_1_a(.in(far_5_5668_0[0]), .out(far_5_5668_1[0]));    relay_conn far_5_5668_1_b(.in(far_5_5668_0[1]), .out(far_5_5668_1[1]));
    wire [1:0] far_5_5668_2;    relay_conn far_5_5668_2_a(.in(far_5_5668_1[0]), .out(far_5_5668_2[0]));    relay_conn far_5_5668_2_b(.in(far_5_5668_1[1]), .out(far_5_5668_2[1]));
    assign layer_5[568] = ~far_5_5668_2[0]; 
    wire [1:0] far_5_5669_0;    relay_conn far_5_5669_0_a(.in(layer_4[482]), .out(far_5_5669_0[0]));    relay_conn far_5_5669_0_b(.in(layer_4[523]), .out(far_5_5669_0[1]));
    assign layer_5[569] = far_5_5669_0[0]; 
    wire [1:0] far_5_5670_0;    relay_conn far_5_5670_0_a(.in(layer_4[388]), .out(far_5_5670_0[0]));    relay_conn far_5_5670_0_b(.in(layer_4[266]), .out(far_5_5670_0[1]));
    wire [1:0] far_5_5670_1;    relay_conn far_5_5670_1_a(.in(far_5_5670_0[0]), .out(far_5_5670_1[0]));    relay_conn far_5_5670_1_b(.in(far_5_5670_0[1]), .out(far_5_5670_1[1]));
    wire [1:0] far_5_5670_2;    relay_conn far_5_5670_2_a(.in(far_5_5670_1[0]), .out(far_5_5670_2[0]));    relay_conn far_5_5670_2_b(.in(far_5_5670_1[1]), .out(far_5_5670_2[1]));
    assign layer_5[570] = far_5_5670_2[1]; 
    assign layer_5[571] = ~(layer_4[723] | layer_4[741]); 
    wire [1:0] far_5_5672_0;    relay_conn far_5_5672_0_a(.in(layer_4[146]), .out(far_5_5672_0[0]));    relay_conn far_5_5672_0_b(.in(layer_4[89]), .out(far_5_5672_0[1]));
    assign layer_5[572] = far_5_5672_0[0]; 
    wire [1:0] far_5_5673_0;    relay_conn far_5_5673_0_a(.in(layer_4[331]), .out(far_5_5673_0[0]));    relay_conn far_5_5673_0_b(.in(layer_4[382]), .out(far_5_5673_0[1]));
    assign layer_5[573] = far_5_5673_0[0] ^ far_5_5673_0[1]; 
    wire [1:0] far_5_5674_0;    relay_conn far_5_5674_0_a(.in(layer_4[850]), .out(far_5_5674_0[0]));    relay_conn far_5_5674_0_b(.in(layer_4[977]), .out(far_5_5674_0[1]));
    wire [1:0] far_5_5674_1;    relay_conn far_5_5674_1_a(.in(far_5_5674_0[0]), .out(far_5_5674_1[0]));    relay_conn far_5_5674_1_b(.in(far_5_5674_0[1]), .out(far_5_5674_1[1]));
    wire [1:0] far_5_5674_2;    relay_conn far_5_5674_2_a(.in(far_5_5674_1[0]), .out(far_5_5674_2[0]));    relay_conn far_5_5674_2_b(.in(far_5_5674_1[1]), .out(far_5_5674_2[1]));
    assign layer_5[574] = ~far_5_5674_2[0] | (far_5_5674_2[0] & far_5_5674_2[1]); 
    wire [1:0] far_5_5675_0;    relay_conn far_5_5675_0_a(.in(layer_4[472]), .out(far_5_5675_0[0]));    relay_conn far_5_5675_0_b(.in(layer_4[417]), .out(far_5_5675_0[1]));
    assign layer_5[575] = ~far_5_5675_0[1]; 
    wire [1:0] far_5_5676_0;    relay_conn far_5_5676_0_a(.in(layer_4[930]), .out(far_5_5676_0[0]));    relay_conn far_5_5676_0_b(.in(layer_4[876]), .out(far_5_5676_0[1]));
    assign layer_5[576] = far_5_5676_0[1]; 
    wire [1:0] far_5_5677_0;    relay_conn far_5_5677_0_a(.in(layer_4[553]), .out(far_5_5677_0[0]));    relay_conn far_5_5677_0_b(.in(layer_4[451]), .out(far_5_5677_0[1]));
    wire [1:0] far_5_5677_1;    relay_conn far_5_5677_1_a(.in(far_5_5677_0[0]), .out(far_5_5677_1[0]));    relay_conn far_5_5677_1_b(.in(far_5_5677_0[1]), .out(far_5_5677_1[1]));
    wire [1:0] far_5_5677_2;    relay_conn far_5_5677_2_a(.in(far_5_5677_1[0]), .out(far_5_5677_2[0]));    relay_conn far_5_5677_2_b(.in(far_5_5677_1[1]), .out(far_5_5677_2[1]));
    assign layer_5[577] = far_5_5677_2[0]; 
    wire [1:0] far_5_5678_0;    relay_conn far_5_5678_0_a(.in(layer_4[528]), .out(far_5_5678_0[0]));    relay_conn far_5_5678_0_b(.in(layer_4[590]), .out(far_5_5678_0[1]));
    assign layer_5[578] = ~far_5_5678_0[0]; 
    wire [1:0] far_5_5679_0;    relay_conn far_5_5679_0_a(.in(layer_4[577]), .out(far_5_5679_0[0]));    relay_conn far_5_5679_0_b(.in(layer_4[489]), .out(far_5_5679_0[1]));
    wire [1:0] far_5_5679_1;    relay_conn far_5_5679_1_a(.in(far_5_5679_0[0]), .out(far_5_5679_1[0]));    relay_conn far_5_5679_1_b(.in(far_5_5679_0[1]), .out(far_5_5679_1[1]));
    assign layer_5[579] = far_5_5679_1[0] | far_5_5679_1[1]; 
    wire [1:0] far_5_5680_0;    relay_conn far_5_5680_0_a(.in(layer_4[632]), .out(far_5_5680_0[0]));    relay_conn far_5_5680_0_b(.in(layer_4[547]), .out(far_5_5680_0[1]));
    wire [1:0] far_5_5680_1;    relay_conn far_5_5680_1_a(.in(far_5_5680_0[0]), .out(far_5_5680_1[0]));    relay_conn far_5_5680_1_b(.in(far_5_5680_0[1]), .out(far_5_5680_1[1]));
    assign layer_5[580] = far_5_5680_1[0] & ~far_5_5680_1[1]; 
    wire [1:0] far_5_5681_0;    relay_conn far_5_5681_0_a(.in(layer_4[222]), .out(far_5_5681_0[0]));    relay_conn far_5_5681_0_b(.in(layer_4[133]), .out(far_5_5681_0[1]));
    wire [1:0] far_5_5681_1;    relay_conn far_5_5681_1_a(.in(far_5_5681_0[0]), .out(far_5_5681_1[0]));    relay_conn far_5_5681_1_b(.in(far_5_5681_0[1]), .out(far_5_5681_1[1]));
    assign layer_5[581] = ~far_5_5681_1[0]; 
    wire [1:0] far_5_5682_0;    relay_conn far_5_5682_0_a(.in(layer_4[13]), .out(far_5_5682_0[0]));    relay_conn far_5_5682_0_b(.in(layer_4[86]), .out(far_5_5682_0[1]));
    wire [1:0] far_5_5682_1;    relay_conn far_5_5682_1_a(.in(far_5_5682_0[0]), .out(far_5_5682_1[0]));    relay_conn far_5_5682_1_b(.in(far_5_5682_0[1]), .out(far_5_5682_1[1]));
    assign layer_5[582] = ~far_5_5682_1[0]; 
    wire [1:0] far_5_5683_0;    relay_conn far_5_5683_0_a(.in(layer_4[483]), .out(far_5_5683_0[0]));    relay_conn far_5_5683_0_b(.in(layer_4[571]), .out(far_5_5683_0[1]));
    wire [1:0] far_5_5683_1;    relay_conn far_5_5683_1_a(.in(far_5_5683_0[0]), .out(far_5_5683_1[0]));    relay_conn far_5_5683_1_b(.in(far_5_5683_0[1]), .out(far_5_5683_1[1]));
    assign layer_5[583] = ~(far_5_5683_1[0] ^ far_5_5683_1[1]); 
    wire [1:0] far_5_5684_0;    relay_conn far_5_5684_0_a(.in(layer_4[608]), .out(far_5_5684_0[0]));    relay_conn far_5_5684_0_b(.in(layer_4[500]), .out(far_5_5684_0[1]));
    wire [1:0] far_5_5684_1;    relay_conn far_5_5684_1_a(.in(far_5_5684_0[0]), .out(far_5_5684_1[0]));    relay_conn far_5_5684_1_b(.in(far_5_5684_0[1]), .out(far_5_5684_1[1]));
    wire [1:0] far_5_5684_2;    relay_conn far_5_5684_2_a(.in(far_5_5684_1[0]), .out(far_5_5684_2[0]));    relay_conn far_5_5684_2_b(.in(far_5_5684_1[1]), .out(far_5_5684_2[1]));
    assign layer_5[584] = ~far_5_5684_2[1]; 
    wire [1:0] far_5_5685_0;    relay_conn far_5_5685_0_a(.in(layer_4[387]), .out(far_5_5685_0[0]));    relay_conn far_5_5685_0_b(.in(layer_4[472]), .out(far_5_5685_0[1]));
    wire [1:0] far_5_5685_1;    relay_conn far_5_5685_1_a(.in(far_5_5685_0[0]), .out(far_5_5685_1[0]));    relay_conn far_5_5685_1_b(.in(far_5_5685_0[1]), .out(far_5_5685_1[1]));
    assign layer_5[585] = ~(far_5_5685_1[0] & far_5_5685_1[1]); 
    wire [1:0] far_5_5686_0;    relay_conn far_5_5686_0_a(.in(layer_4[450]), .out(far_5_5686_0[0]));    relay_conn far_5_5686_0_b(.in(layer_4[514]), .out(far_5_5686_0[1]));
    wire [1:0] far_5_5686_1;    relay_conn far_5_5686_1_a(.in(far_5_5686_0[0]), .out(far_5_5686_1[0]));    relay_conn far_5_5686_1_b(.in(far_5_5686_0[1]), .out(far_5_5686_1[1]));
    assign layer_5[586] = far_5_5686_1[0] & ~far_5_5686_1[1]; 
    wire [1:0] far_5_5687_0;    relay_conn far_5_5687_0_a(.in(layer_4[945]), .out(far_5_5687_0[0]));    relay_conn far_5_5687_0_b(.in(layer_4[992]), .out(far_5_5687_0[1]));
    assign layer_5[587] = ~far_5_5687_0[0]; 
    assign layer_5[588] = ~layer_4[141]; 
    assign layer_5[589] = ~layer_4[45]; 
    assign layer_5[590] = layer_4[795] ^ layer_4[789]; 
    wire [1:0] far_5_5691_0;    relay_conn far_5_5691_0_a(.in(layer_4[386]), .out(far_5_5691_0[0]));    relay_conn far_5_5691_0_b(.in(layer_4[480]), .out(far_5_5691_0[1]));
    wire [1:0] far_5_5691_1;    relay_conn far_5_5691_1_a(.in(far_5_5691_0[0]), .out(far_5_5691_1[0]));    relay_conn far_5_5691_1_b(.in(far_5_5691_0[1]), .out(far_5_5691_1[1]));
    assign layer_5[591] = far_5_5691_1[0] & far_5_5691_1[1]; 
    wire [1:0] far_5_5692_0;    relay_conn far_5_5692_0_a(.in(layer_4[59]), .out(far_5_5692_0[0]));    relay_conn far_5_5692_0_b(.in(layer_4[124]), .out(far_5_5692_0[1]));
    wire [1:0] far_5_5692_1;    relay_conn far_5_5692_1_a(.in(far_5_5692_0[0]), .out(far_5_5692_1[0]));    relay_conn far_5_5692_1_b(.in(far_5_5692_0[1]), .out(far_5_5692_1[1]));
    assign layer_5[592] = ~(far_5_5692_1[0] | far_5_5692_1[1]); 
    wire [1:0] far_5_5693_0;    relay_conn far_5_5693_0_a(.in(layer_4[286]), .out(far_5_5693_0[0]));    relay_conn far_5_5693_0_b(.in(layer_4[188]), .out(far_5_5693_0[1]));
    wire [1:0] far_5_5693_1;    relay_conn far_5_5693_1_a(.in(far_5_5693_0[0]), .out(far_5_5693_1[0]));    relay_conn far_5_5693_1_b(.in(far_5_5693_0[1]), .out(far_5_5693_1[1]));
    wire [1:0] far_5_5693_2;    relay_conn far_5_5693_2_a(.in(far_5_5693_1[0]), .out(far_5_5693_2[0]));    relay_conn far_5_5693_2_b(.in(far_5_5693_1[1]), .out(far_5_5693_2[1]));
    assign layer_5[593] = ~(far_5_5693_2[0] | far_5_5693_2[1]); 
    wire [1:0] far_5_5694_0;    relay_conn far_5_5694_0_a(.in(layer_4[402]), .out(far_5_5694_0[0]));    relay_conn far_5_5694_0_b(.in(layer_4[288]), .out(far_5_5694_0[1]));
    wire [1:0] far_5_5694_1;    relay_conn far_5_5694_1_a(.in(far_5_5694_0[0]), .out(far_5_5694_1[0]));    relay_conn far_5_5694_1_b(.in(far_5_5694_0[1]), .out(far_5_5694_1[1]));
    wire [1:0] far_5_5694_2;    relay_conn far_5_5694_2_a(.in(far_5_5694_1[0]), .out(far_5_5694_2[0]));    relay_conn far_5_5694_2_b(.in(far_5_5694_1[1]), .out(far_5_5694_2[1]));
    assign layer_5[594] = ~(far_5_5694_2[0] | far_5_5694_2[1]); 
    wire [1:0] far_5_5695_0;    relay_conn far_5_5695_0_a(.in(layer_4[306]), .out(far_5_5695_0[0]));    relay_conn far_5_5695_0_b(.in(layer_4[224]), .out(far_5_5695_0[1]));
    wire [1:0] far_5_5695_1;    relay_conn far_5_5695_1_a(.in(far_5_5695_0[0]), .out(far_5_5695_1[0]));    relay_conn far_5_5695_1_b(.in(far_5_5695_0[1]), .out(far_5_5695_1[1]));
    assign layer_5[595] = ~(far_5_5695_1[0] & far_5_5695_1[1]); 
    assign layer_5[596] = ~(layer_4[642] | layer_4[661]); 
    wire [1:0] far_5_5697_0;    relay_conn far_5_5697_0_a(.in(layer_4[604]), .out(far_5_5697_0[0]));    relay_conn far_5_5697_0_b(.in(layer_4[678]), .out(far_5_5697_0[1]));
    wire [1:0] far_5_5697_1;    relay_conn far_5_5697_1_a(.in(far_5_5697_0[0]), .out(far_5_5697_1[0]));    relay_conn far_5_5697_1_b(.in(far_5_5697_0[1]), .out(far_5_5697_1[1]));
    assign layer_5[597] = far_5_5697_1[1] & ~far_5_5697_1[0]; 
    assign layer_5[598] = ~layer_4[864] | (layer_4[864] & layer_4[877]); 
    wire [1:0] far_5_5699_0;    relay_conn far_5_5699_0_a(.in(layer_4[45]), .out(far_5_5699_0[0]));    relay_conn far_5_5699_0_b(.in(layer_4[169]), .out(far_5_5699_0[1]));
    wire [1:0] far_5_5699_1;    relay_conn far_5_5699_1_a(.in(far_5_5699_0[0]), .out(far_5_5699_1[0]));    relay_conn far_5_5699_1_b(.in(far_5_5699_0[1]), .out(far_5_5699_1[1]));
    wire [1:0] far_5_5699_2;    relay_conn far_5_5699_2_a(.in(far_5_5699_1[0]), .out(far_5_5699_2[0]));    relay_conn far_5_5699_2_b(.in(far_5_5699_1[1]), .out(far_5_5699_2[1]));
    assign layer_5[599] = far_5_5699_2[0] & far_5_5699_2[1]; 
    wire [1:0] far_5_5700_0;    relay_conn far_5_5700_0_a(.in(layer_4[642]), .out(far_5_5700_0[0]));    relay_conn far_5_5700_0_b(.in(layer_4[675]), .out(far_5_5700_0[1]));
    assign layer_5[600] = ~far_5_5700_0[0]; 
    wire [1:0] far_5_5701_0;    relay_conn far_5_5701_0_a(.in(layer_4[754]), .out(far_5_5701_0[0]));    relay_conn far_5_5701_0_b(.in(layer_4[666]), .out(far_5_5701_0[1]));
    wire [1:0] far_5_5701_1;    relay_conn far_5_5701_1_a(.in(far_5_5701_0[0]), .out(far_5_5701_1[0]));    relay_conn far_5_5701_1_b(.in(far_5_5701_0[1]), .out(far_5_5701_1[1]));
    assign layer_5[601] = far_5_5701_1[0] | far_5_5701_1[1]; 
    assign layer_5[602] = ~layer_4[945]; 
    wire [1:0] far_5_5703_0;    relay_conn far_5_5703_0_a(.in(layer_4[910]), .out(far_5_5703_0[0]));    relay_conn far_5_5703_0_b(.in(layer_4[806]), .out(far_5_5703_0[1]));
    wire [1:0] far_5_5703_1;    relay_conn far_5_5703_1_a(.in(far_5_5703_0[0]), .out(far_5_5703_1[0]));    relay_conn far_5_5703_1_b(.in(far_5_5703_0[1]), .out(far_5_5703_1[1]));
    wire [1:0] far_5_5703_2;    relay_conn far_5_5703_2_a(.in(far_5_5703_1[0]), .out(far_5_5703_2[0]));    relay_conn far_5_5703_2_b(.in(far_5_5703_1[1]), .out(far_5_5703_2[1]));
    assign layer_5[603] = far_5_5703_2[1]; 
    wire [1:0] far_5_5704_0;    relay_conn far_5_5704_0_a(.in(layer_4[231]), .out(far_5_5704_0[0]));    relay_conn far_5_5704_0_b(.in(layer_4[186]), .out(far_5_5704_0[1]));
    assign layer_5[604] = far_5_5704_0[0] | far_5_5704_0[1]; 
    wire [1:0] far_5_5705_0;    relay_conn far_5_5705_0_a(.in(layer_4[545]), .out(far_5_5705_0[0]));    relay_conn far_5_5705_0_b(.in(layer_4[610]), .out(far_5_5705_0[1]));
    wire [1:0] far_5_5705_1;    relay_conn far_5_5705_1_a(.in(far_5_5705_0[0]), .out(far_5_5705_1[0]));    relay_conn far_5_5705_1_b(.in(far_5_5705_0[1]), .out(far_5_5705_1[1]));
    assign layer_5[605] = far_5_5705_1[0] | far_5_5705_1[1]; 
    wire [1:0] far_5_5706_0;    relay_conn far_5_5706_0_a(.in(layer_4[644]), .out(far_5_5706_0[0]));    relay_conn far_5_5706_0_b(.in(layer_4[608]), .out(far_5_5706_0[1]));
    assign layer_5[606] = far_5_5706_0[0] & ~far_5_5706_0[1]; 
    wire [1:0] far_5_5707_0;    relay_conn far_5_5707_0_a(.in(layer_4[876]), .out(far_5_5707_0[0]));    relay_conn far_5_5707_0_b(.in(layer_4[944]), .out(far_5_5707_0[1]));
    wire [1:0] far_5_5707_1;    relay_conn far_5_5707_1_a(.in(far_5_5707_0[0]), .out(far_5_5707_1[0]));    relay_conn far_5_5707_1_b(.in(far_5_5707_0[1]), .out(far_5_5707_1[1]));
    assign layer_5[607] = ~(far_5_5707_1[0] ^ far_5_5707_1[1]); 
    wire [1:0] far_5_5708_0;    relay_conn far_5_5708_0_a(.in(layer_4[285]), .out(far_5_5708_0[0]));    relay_conn far_5_5708_0_b(.in(layer_4[217]), .out(far_5_5708_0[1]));
    wire [1:0] far_5_5708_1;    relay_conn far_5_5708_1_a(.in(far_5_5708_0[0]), .out(far_5_5708_1[0]));    relay_conn far_5_5708_1_b(.in(far_5_5708_0[1]), .out(far_5_5708_1[1]));
    assign layer_5[608] = ~far_5_5708_1[0] | (far_5_5708_1[0] & far_5_5708_1[1]); 
    wire [1:0] far_5_5709_0;    relay_conn far_5_5709_0_a(.in(layer_4[181]), .out(far_5_5709_0[0]));    relay_conn far_5_5709_0_b(.in(layer_4[89]), .out(far_5_5709_0[1]));
    wire [1:0] far_5_5709_1;    relay_conn far_5_5709_1_a(.in(far_5_5709_0[0]), .out(far_5_5709_1[0]));    relay_conn far_5_5709_1_b(.in(far_5_5709_0[1]), .out(far_5_5709_1[1]));
    assign layer_5[609] = far_5_5709_1[0] | far_5_5709_1[1]; 
    assign layer_5[610] = layer_4[357] & ~layer_4[350]; 
    wire [1:0] far_5_5711_0;    relay_conn far_5_5711_0_a(.in(layer_4[521]), .out(far_5_5711_0[0]));    relay_conn far_5_5711_0_b(.in(layer_4[645]), .out(far_5_5711_0[1]));
    wire [1:0] far_5_5711_1;    relay_conn far_5_5711_1_a(.in(far_5_5711_0[0]), .out(far_5_5711_1[0]));    relay_conn far_5_5711_1_b(.in(far_5_5711_0[1]), .out(far_5_5711_1[1]));
    wire [1:0] far_5_5711_2;    relay_conn far_5_5711_2_a(.in(far_5_5711_1[0]), .out(far_5_5711_2[0]));    relay_conn far_5_5711_2_b(.in(far_5_5711_1[1]), .out(far_5_5711_2[1]));
    assign layer_5[611] = ~far_5_5711_2[1] | (far_5_5711_2[0] & far_5_5711_2[1]); 
    wire [1:0] far_5_5712_0;    relay_conn far_5_5712_0_a(.in(layer_4[130]), .out(far_5_5712_0[0]));    relay_conn far_5_5712_0_b(.in(layer_4[72]), .out(far_5_5712_0[1]));
    assign layer_5[612] = ~far_5_5712_0[1] | (far_5_5712_0[0] & far_5_5712_0[1]); 
    wire [1:0] far_5_5713_0;    relay_conn far_5_5713_0_a(.in(layer_4[363]), .out(far_5_5713_0[0]));    relay_conn far_5_5713_0_b(.in(layer_4[472]), .out(far_5_5713_0[1]));
    wire [1:0] far_5_5713_1;    relay_conn far_5_5713_1_a(.in(far_5_5713_0[0]), .out(far_5_5713_1[0]));    relay_conn far_5_5713_1_b(.in(far_5_5713_0[1]), .out(far_5_5713_1[1]));
    wire [1:0] far_5_5713_2;    relay_conn far_5_5713_2_a(.in(far_5_5713_1[0]), .out(far_5_5713_2[0]));    relay_conn far_5_5713_2_b(.in(far_5_5713_1[1]), .out(far_5_5713_2[1]));
    assign layer_5[613] = far_5_5713_2[0] & ~far_5_5713_2[1]; 
    assign layer_5[614] = ~layer_4[443]; 
    wire [1:0] far_5_5715_0;    relay_conn far_5_5715_0_a(.in(layer_4[149]), .out(far_5_5715_0[0]));    relay_conn far_5_5715_0_b(.in(layer_4[249]), .out(far_5_5715_0[1]));
    wire [1:0] far_5_5715_1;    relay_conn far_5_5715_1_a(.in(far_5_5715_0[0]), .out(far_5_5715_1[0]));    relay_conn far_5_5715_1_b(.in(far_5_5715_0[1]), .out(far_5_5715_1[1]));
    wire [1:0] far_5_5715_2;    relay_conn far_5_5715_2_a(.in(far_5_5715_1[0]), .out(far_5_5715_2[0]));    relay_conn far_5_5715_2_b(.in(far_5_5715_1[1]), .out(far_5_5715_2[1]));
    assign layer_5[615] = far_5_5715_2[1] & ~far_5_5715_2[0]; 
    wire [1:0] far_5_5716_0;    relay_conn far_5_5716_0_a(.in(layer_4[806]), .out(far_5_5716_0[0]));    relay_conn far_5_5716_0_b(.in(layer_4[861]), .out(far_5_5716_0[1]));
    assign layer_5[616] = ~far_5_5716_0[0] | (far_5_5716_0[0] & far_5_5716_0[1]); 
    wire [1:0] far_5_5717_0;    relay_conn far_5_5717_0_a(.in(layer_4[982]), .out(far_5_5717_0[0]));    relay_conn far_5_5717_0_b(.in(layer_4[867]), .out(far_5_5717_0[1]));
    wire [1:0] far_5_5717_1;    relay_conn far_5_5717_1_a(.in(far_5_5717_0[0]), .out(far_5_5717_1[0]));    relay_conn far_5_5717_1_b(.in(far_5_5717_0[1]), .out(far_5_5717_1[1]));
    wire [1:0] far_5_5717_2;    relay_conn far_5_5717_2_a(.in(far_5_5717_1[0]), .out(far_5_5717_2[0]));    relay_conn far_5_5717_2_b(.in(far_5_5717_1[1]), .out(far_5_5717_2[1]));
    assign layer_5[617] = ~(far_5_5717_2[0] ^ far_5_5717_2[1]); 
    wire [1:0] far_5_5718_0;    relay_conn far_5_5718_0_a(.in(layer_4[315]), .out(far_5_5718_0[0]));    relay_conn far_5_5718_0_b(.in(layer_4[383]), .out(far_5_5718_0[1]));
    wire [1:0] far_5_5718_1;    relay_conn far_5_5718_1_a(.in(far_5_5718_0[0]), .out(far_5_5718_1[0]));    relay_conn far_5_5718_1_b(.in(far_5_5718_0[1]), .out(far_5_5718_1[1]));
    assign layer_5[618] = ~(far_5_5718_1[0] & far_5_5718_1[1]); 
    wire [1:0] far_5_5719_0;    relay_conn far_5_5719_0_a(.in(layer_4[884]), .out(far_5_5719_0[0]));    relay_conn far_5_5719_0_b(.in(layer_4[975]), .out(far_5_5719_0[1]));
    wire [1:0] far_5_5719_1;    relay_conn far_5_5719_1_a(.in(far_5_5719_0[0]), .out(far_5_5719_1[0]));    relay_conn far_5_5719_1_b(.in(far_5_5719_0[1]), .out(far_5_5719_1[1]));
    assign layer_5[619] = ~(far_5_5719_1[0] | far_5_5719_1[1]); 
    wire [1:0] far_5_5720_0;    relay_conn far_5_5720_0_a(.in(layer_4[958]), .out(far_5_5720_0[0]));    relay_conn far_5_5720_0_b(.in(layer_4[838]), .out(far_5_5720_0[1]));
    wire [1:0] far_5_5720_1;    relay_conn far_5_5720_1_a(.in(far_5_5720_0[0]), .out(far_5_5720_1[0]));    relay_conn far_5_5720_1_b(.in(far_5_5720_0[1]), .out(far_5_5720_1[1]));
    wire [1:0] far_5_5720_2;    relay_conn far_5_5720_2_a(.in(far_5_5720_1[0]), .out(far_5_5720_2[0]));    relay_conn far_5_5720_2_b(.in(far_5_5720_1[1]), .out(far_5_5720_2[1]));
    assign layer_5[620] = far_5_5720_2[0]; 
    wire [1:0] far_5_5721_0;    relay_conn far_5_5721_0_a(.in(layer_4[103]), .out(far_5_5721_0[0]));    relay_conn far_5_5721_0_b(.in(layer_4[12]), .out(far_5_5721_0[1]));
    wire [1:0] far_5_5721_1;    relay_conn far_5_5721_1_a(.in(far_5_5721_0[0]), .out(far_5_5721_1[0]));    relay_conn far_5_5721_1_b(.in(far_5_5721_0[1]), .out(far_5_5721_1[1]));
    assign layer_5[621] = ~far_5_5721_1[0]; 
    assign layer_5[622] = ~layer_4[886]; 
    wire [1:0] far_5_5723_0;    relay_conn far_5_5723_0_a(.in(layer_4[541]), .out(far_5_5723_0[0]));    relay_conn far_5_5723_0_b(.in(layer_4[602]), .out(far_5_5723_0[1]));
    assign layer_5[623] = ~(far_5_5723_0[0] | far_5_5723_0[1]); 
    wire [1:0] far_5_5724_0;    relay_conn far_5_5724_0_a(.in(layer_4[759]), .out(far_5_5724_0[0]));    relay_conn far_5_5724_0_b(.in(layer_4[644]), .out(far_5_5724_0[1]));
    wire [1:0] far_5_5724_1;    relay_conn far_5_5724_1_a(.in(far_5_5724_0[0]), .out(far_5_5724_1[0]));    relay_conn far_5_5724_1_b(.in(far_5_5724_0[1]), .out(far_5_5724_1[1]));
    wire [1:0] far_5_5724_2;    relay_conn far_5_5724_2_a(.in(far_5_5724_1[0]), .out(far_5_5724_2[0]));    relay_conn far_5_5724_2_b(.in(far_5_5724_1[1]), .out(far_5_5724_2[1]));
    assign layer_5[624] = ~far_5_5724_2[1]; 
    wire [1:0] far_5_5725_0;    relay_conn far_5_5725_0_a(.in(layer_4[185]), .out(far_5_5725_0[0]));    relay_conn far_5_5725_0_b(.in(layer_4[298]), .out(far_5_5725_0[1]));
    wire [1:0] far_5_5725_1;    relay_conn far_5_5725_1_a(.in(far_5_5725_0[0]), .out(far_5_5725_1[0]));    relay_conn far_5_5725_1_b(.in(far_5_5725_0[1]), .out(far_5_5725_1[1]));
    wire [1:0] far_5_5725_2;    relay_conn far_5_5725_2_a(.in(far_5_5725_1[0]), .out(far_5_5725_2[0]));    relay_conn far_5_5725_2_b(.in(far_5_5725_1[1]), .out(far_5_5725_2[1]));
    assign layer_5[625] = far_5_5725_2[0] & ~far_5_5725_2[1]; 
    assign layer_5[626] = layer_4[730] & layer_4[728]; 
    wire [1:0] far_5_5727_0;    relay_conn far_5_5727_0_a(.in(layer_4[62]), .out(far_5_5727_0[0]));    relay_conn far_5_5727_0_b(.in(layer_4[115]), .out(far_5_5727_0[1]));
    assign layer_5[627] = ~far_5_5727_0[0]; 
    assign layer_5[628] = layer_4[905] & layer_4[931]; 
    wire [1:0] far_5_5729_0;    relay_conn far_5_5729_0_a(.in(layer_4[408]), .out(far_5_5729_0[0]));    relay_conn far_5_5729_0_b(.in(layer_4[323]), .out(far_5_5729_0[1]));
    wire [1:0] far_5_5729_1;    relay_conn far_5_5729_1_a(.in(far_5_5729_0[0]), .out(far_5_5729_1[0]));    relay_conn far_5_5729_1_b(.in(far_5_5729_0[1]), .out(far_5_5729_1[1]));
    assign layer_5[629] = ~far_5_5729_1[0]; 
    wire [1:0] far_5_5730_0;    relay_conn far_5_5730_0_a(.in(layer_4[983]), .out(far_5_5730_0[0]));    relay_conn far_5_5730_0_b(.in(layer_4[882]), .out(far_5_5730_0[1]));
    wire [1:0] far_5_5730_1;    relay_conn far_5_5730_1_a(.in(far_5_5730_0[0]), .out(far_5_5730_1[0]));    relay_conn far_5_5730_1_b(.in(far_5_5730_0[1]), .out(far_5_5730_1[1]));
    wire [1:0] far_5_5730_2;    relay_conn far_5_5730_2_a(.in(far_5_5730_1[0]), .out(far_5_5730_2[0]));    relay_conn far_5_5730_2_b(.in(far_5_5730_1[1]), .out(far_5_5730_2[1]));
    assign layer_5[630] = ~far_5_5730_2[1] | (far_5_5730_2[0] & far_5_5730_2[1]); 
    wire [1:0] far_5_5731_0;    relay_conn far_5_5731_0_a(.in(layer_4[327]), .out(far_5_5731_0[0]));    relay_conn far_5_5731_0_b(.in(layer_4[379]), .out(far_5_5731_0[1]));
    assign layer_5[631] = far_5_5731_0[1]; 
    wire [1:0] far_5_5732_0;    relay_conn far_5_5732_0_a(.in(layer_4[185]), .out(far_5_5732_0[0]));    relay_conn far_5_5732_0_b(.in(layer_4[279]), .out(far_5_5732_0[1]));
    wire [1:0] far_5_5732_1;    relay_conn far_5_5732_1_a(.in(far_5_5732_0[0]), .out(far_5_5732_1[0]));    relay_conn far_5_5732_1_b(.in(far_5_5732_0[1]), .out(far_5_5732_1[1]));
    assign layer_5[632] = ~far_5_5732_1[0]; 
    assign layer_5[633] = ~layer_4[13] | (layer_4[13] & layer_4[20]); 
    wire [1:0] far_5_5734_0;    relay_conn far_5_5734_0_a(.in(layer_4[536]), .out(far_5_5734_0[0]));    relay_conn far_5_5734_0_b(.in(layer_4[428]), .out(far_5_5734_0[1]));
    wire [1:0] far_5_5734_1;    relay_conn far_5_5734_1_a(.in(far_5_5734_0[0]), .out(far_5_5734_1[0]));    relay_conn far_5_5734_1_b(.in(far_5_5734_0[1]), .out(far_5_5734_1[1]));
    wire [1:0] far_5_5734_2;    relay_conn far_5_5734_2_a(.in(far_5_5734_1[0]), .out(far_5_5734_2[0]));    relay_conn far_5_5734_2_b(.in(far_5_5734_1[1]), .out(far_5_5734_2[1]));
    assign layer_5[634] = far_5_5734_2[0] | far_5_5734_2[1]; 
    wire [1:0] far_5_5735_0;    relay_conn far_5_5735_0_a(.in(layer_4[654]), .out(far_5_5735_0[0]));    relay_conn far_5_5735_0_b(.in(layer_4[569]), .out(far_5_5735_0[1]));
    wire [1:0] far_5_5735_1;    relay_conn far_5_5735_1_a(.in(far_5_5735_0[0]), .out(far_5_5735_1[0]));    relay_conn far_5_5735_1_b(.in(far_5_5735_0[1]), .out(far_5_5735_1[1]));
    assign layer_5[635] = ~(far_5_5735_1[0] ^ far_5_5735_1[1]); 
    wire [1:0] far_5_5736_0;    relay_conn far_5_5736_0_a(.in(layer_4[775]), .out(far_5_5736_0[0]));    relay_conn far_5_5736_0_b(.in(layer_4[884]), .out(far_5_5736_0[1]));
    wire [1:0] far_5_5736_1;    relay_conn far_5_5736_1_a(.in(far_5_5736_0[0]), .out(far_5_5736_1[0]));    relay_conn far_5_5736_1_b(.in(far_5_5736_0[1]), .out(far_5_5736_1[1]));
    wire [1:0] far_5_5736_2;    relay_conn far_5_5736_2_a(.in(far_5_5736_1[0]), .out(far_5_5736_2[0]));    relay_conn far_5_5736_2_b(.in(far_5_5736_1[1]), .out(far_5_5736_2[1]));
    assign layer_5[636] = ~far_5_5736_2[0]; 
    wire [1:0] far_5_5737_0;    relay_conn far_5_5737_0_a(.in(layer_4[855]), .out(far_5_5737_0[0]));    relay_conn far_5_5737_0_b(.in(layer_4[795]), .out(far_5_5737_0[1]));
    assign layer_5[637] = ~far_5_5737_0[0]; 
    assign layer_5[638] = layer_4[655] ^ layer_4[650]; 
    assign layer_5[639] = layer_4[167]; 
    wire [1:0] far_5_5740_0;    relay_conn far_5_5740_0_a(.in(layer_4[11]), .out(far_5_5740_0[0]));    relay_conn far_5_5740_0_b(.in(layer_4[45]), .out(far_5_5740_0[1]));
    assign layer_5[640] = far_5_5740_0[0]; 
    wire [1:0] far_5_5741_0;    relay_conn far_5_5741_0_a(.in(layer_4[991]), .out(far_5_5741_0[0]));    relay_conn far_5_5741_0_b(.in(layer_4[919]), .out(far_5_5741_0[1]));
    wire [1:0] far_5_5741_1;    relay_conn far_5_5741_1_a(.in(far_5_5741_0[0]), .out(far_5_5741_1[0]));    relay_conn far_5_5741_1_b(.in(far_5_5741_0[1]), .out(far_5_5741_1[1]));
    assign layer_5[641] = ~far_5_5741_1[1] | (far_5_5741_1[0] & far_5_5741_1[1]); 
    wire [1:0] far_5_5742_0;    relay_conn far_5_5742_0_a(.in(layer_4[221]), .out(far_5_5742_0[0]));    relay_conn far_5_5742_0_b(.in(layer_4[150]), .out(far_5_5742_0[1]));
    wire [1:0] far_5_5742_1;    relay_conn far_5_5742_1_a(.in(far_5_5742_0[0]), .out(far_5_5742_1[0]));    relay_conn far_5_5742_1_b(.in(far_5_5742_0[1]), .out(far_5_5742_1[1]));
    assign layer_5[642] = far_5_5742_1[1]; 
    wire [1:0] far_5_5743_0;    relay_conn far_5_5743_0_a(.in(layer_4[114]), .out(far_5_5743_0[0]));    relay_conn far_5_5743_0_b(.in(layer_4[188]), .out(far_5_5743_0[1]));
    wire [1:0] far_5_5743_1;    relay_conn far_5_5743_1_a(.in(far_5_5743_0[0]), .out(far_5_5743_1[0]));    relay_conn far_5_5743_1_b(.in(far_5_5743_0[1]), .out(far_5_5743_1[1]));
    assign layer_5[643] = far_5_5743_1[0] | far_5_5743_1[1]; 
    assign layer_5[644] = ~layer_4[88]; 
    assign layer_5[645] = layer_4[62] & ~layer_4[68]; 
    wire [1:0] far_5_5746_0;    relay_conn far_5_5746_0_a(.in(layer_4[929]), .out(far_5_5746_0[0]));    relay_conn far_5_5746_0_b(.in(layer_4[1013]), .out(far_5_5746_0[1]));
    wire [1:0] far_5_5746_1;    relay_conn far_5_5746_1_a(.in(far_5_5746_0[0]), .out(far_5_5746_1[0]));    relay_conn far_5_5746_1_b(.in(far_5_5746_0[1]), .out(far_5_5746_1[1]));
    assign layer_5[646] = far_5_5746_1[0] & far_5_5746_1[1]; 
    wire [1:0] far_5_5747_0;    relay_conn far_5_5747_0_a(.in(layer_4[759]), .out(far_5_5747_0[0]));    relay_conn far_5_5747_0_b(.in(layer_4[652]), .out(far_5_5747_0[1]));
    wire [1:0] far_5_5747_1;    relay_conn far_5_5747_1_a(.in(far_5_5747_0[0]), .out(far_5_5747_1[0]));    relay_conn far_5_5747_1_b(.in(far_5_5747_0[1]), .out(far_5_5747_1[1]));
    wire [1:0] far_5_5747_2;    relay_conn far_5_5747_2_a(.in(far_5_5747_1[0]), .out(far_5_5747_2[0]));    relay_conn far_5_5747_2_b(.in(far_5_5747_1[1]), .out(far_5_5747_2[1]));
    assign layer_5[647] = far_5_5747_2[0] ^ far_5_5747_2[1]; 
    wire [1:0] far_5_5748_0;    relay_conn far_5_5748_0_a(.in(layer_4[325]), .out(far_5_5748_0[0]));    relay_conn far_5_5748_0_b(.in(layer_4[223]), .out(far_5_5748_0[1]));
    wire [1:0] far_5_5748_1;    relay_conn far_5_5748_1_a(.in(far_5_5748_0[0]), .out(far_5_5748_1[0]));    relay_conn far_5_5748_1_b(.in(far_5_5748_0[1]), .out(far_5_5748_1[1]));
    wire [1:0] far_5_5748_2;    relay_conn far_5_5748_2_a(.in(far_5_5748_1[0]), .out(far_5_5748_2[0]));    relay_conn far_5_5748_2_b(.in(far_5_5748_1[1]), .out(far_5_5748_2[1]));
    assign layer_5[648] = ~far_5_5748_2[0]; 
    assign layer_5[649] = ~layer_4[757]; 
    wire [1:0] far_5_5750_0;    relay_conn far_5_5750_0_a(.in(layer_4[992]), .out(far_5_5750_0[0]));    relay_conn far_5_5750_0_b(.in(layer_4[951]), .out(far_5_5750_0[1]));
    assign layer_5[650] = ~far_5_5750_0[1] | (far_5_5750_0[0] & far_5_5750_0[1]); 
    wire [1:0] far_5_5751_0;    relay_conn far_5_5751_0_a(.in(layer_4[608]), .out(far_5_5751_0[0]));    relay_conn far_5_5751_0_b(.in(layer_4[556]), .out(far_5_5751_0[1]));
    assign layer_5[651] = ~far_5_5751_0[0]; 
    wire [1:0] far_5_5752_0;    relay_conn far_5_5752_0_a(.in(layer_4[515]), .out(far_5_5752_0[0]));    relay_conn far_5_5752_0_b(.in(layer_4[596]), .out(far_5_5752_0[1]));
    wire [1:0] far_5_5752_1;    relay_conn far_5_5752_1_a(.in(far_5_5752_0[0]), .out(far_5_5752_1[0]));    relay_conn far_5_5752_1_b(.in(far_5_5752_0[1]), .out(far_5_5752_1[1]));
    assign layer_5[652] = ~(far_5_5752_1[0] ^ far_5_5752_1[1]); 
    wire [1:0] far_5_5753_0;    relay_conn far_5_5753_0_a(.in(layer_4[802]), .out(far_5_5753_0[0]));    relay_conn far_5_5753_0_b(.in(layer_4[890]), .out(far_5_5753_0[1]));
    wire [1:0] far_5_5753_1;    relay_conn far_5_5753_1_a(.in(far_5_5753_0[0]), .out(far_5_5753_1[0]));    relay_conn far_5_5753_1_b(.in(far_5_5753_0[1]), .out(far_5_5753_1[1]));
    assign layer_5[653] = far_5_5753_1[1] & ~far_5_5753_1[0]; 
    wire [1:0] far_5_5754_0;    relay_conn far_5_5754_0_a(.in(layer_4[464]), .out(far_5_5754_0[0]));    relay_conn far_5_5754_0_b(.in(layer_4[567]), .out(far_5_5754_0[1]));
    wire [1:0] far_5_5754_1;    relay_conn far_5_5754_1_a(.in(far_5_5754_0[0]), .out(far_5_5754_1[0]));    relay_conn far_5_5754_1_b(.in(far_5_5754_0[1]), .out(far_5_5754_1[1]));
    wire [1:0] far_5_5754_2;    relay_conn far_5_5754_2_a(.in(far_5_5754_1[0]), .out(far_5_5754_2[0]));    relay_conn far_5_5754_2_b(.in(far_5_5754_1[1]), .out(far_5_5754_2[1]));
    assign layer_5[654] = ~far_5_5754_2[0] | (far_5_5754_2[0] & far_5_5754_2[1]); 
    wire [1:0] far_5_5755_0;    relay_conn far_5_5755_0_a(.in(layer_4[94]), .out(far_5_5755_0[0]));    relay_conn far_5_5755_0_b(.in(layer_4[166]), .out(far_5_5755_0[1]));
    wire [1:0] far_5_5755_1;    relay_conn far_5_5755_1_a(.in(far_5_5755_0[0]), .out(far_5_5755_1[0]));    relay_conn far_5_5755_1_b(.in(far_5_5755_0[1]), .out(far_5_5755_1[1]));
    assign layer_5[655] = far_5_5755_1[1] & ~far_5_5755_1[0]; 
    wire [1:0] far_5_5756_0;    relay_conn far_5_5756_0_a(.in(layer_4[428]), .out(far_5_5756_0[0]));    relay_conn far_5_5756_0_b(.in(layer_4[553]), .out(far_5_5756_0[1]));
    wire [1:0] far_5_5756_1;    relay_conn far_5_5756_1_a(.in(far_5_5756_0[0]), .out(far_5_5756_1[0]));    relay_conn far_5_5756_1_b(.in(far_5_5756_0[1]), .out(far_5_5756_1[1]));
    wire [1:0] far_5_5756_2;    relay_conn far_5_5756_2_a(.in(far_5_5756_1[0]), .out(far_5_5756_2[0]));    relay_conn far_5_5756_2_b(.in(far_5_5756_1[1]), .out(far_5_5756_2[1]));
    assign layer_5[656] = far_5_5756_2[1]; 
    assign layer_5[657] = ~layer_4[1005] | (layer_4[997] & layer_4[1005]); 
    wire [1:0] far_5_5758_0;    relay_conn far_5_5758_0_a(.in(layer_4[730]), .out(far_5_5758_0[0]));    relay_conn far_5_5758_0_b(.in(layer_4[629]), .out(far_5_5758_0[1]));
    wire [1:0] far_5_5758_1;    relay_conn far_5_5758_1_a(.in(far_5_5758_0[0]), .out(far_5_5758_1[0]));    relay_conn far_5_5758_1_b(.in(far_5_5758_0[1]), .out(far_5_5758_1[1]));
    wire [1:0] far_5_5758_2;    relay_conn far_5_5758_2_a(.in(far_5_5758_1[0]), .out(far_5_5758_2[0]));    relay_conn far_5_5758_2_b(.in(far_5_5758_1[1]), .out(far_5_5758_2[1]));
    assign layer_5[658] = ~(far_5_5758_2[0] | far_5_5758_2[1]); 
    wire [1:0] far_5_5759_0;    relay_conn far_5_5759_0_a(.in(layer_4[830]), .out(far_5_5759_0[0]));    relay_conn far_5_5759_0_b(.in(layer_4[876]), .out(far_5_5759_0[1]));
    assign layer_5[659] = ~far_5_5759_0[1] | (far_5_5759_0[0] & far_5_5759_0[1]); 
    assign layer_5[660] = layer_4[859] & layer_4[858]; 
    wire [1:0] far_5_5761_0;    relay_conn far_5_5761_0_a(.in(layer_4[92]), .out(far_5_5761_0[0]));    relay_conn far_5_5761_0_b(.in(layer_4[168]), .out(far_5_5761_0[1]));
    wire [1:0] far_5_5761_1;    relay_conn far_5_5761_1_a(.in(far_5_5761_0[0]), .out(far_5_5761_1[0]));    relay_conn far_5_5761_1_b(.in(far_5_5761_0[1]), .out(far_5_5761_1[1]));
    assign layer_5[661] = ~(far_5_5761_1[0] & far_5_5761_1[1]); 
    wire [1:0] far_5_5762_0;    relay_conn far_5_5762_0_a(.in(layer_4[424]), .out(far_5_5762_0[0]));    relay_conn far_5_5762_0_b(.in(layer_4[383]), .out(far_5_5762_0[1]));
    assign layer_5[662] = far_5_5762_0[1]; 
    wire [1:0] far_5_5763_0;    relay_conn far_5_5763_0_a(.in(layer_4[171]), .out(far_5_5763_0[0]));    relay_conn far_5_5763_0_b(.in(layer_4[114]), .out(far_5_5763_0[1]));
    assign layer_5[663] = ~(far_5_5763_0[0] & far_5_5763_0[1]); 
    assign layer_5[664] = layer_4[424] & ~layer_4[438]; 
    wire [1:0] far_5_5765_0;    relay_conn far_5_5765_0_a(.in(layer_4[202]), .out(far_5_5765_0[0]));    relay_conn far_5_5765_0_b(.in(layer_4[130]), .out(far_5_5765_0[1]));
    wire [1:0] far_5_5765_1;    relay_conn far_5_5765_1_a(.in(far_5_5765_0[0]), .out(far_5_5765_1[0]));    relay_conn far_5_5765_1_b(.in(far_5_5765_0[1]), .out(far_5_5765_1[1]));
    assign layer_5[665] = ~(far_5_5765_1[0] | far_5_5765_1[1]); 
    wire [1:0] far_5_5766_0;    relay_conn far_5_5766_0_a(.in(layer_4[645]), .out(far_5_5766_0[0]));    relay_conn far_5_5766_0_b(.in(layer_4[559]), .out(far_5_5766_0[1]));
    wire [1:0] far_5_5766_1;    relay_conn far_5_5766_1_a(.in(far_5_5766_0[0]), .out(far_5_5766_1[0]));    relay_conn far_5_5766_1_b(.in(far_5_5766_0[1]), .out(far_5_5766_1[1]));
    assign layer_5[666] = far_5_5766_1[1]; 
    wire [1:0] far_5_5767_0;    relay_conn far_5_5767_0_a(.in(layer_4[325]), .out(far_5_5767_0[0]));    relay_conn far_5_5767_0_b(.in(layer_4[365]), .out(far_5_5767_0[1]));
    assign layer_5[667] = ~far_5_5767_0[1]; 
    wire [1:0] far_5_5768_0;    relay_conn far_5_5768_0_a(.in(layer_4[267]), .out(far_5_5768_0[0]));    relay_conn far_5_5768_0_b(.in(layer_4[319]), .out(far_5_5768_0[1]));
    assign layer_5[668] = ~far_5_5768_0[1]; 
    wire [1:0] far_5_5769_0;    relay_conn far_5_5769_0_a(.in(layer_4[186]), .out(far_5_5769_0[0]));    relay_conn far_5_5769_0_b(.in(layer_4[94]), .out(far_5_5769_0[1]));
    wire [1:0] far_5_5769_1;    relay_conn far_5_5769_1_a(.in(far_5_5769_0[0]), .out(far_5_5769_1[0]));    relay_conn far_5_5769_1_b(.in(far_5_5769_0[1]), .out(far_5_5769_1[1]));
    assign layer_5[669] = ~far_5_5769_1[1] | (far_5_5769_1[0] & far_5_5769_1[1]); 
    wire [1:0] far_5_5770_0;    relay_conn far_5_5770_0_a(.in(layer_4[485]), .out(far_5_5770_0[0]));    relay_conn far_5_5770_0_b(.in(layer_4[398]), .out(far_5_5770_0[1]));
    wire [1:0] far_5_5770_1;    relay_conn far_5_5770_1_a(.in(far_5_5770_0[0]), .out(far_5_5770_1[0]));    relay_conn far_5_5770_1_b(.in(far_5_5770_0[1]), .out(far_5_5770_1[1]));
    assign layer_5[670] = ~far_5_5770_1[1]; 
    assign layer_5[671] = ~layer_4[330]; 
    wire [1:0] far_5_5772_0;    relay_conn far_5_5772_0_a(.in(layer_4[451]), .out(far_5_5772_0[0]));    relay_conn far_5_5772_0_b(.in(layer_4[483]), .out(far_5_5772_0[1]));
    assign layer_5[672] = ~far_5_5772_0[1]; 
    assign layer_5[673] = layer_4[845] & layer_4[823]; 
    assign layer_5[674] = layer_4[429] | layer_4[415]; 
    assign layer_5[675] = ~layer_4[1012]; 
    wire [1:0] far_5_5776_0;    relay_conn far_5_5776_0_a(.in(layer_4[387]), .out(far_5_5776_0[0]));    relay_conn far_5_5776_0_b(.in(layer_4[267]), .out(far_5_5776_0[1]));
    wire [1:0] far_5_5776_1;    relay_conn far_5_5776_1_a(.in(far_5_5776_0[0]), .out(far_5_5776_1[0]));    relay_conn far_5_5776_1_b(.in(far_5_5776_0[1]), .out(far_5_5776_1[1]));
    wire [1:0] far_5_5776_2;    relay_conn far_5_5776_2_a(.in(far_5_5776_1[0]), .out(far_5_5776_2[0]));    relay_conn far_5_5776_2_b(.in(far_5_5776_1[1]), .out(far_5_5776_2[1]));
    assign layer_5[676] = far_5_5776_2[0] ^ far_5_5776_2[1]; 
    wire [1:0] far_5_5777_0;    relay_conn far_5_5777_0_a(.in(layer_4[763]), .out(far_5_5777_0[0]));    relay_conn far_5_5777_0_b(.in(layer_4[716]), .out(far_5_5777_0[1]));
    assign layer_5[677] = far_5_5777_0[0] & ~far_5_5777_0[1]; 
    wire [1:0] far_5_5778_0;    relay_conn far_5_5778_0_a(.in(layer_4[74]), .out(far_5_5778_0[0]));    relay_conn far_5_5778_0_b(.in(layer_4[13]), .out(far_5_5778_0[1]));
    assign layer_5[678] = ~far_5_5778_0[1] | (far_5_5778_0[0] & far_5_5778_0[1]); 
    wire [1:0] far_5_5779_0;    relay_conn far_5_5779_0_a(.in(layer_4[502]), .out(far_5_5779_0[0]));    relay_conn far_5_5779_0_b(.in(layer_4[553]), .out(far_5_5779_0[1]));
    assign layer_5[679] = ~(far_5_5779_0[0] | far_5_5779_0[1]); 
    assign layer_5[680] = ~layer_4[967] | (layer_4[967] & layer_4[994]); 
    wire [1:0] far_5_5781_0;    relay_conn far_5_5781_0_a(.in(layer_4[636]), .out(far_5_5781_0[0]));    relay_conn far_5_5781_0_b(.in(layer_4[718]), .out(far_5_5781_0[1]));
    wire [1:0] far_5_5781_1;    relay_conn far_5_5781_1_a(.in(far_5_5781_0[0]), .out(far_5_5781_1[0]));    relay_conn far_5_5781_1_b(.in(far_5_5781_0[1]), .out(far_5_5781_1[1]));
    assign layer_5[681] = ~far_5_5781_1[1]; 
    assign layer_5[682] = ~layer_4[901]; 
    wire [1:0] far_5_5783_0;    relay_conn far_5_5783_0_a(.in(layer_4[40]), .out(far_5_5783_0[0]));    relay_conn far_5_5783_0_b(.in(layer_4[132]), .out(far_5_5783_0[1]));
    wire [1:0] far_5_5783_1;    relay_conn far_5_5783_1_a(.in(far_5_5783_0[0]), .out(far_5_5783_1[0]));    relay_conn far_5_5783_1_b(.in(far_5_5783_0[1]), .out(far_5_5783_1[1]));
    assign layer_5[683] = ~far_5_5783_1[0] | (far_5_5783_1[0] & far_5_5783_1[1]); 
    wire [1:0] far_5_5784_0;    relay_conn far_5_5784_0_a(.in(layer_4[502]), .out(far_5_5784_0[0]));    relay_conn far_5_5784_0_b(.in(layer_4[546]), .out(far_5_5784_0[1]));
    assign layer_5[684] = far_5_5784_0[0] | far_5_5784_0[1]; 
    wire [1:0] far_5_5785_0;    relay_conn far_5_5785_0_a(.in(layer_4[25]), .out(far_5_5785_0[0]));    relay_conn far_5_5785_0_b(.in(layer_4[129]), .out(far_5_5785_0[1]));
    wire [1:0] far_5_5785_1;    relay_conn far_5_5785_1_a(.in(far_5_5785_0[0]), .out(far_5_5785_1[0]));    relay_conn far_5_5785_1_b(.in(far_5_5785_0[1]), .out(far_5_5785_1[1]));
    wire [1:0] far_5_5785_2;    relay_conn far_5_5785_2_a(.in(far_5_5785_1[0]), .out(far_5_5785_2[0]));    relay_conn far_5_5785_2_b(.in(far_5_5785_1[1]), .out(far_5_5785_2[1]));
    assign layer_5[685] = ~far_5_5785_2[1] | (far_5_5785_2[0] & far_5_5785_2[1]); 
    assign layer_5[686] = layer_4[759]; 
    assign layer_5[687] = layer_4[836] & ~layer_4[846]; 
    wire [1:0] far_5_5788_0;    relay_conn far_5_5788_0_a(.in(layer_4[530]), .out(far_5_5788_0[0]));    relay_conn far_5_5788_0_b(.in(layer_4[419]), .out(far_5_5788_0[1]));
    wire [1:0] far_5_5788_1;    relay_conn far_5_5788_1_a(.in(far_5_5788_0[0]), .out(far_5_5788_1[0]));    relay_conn far_5_5788_1_b(.in(far_5_5788_0[1]), .out(far_5_5788_1[1]));
    wire [1:0] far_5_5788_2;    relay_conn far_5_5788_2_a(.in(far_5_5788_1[0]), .out(far_5_5788_2[0]));    relay_conn far_5_5788_2_b(.in(far_5_5788_1[1]), .out(far_5_5788_2[1]));
    assign layer_5[688] = ~far_5_5788_2[0]; 
    assign layer_5[689] = ~layer_4[322] | (layer_4[300] & layer_4[322]); 
    wire [1:0] far_5_5790_0;    relay_conn far_5_5790_0_a(.in(layer_4[267]), .out(far_5_5790_0[0]));    relay_conn far_5_5790_0_b(.in(layer_4[142]), .out(far_5_5790_0[1]));
    wire [1:0] far_5_5790_1;    relay_conn far_5_5790_1_a(.in(far_5_5790_0[0]), .out(far_5_5790_1[0]));    relay_conn far_5_5790_1_b(.in(far_5_5790_0[1]), .out(far_5_5790_1[1]));
    wire [1:0] far_5_5790_2;    relay_conn far_5_5790_2_a(.in(far_5_5790_1[0]), .out(far_5_5790_2[0]));    relay_conn far_5_5790_2_b(.in(far_5_5790_1[1]), .out(far_5_5790_2[1]));
    assign layer_5[690] = ~far_5_5790_2[0] | (far_5_5790_2[0] & far_5_5790_2[1]); 
    assign layer_5[691] = layer_4[620]; 
    assign layer_5[692] = layer_4[644] & ~layer_4[615]; 
    wire [1:0] far_5_5793_0;    relay_conn far_5_5793_0_a(.in(layer_4[665]), .out(far_5_5793_0[0]));    relay_conn far_5_5793_0_b(.in(layer_4[619]), .out(far_5_5793_0[1]));
    assign layer_5[693] = ~far_5_5793_0[1] | (far_5_5793_0[0] & far_5_5793_0[1]); 
    assign layer_5[694] = layer_4[96] & ~layer_4[94]; 
    wire [1:0] far_5_5795_0;    relay_conn far_5_5795_0_a(.in(layer_4[768]), .out(far_5_5795_0[0]));    relay_conn far_5_5795_0_b(.in(layer_4[850]), .out(far_5_5795_0[1]));
    wire [1:0] far_5_5795_1;    relay_conn far_5_5795_1_a(.in(far_5_5795_0[0]), .out(far_5_5795_1[0]));    relay_conn far_5_5795_1_b(.in(far_5_5795_0[1]), .out(far_5_5795_1[1]));
    assign layer_5[695] = far_5_5795_1[0] & ~far_5_5795_1[1]; 
    assign layer_5[696] = layer_4[437] | layer_4[436]; 
    wire [1:0] far_5_5797_0;    relay_conn far_5_5797_0_a(.in(layer_4[190]), .out(far_5_5797_0[0]));    relay_conn far_5_5797_0_b(.in(layer_4[142]), .out(far_5_5797_0[1]));
    assign layer_5[697] = far_5_5797_0[0]; 
    assign layer_5[698] = layer_4[640]; 
    wire [1:0] far_5_5799_0;    relay_conn far_5_5799_0_a(.in(layer_4[382]), .out(far_5_5799_0[0]));    relay_conn far_5_5799_0_b(.in(layer_4[435]), .out(far_5_5799_0[1]));
    assign layer_5[699] = far_5_5799_0[0]; 
    wire [1:0] far_5_5800_0;    relay_conn far_5_5800_0_a(.in(layer_4[430]), .out(far_5_5800_0[0]));    relay_conn far_5_5800_0_b(.in(layer_4[343]), .out(far_5_5800_0[1]));
    wire [1:0] far_5_5800_1;    relay_conn far_5_5800_1_a(.in(far_5_5800_0[0]), .out(far_5_5800_1[0]));    relay_conn far_5_5800_1_b(.in(far_5_5800_0[1]), .out(far_5_5800_1[1]));
    assign layer_5[700] = far_5_5800_1[1]; 
    wire [1:0] far_5_5801_0;    relay_conn far_5_5801_0_a(.in(layer_4[401]), .out(far_5_5801_0[0]));    relay_conn far_5_5801_0_b(.in(layer_4[442]), .out(far_5_5801_0[1]));
    assign layer_5[701] = ~far_5_5801_0[0] | (far_5_5801_0[0] & far_5_5801_0[1]); 
    wire [1:0] far_5_5802_0;    relay_conn far_5_5802_0_a(.in(layer_4[950]), .out(far_5_5802_0[0]));    relay_conn far_5_5802_0_b(.in(layer_4[1008]), .out(far_5_5802_0[1]));
    assign layer_5[702] = ~(far_5_5802_0[0] & far_5_5802_0[1]); 
    wire [1:0] far_5_5803_0;    relay_conn far_5_5803_0_a(.in(layer_4[911]), .out(far_5_5803_0[0]));    relay_conn far_5_5803_0_b(.in(layer_4[953]), .out(far_5_5803_0[1]));
    assign layer_5[703] = ~far_5_5803_0[0] | (far_5_5803_0[0] & far_5_5803_0[1]); 
    wire [1:0] far_5_5804_0;    relay_conn far_5_5804_0_a(.in(layer_4[215]), .out(far_5_5804_0[0]));    relay_conn far_5_5804_0_b(.in(layer_4[307]), .out(far_5_5804_0[1]));
    wire [1:0] far_5_5804_1;    relay_conn far_5_5804_1_a(.in(far_5_5804_0[0]), .out(far_5_5804_1[0]));    relay_conn far_5_5804_1_b(.in(far_5_5804_0[1]), .out(far_5_5804_1[1]));
    assign layer_5[704] = far_5_5804_1[0]; 
    wire [1:0] far_5_5805_0;    relay_conn far_5_5805_0_a(.in(layer_4[910]), .out(far_5_5805_0[0]));    relay_conn far_5_5805_0_b(.in(layer_4[830]), .out(far_5_5805_0[1]));
    wire [1:0] far_5_5805_1;    relay_conn far_5_5805_1_a(.in(far_5_5805_0[0]), .out(far_5_5805_1[0]));    relay_conn far_5_5805_1_b(.in(far_5_5805_0[1]), .out(far_5_5805_1[1]));
    assign layer_5[705] = far_5_5805_1[1]; 
    wire [1:0] far_5_5806_0;    relay_conn far_5_5806_0_a(.in(layer_4[62]), .out(far_5_5806_0[0]));    relay_conn far_5_5806_0_b(.in(layer_4[182]), .out(far_5_5806_0[1]));
    wire [1:0] far_5_5806_1;    relay_conn far_5_5806_1_a(.in(far_5_5806_0[0]), .out(far_5_5806_1[0]));    relay_conn far_5_5806_1_b(.in(far_5_5806_0[1]), .out(far_5_5806_1[1]));
    wire [1:0] far_5_5806_2;    relay_conn far_5_5806_2_a(.in(far_5_5806_1[0]), .out(far_5_5806_2[0]));    relay_conn far_5_5806_2_b(.in(far_5_5806_1[1]), .out(far_5_5806_2[1]));
    assign layer_5[706] = far_5_5806_2[1]; 
    assign layer_5[707] = ~layer_4[650] | (layer_4[679] & layer_4[650]); 
    wire [1:0] far_5_5808_0;    relay_conn far_5_5808_0_a(.in(layer_4[429]), .out(far_5_5808_0[0]));    relay_conn far_5_5808_0_b(.in(layer_4[477]), .out(far_5_5808_0[1]));
    assign layer_5[708] = far_5_5808_0[1] & ~far_5_5808_0[0]; 
    wire [1:0] far_5_5809_0;    relay_conn far_5_5809_0_a(.in(layer_4[253]), .out(far_5_5809_0[0]));    relay_conn far_5_5809_0_b(.in(layer_4[301]), .out(far_5_5809_0[1]));
    assign layer_5[709] = far_5_5809_0[0]; 
    wire [1:0] far_5_5810_0;    relay_conn far_5_5810_0_a(.in(layer_4[293]), .out(far_5_5810_0[0]));    relay_conn far_5_5810_0_b(.in(layer_4[369]), .out(far_5_5810_0[1]));
    wire [1:0] far_5_5810_1;    relay_conn far_5_5810_1_a(.in(far_5_5810_0[0]), .out(far_5_5810_1[0]));    relay_conn far_5_5810_1_b(.in(far_5_5810_0[1]), .out(far_5_5810_1[1]));
    assign layer_5[710] = ~far_5_5810_1[0] | (far_5_5810_1[0] & far_5_5810_1[1]); 
    wire [1:0] far_5_5811_0;    relay_conn far_5_5811_0_a(.in(layer_4[580]), .out(far_5_5811_0[0]));    relay_conn far_5_5811_0_b(.in(layer_4[680]), .out(far_5_5811_0[1]));
    wire [1:0] far_5_5811_1;    relay_conn far_5_5811_1_a(.in(far_5_5811_0[0]), .out(far_5_5811_1[0]));    relay_conn far_5_5811_1_b(.in(far_5_5811_0[1]), .out(far_5_5811_1[1]));
    wire [1:0] far_5_5811_2;    relay_conn far_5_5811_2_a(.in(far_5_5811_1[0]), .out(far_5_5811_2[0]));    relay_conn far_5_5811_2_b(.in(far_5_5811_1[1]), .out(far_5_5811_2[1]));
    assign layer_5[711] = far_5_5811_2[1] & ~far_5_5811_2[0]; 
    wire [1:0] far_5_5812_0;    relay_conn far_5_5812_0_a(.in(layer_4[274]), .out(far_5_5812_0[0]));    relay_conn far_5_5812_0_b(.in(layer_4[325]), .out(far_5_5812_0[1]));
    assign layer_5[712] = ~far_5_5812_0[0]; 
    assign layer_5[713] = layer_4[16] | layer_4[13]; 
    wire [1:0] far_5_5814_0;    relay_conn far_5_5814_0_a(.in(layer_4[690]), .out(far_5_5814_0[0]));    relay_conn far_5_5814_0_b(.in(layer_4[743]), .out(far_5_5814_0[1]));
    assign layer_5[714] = ~(far_5_5814_0[0] & far_5_5814_0[1]); 
    wire [1:0] far_5_5815_0;    relay_conn far_5_5815_0_a(.in(layer_4[52]), .out(far_5_5815_0[0]));    relay_conn far_5_5815_0_b(.in(layer_4[6]), .out(far_5_5815_0[1]));
    assign layer_5[715] = ~far_5_5815_0[1]; 
    wire [1:0] far_5_5816_0;    relay_conn far_5_5816_0_a(.in(layer_4[656]), .out(far_5_5816_0[0]));    relay_conn far_5_5816_0_b(.in(layer_4[594]), .out(far_5_5816_0[1]));
    assign layer_5[716] = far_5_5816_0[1] & ~far_5_5816_0[0]; 
    wire [1:0] far_5_5817_0;    relay_conn far_5_5817_0_a(.in(layer_4[438]), .out(far_5_5817_0[0]));    relay_conn far_5_5817_0_b(.in(layer_4[370]), .out(far_5_5817_0[1]));
    wire [1:0] far_5_5817_1;    relay_conn far_5_5817_1_a(.in(far_5_5817_0[0]), .out(far_5_5817_1[0]));    relay_conn far_5_5817_1_b(.in(far_5_5817_0[1]), .out(far_5_5817_1[1]));
    assign layer_5[717] = far_5_5817_1[0]; 
    wire [1:0] far_5_5818_0;    relay_conn far_5_5818_0_a(.in(layer_4[650]), .out(far_5_5818_0[0]));    relay_conn far_5_5818_0_b(.in(layer_4[583]), .out(far_5_5818_0[1]));
    wire [1:0] far_5_5818_1;    relay_conn far_5_5818_1_a(.in(far_5_5818_0[0]), .out(far_5_5818_1[0]));    relay_conn far_5_5818_1_b(.in(far_5_5818_0[1]), .out(far_5_5818_1[1]));
    assign layer_5[718] = far_5_5818_1[0] | far_5_5818_1[1]; 
    wire [1:0] far_5_5819_0;    relay_conn far_5_5819_0_a(.in(layer_4[200]), .out(far_5_5819_0[0]));    relay_conn far_5_5819_0_b(.in(layer_4[78]), .out(far_5_5819_0[1]));
    wire [1:0] far_5_5819_1;    relay_conn far_5_5819_1_a(.in(far_5_5819_0[0]), .out(far_5_5819_1[0]));    relay_conn far_5_5819_1_b(.in(far_5_5819_0[1]), .out(far_5_5819_1[1]));
    wire [1:0] far_5_5819_2;    relay_conn far_5_5819_2_a(.in(far_5_5819_1[0]), .out(far_5_5819_2[0]));    relay_conn far_5_5819_2_b(.in(far_5_5819_1[1]), .out(far_5_5819_2[1]));
    assign layer_5[719] = ~far_5_5819_2[1]; 
    assign layer_5[720] = ~layer_4[133] | (layer_4[145] & layer_4[133]); 
    assign layer_5[721] = layer_4[997] & ~layer_4[984]; 
    assign layer_5[722] = layer_4[598] & ~layer_4[576]; 
    wire [1:0] far_5_5823_0;    relay_conn far_5_5823_0_a(.in(layer_4[164]), .out(far_5_5823_0[0]));    relay_conn far_5_5823_0_b(.in(layer_4[266]), .out(far_5_5823_0[1]));
    wire [1:0] far_5_5823_1;    relay_conn far_5_5823_1_a(.in(far_5_5823_0[0]), .out(far_5_5823_1[0]));    relay_conn far_5_5823_1_b(.in(far_5_5823_0[1]), .out(far_5_5823_1[1]));
    wire [1:0] far_5_5823_2;    relay_conn far_5_5823_2_a(.in(far_5_5823_1[0]), .out(far_5_5823_2[0]));    relay_conn far_5_5823_2_b(.in(far_5_5823_1[1]), .out(far_5_5823_2[1]));
    assign layer_5[723] = ~far_5_5823_2[1]; 
    assign layer_5[724] = ~(layer_4[66] | layer_4[88]); 
    wire [1:0] far_5_5825_0;    relay_conn far_5_5825_0_a(.in(layer_4[454]), .out(far_5_5825_0[0]));    relay_conn far_5_5825_0_b(.in(layer_4[400]), .out(far_5_5825_0[1]));
    assign layer_5[725] = far_5_5825_0[0] | far_5_5825_0[1]; 
    wire [1:0] far_5_5826_0;    relay_conn far_5_5826_0_a(.in(layer_4[650]), .out(far_5_5826_0[0]));    relay_conn far_5_5826_0_b(.in(layer_4[718]), .out(far_5_5826_0[1]));
    wire [1:0] far_5_5826_1;    relay_conn far_5_5826_1_a(.in(far_5_5826_0[0]), .out(far_5_5826_1[0]));    relay_conn far_5_5826_1_b(.in(far_5_5826_0[1]), .out(far_5_5826_1[1]));
    assign layer_5[726] = ~(far_5_5826_1[0] & far_5_5826_1[1]); 
    wire [1:0] far_5_5827_0;    relay_conn far_5_5827_0_a(.in(layer_4[958]), .out(far_5_5827_0[0]));    relay_conn far_5_5827_0_b(.in(layer_4[875]), .out(far_5_5827_0[1]));
    wire [1:0] far_5_5827_1;    relay_conn far_5_5827_1_a(.in(far_5_5827_0[0]), .out(far_5_5827_1[0]));    relay_conn far_5_5827_1_b(.in(far_5_5827_0[1]), .out(far_5_5827_1[1]));
    assign layer_5[727] = far_5_5827_1[1]; 
    wire [1:0] far_5_5828_0;    relay_conn far_5_5828_0_a(.in(layer_4[235]), .out(far_5_5828_0[0]));    relay_conn far_5_5828_0_b(.in(layer_4[354]), .out(far_5_5828_0[1]));
    wire [1:0] far_5_5828_1;    relay_conn far_5_5828_1_a(.in(far_5_5828_0[0]), .out(far_5_5828_1[0]));    relay_conn far_5_5828_1_b(.in(far_5_5828_0[1]), .out(far_5_5828_1[1]));
    wire [1:0] far_5_5828_2;    relay_conn far_5_5828_2_a(.in(far_5_5828_1[0]), .out(far_5_5828_2[0]));    relay_conn far_5_5828_2_b(.in(far_5_5828_1[1]), .out(far_5_5828_2[1]));
    assign layer_5[728] = ~(far_5_5828_2[0] & far_5_5828_2[1]); 
    wire [1:0] far_5_5829_0;    relay_conn far_5_5829_0_a(.in(layer_4[468]), .out(far_5_5829_0[0]));    relay_conn far_5_5829_0_b(.in(layer_4[543]), .out(far_5_5829_0[1]));
    wire [1:0] far_5_5829_1;    relay_conn far_5_5829_1_a(.in(far_5_5829_0[0]), .out(far_5_5829_1[0]));    relay_conn far_5_5829_1_b(.in(far_5_5829_0[1]), .out(far_5_5829_1[1]));
    assign layer_5[729] = far_5_5829_1[0] | far_5_5829_1[1]; 
    wire [1:0] far_5_5830_0;    relay_conn far_5_5830_0_a(.in(layer_4[765]), .out(far_5_5830_0[0]));    relay_conn far_5_5830_0_b(.in(layer_4[653]), .out(far_5_5830_0[1]));
    wire [1:0] far_5_5830_1;    relay_conn far_5_5830_1_a(.in(far_5_5830_0[0]), .out(far_5_5830_1[0]));    relay_conn far_5_5830_1_b(.in(far_5_5830_0[1]), .out(far_5_5830_1[1]));
    wire [1:0] far_5_5830_2;    relay_conn far_5_5830_2_a(.in(far_5_5830_1[0]), .out(far_5_5830_2[0]));    relay_conn far_5_5830_2_b(.in(far_5_5830_1[1]), .out(far_5_5830_2[1]));
    assign layer_5[730] = far_5_5830_2[0] & far_5_5830_2[1]; 
    wire [1:0] far_5_5831_0;    relay_conn far_5_5831_0_a(.in(layer_4[644]), .out(far_5_5831_0[0]));    relay_conn far_5_5831_0_b(.in(layer_4[736]), .out(far_5_5831_0[1]));
    wire [1:0] far_5_5831_1;    relay_conn far_5_5831_1_a(.in(far_5_5831_0[0]), .out(far_5_5831_1[0]));    relay_conn far_5_5831_1_b(.in(far_5_5831_0[1]), .out(far_5_5831_1[1]));
    assign layer_5[731] = far_5_5831_1[0] & ~far_5_5831_1[1]; 
    wire [1:0] far_5_5832_0;    relay_conn far_5_5832_0_a(.in(layer_4[783]), .out(far_5_5832_0[0]));    relay_conn far_5_5832_0_b(.in(layer_4[850]), .out(far_5_5832_0[1]));
    wire [1:0] far_5_5832_1;    relay_conn far_5_5832_1_a(.in(far_5_5832_0[0]), .out(far_5_5832_1[0]));    relay_conn far_5_5832_1_b(.in(far_5_5832_0[1]), .out(far_5_5832_1[1]));
    assign layer_5[732] = ~far_5_5832_1[0]; 
    wire [1:0] far_5_5833_0;    relay_conn far_5_5833_0_a(.in(layer_4[26]), .out(far_5_5833_0[0]));    relay_conn far_5_5833_0_b(.in(layer_4[97]), .out(far_5_5833_0[1]));
    wire [1:0] far_5_5833_1;    relay_conn far_5_5833_1_a(.in(far_5_5833_0[0]), .out(far_5_5833_1[0]));    relay_conn far_5_5833_1_b(.in(far_5_5833_0[1]), .out(far_5_5833_1[1]));
    assign layer_5[733] = far_5_5833_1[0] | far_5_5833_1[1]; 
    assign layer_5[734] = layer_4[103] | layer_4[129]; 
    wire [1:0] far_5_5835_0;    relay_conn far_5_5835_0_a(.in(layer_4[310]), .out(far_5_5835_0[0]));    relay_conn far_5_5835_0_b(.in(layer_4[202]), .out(far_5_5835_0[1]));
    wire [1:0] far_5_5835_1;    relay_conn far_5_5835_1_a(.in(far_5_5835_0[0]), .out(far_5_5835_1[0]));    relay_conn far_5_5835_1_b(.in(far_5_5835_0[1]), .out(far_5_5835_1[1]));
    wire [1:0] far_5_5835_2;    relay_conn far_5_5835_2_a(.in(far_5_5835_1[0]), .out(far_5_5835_2[0]));    relay_conn far_5_5835_2_b(.in(far_5_5835_1[1]), .out(far_5_5835_2[1]));
    assign layer_5[735] = far_5_5835_2[0] | far_5_5835_2[1]; 
    wire [1:0] far_5_5836_0;    relay_conn far_5_5836_0_a(.in(layer_4[381]), .out(far_5_5836_0[0]));    relay_conn far_5_5836_0_b(.in(layer_4[294]), .out(far_5_5836_0[1]));
    wire [1:0] far_5_5836_1;    relay_conn far_5_5836_1_a(.in(far_5_5836_0[0]), .out(far_5_5836_1[0]));    relay_conn far_5_5836_1_b(.in(far_5_5836_0[1]), .out(far_5_5836_1[1]));
    assign layer_5[736] = ~far_5_5836_1[1]; 
    assign layer_5[737] = ~(layer_4[692] | layer_4[684]); 
    assign layer_5[738] = ~(layer_4[360] & layer_4[337]); 
    assign layer_5[739] = ~layer_4[654]; 
    wire [1:0] far_5_5840_0;    relay_conn far_5_5840_0_a(.in(layer_4[341]), .out(far_5_5840_0[0]));    relay_conn far_5_5840_0_b(.in(layer_4[266]), .out(far_5_5840_0[1]));
    wire [1:0] far_5_5840_1;    relay_conn far_5_5840_1_a(.in(far_5_5840_0[0]), .out(far_5_5840_1[0]));    relay_conn far_5_5840_1_b(.in(far_5_5840_0[1]), .out(far_5_5840_1[1]));
    assign layer_5[740] = far_5_5840_1[0] & far_5_5840_1[1]; 
    wire [1:0] far_5_5841_0;    relay_conn far_5_5841_0_a(.in(layer_4[789]), .out(far_5_5841_0[0]));    relay_conn far_5_5841_0_b(.in(layer_4[665]), .out(far_5_5841_0[1]));
    wire [1:0] far_5_5841_1;    relay_conn far_5_5841_1_a(.in(far_5_5841_0[0]), .out(far_5_5841_1[0]));    relay_conn far_5_5841_1_b(.in(far_5_5841_0[1]), .out(far_5_5841_1[1]));
    wire [1:0] far_5_5841_2;    relay_conn far_5_5841_2_a(.in(far_5_5841_1[0]), .out(far_5_5841_2[0]));    relay_conn far_5_5841_2_b(.in(far_5_5841_1[1]), .out(far_5_5841_2[1]));
    assign layer_5[741] = ~(far_5_5841_2[0] ^ far_5_5841_2[1]); 
    wire [1:0] far_5_5842_0;    relay_conn far_5_5842_0_a(.in(layer_4[286]), .out(far_5_5842_0[0]));    relay_conn far_5_5842_0_b(.in(layer_4[409]), .out(far_5_5842_0[1]));
    wire [1:0] far_5_5842_1;    relay_conn far_5_5842_1_a(.in(far_5_5842_0[0]), .out(far_5_5842_1[0]));    relay_conn far_5_5842_1_b(.in(far_5_5842_0[1]), .out(far_5_5842_1[1]));
    wire [1:0] far_5_5842_2;    relay_conn far_5_5842_2_a(.in(far_5_5842_1[0]), .out(far_5_5842_2[0]));    relay_conn far_5_5842_2_b(.in(far_5_5842_1[1]), .out(far_5_5842_2[1]));
    assign layer_5[742] = ~far_5_5842_2[0]; 
    wire [1:0] far_5_5843_0;    relay_conn far_5_5843_0_a(.in(layer_4[339]), .out(far_5_5843_0[0]));    relay_conn far_5_5843_0_b(.in(layer_4[301]), .out(far_5_5843_0[1]));
    assign layer_5[743] = ~(far_5_5843_0[0] | far_5_5843_0[1]); 
    assign layer_5[744] = ~layer_4[936] | (layer_4[936] & layer_4[922]); 
    assign layer_5[745] = ~(layer_4[746] & layer_4[718]); 
    wire [1:0] far_5_5846_0;    relay_conn far_5_5846_0_a(.in(layer_4[300]), .out(far_5_5846_0[0]));    relay_conn far_5_5846_0_b(.in(layer_4[403]), .out(far_5_5846_0[1]));
    wire [1:0] far_5_5846_1;    relay_conn far_5_5846_1_a(.in(far_5_5846_0[0]), .out(far_5_5846_1[0]));    relay_conn far_5_5846_1_b(.in(far_5_5846_0[1]), .out(far_5_5846_1[1]));
    wire [1:0] far_5_5846_2;    relay_conn far_5_5846_2_a(.in(far_5_5846_1[0]), .out(far_5_5846_2[0]));    relay_conn far_5_5846_2_b(.in(far_5_5846_1[1]), .out(far_5_5846_2[1]));
    assign layer_5[746] = ~far_5_5846_2[1]; 
    wire [1:0] far_5_5847_0;    relay_conn far_5_5847_0_a(.in(layer_4[127]), .out(far_5_5847_0[0]));    relay_conn far_5_5847_0_b(.in(layer_4[89]), .out(far_5_5847_0[1]));
    assign layer_5[747] = ~far_5_5847_0[0] | (far_5_5847_0[0] & far_5_5847_0[1]); 
    wire [1:0] far_5_5848_0;    relay_conn far_5_5848_0_a(.in(layer_4[755]), .out(far_5_5848_0[0]));    relay_conn far_5_5848_0_b(.in(layer_4[650]), .out(far_5_5848_0[1]));
    wire [1:0] far_5_5848_1;    relay_conn far_5_5848_1_a(.in(far_5_5848_0[0]), .out(far_5_5848_1[0]));    relay_conn far_5_5848_1_b(.in(far_5_5848_0[1]), .out(far_5_5848_1[1]));
    wire [1:0] far_5_5848_2;    relay_conn far_5_5848_2_a(.in(far_5_5848_1[0]), .out(far_5_5848_2[0]));    relay_conn far_5_5848_2_b(.in(far_5_5848_1[1]), .out(far_5_5848_2[1]));
    assign layer_5[748] = ~far_5_5848_2[1]; 
    wire [1:0] far_5_5849_0;    relay_conn far_5_5849_0_a(.in(layer_4[22]), .out(far_5_5849_0[0]));    relay_conn far_5_5849_0_b(.in(layer_4[141]), .out(far_5_5849_0[1]));
    wire [1:0] far_5_5849_1;    relay_conn far_5_5849_1_a(.in(far_5_5849_0[0]), .out(far_5_5849_1[0]));    relay_conn far_5_5849_1_b(.in(far_5_5849_0[1]), .out(far_5_5849_1[1]));
    wire [1:0] far_5_5849_2;    relay_conn far_5_5849_2_a(.in(far_5_5849_1[0]), .out(far_5_5849_2[0]));    relay_conn far_5_5849_2_b(.in(far_5_5849_1[1]), .out(far_5_5849_2[1]));
    assign layer_5[749] = ~far_5_5849_2[1] | (far_5_5849_2[0] & far_5_5849_2[1]); 
    wire [1:0] far_5_5850_0;    relay_conn far_5_5850_0_a(.in(layer_4[472]), .out(far_5_5850_0[0]));    relay_conn far_5_5850_0_b(.in(layer_4[523]), .out(far_5_5850_0[1]));
    assign layer_5[750] = ~far_5_5850_0[0]; 
    wire [1:0] far_5_5851_0;    relay_conn far_5_5851_0_a(.in(layer_4[536]), .out(far_5_5851_0[0]));    relay_conn far_5_5851_0_b(.in(layer_4[419]), .out(far_5_5851_0[1]));
    wire [1:0] far_5_5851_1;    relay_conn far_5_5851_1_a(.in(far_5_5851_0[0]), .out(far_5_5851_1[0]));    relay_conn far_5_5851_1_b(.in(far_5_5851_0[1]), .out(far_5_5851_1[1]));
    wire [1:0] far_5_5851_2;    relay_conn far_5_5851_2_a(.in(far_5_5851_1[0]), .out(far_5_5851_2[0]));    relay_conn far_5_5851_2_b(.in(far_5_5851_1[1]), .out(far_5_5851_2[1]));
    assign layer_5[751] = far_5_5851_2[1] & ~far_5_5851_2[0]; 
    wire [1:0] far_5_5852_0;    relay_conn far_5_5852_0_a(.in(layer_4[656]), .out(far_5_5852_0[0]));    relay_conn far_5_5852_0_b(.in(layer_4[780]), .out(far_5_5852_0[1]));
    wire [1:0] far_5_5852_1;    relay_conn far_5_5852_1_a(.in(far_5_5852_0[0]), .out(far_5_5852_1[0]));    relay_conn far_5_5852_1_b(.in(far_5_5852_0[1]), .out(far_5_5852_1[1]));
    wire [1:0] far_5_5852_2;    relay_conn far_5_5852_2_a(.in(far_5_5852_1[0]), .out(far_5_5852_2[0]));    relay_conn far_5_5852_2_b(.in(far_5_5852_1[1]), .out(far_5_5852_2[1]));
    assign layer_5[752] = ~(far_5_5852_2[0] & far_5_5852_2[1]); 
    wire [1:0] far_5_5853_0;    relay_conn far_5_5853_0_a(.in(layer_4[186]), .out(far_5_5853_0[0]));    relay_conn far_5_5853_0_b(.in(layer_4[123]), .out(far_5_5853_0[1]));
    assign layer_5[753] = ~far_5_5853_0[1]; 
    wire [1:0] far_5_5854_0;    relay_conn far_5_5854_0_a(.in(layer_4[264]), .out(far_5_5854_0[0]));    relay_conn far_5_5854_0_b(.in(layer_4[301]), .out(far_5_5854_0[1]));
    assign layer_5[754] = ~far_5_5854_0[0]; 
    wire [1:0] far_5_5855_0;    relay_conn far_5_5855_0_a(.in(layer_4[207]), .out(far_5_5855_0[0]));    relay_conn far_5_5855_0_b(.in(layer_4[171]), .out(far_5_5855_0[1]));
    assign layer_5[755] = far_5_5855_0[1]; 
    wire [1:0] far_5_5856_0;    relay_conn far_5_5856_0_a(.in(layer_4[768]), .out(far_5_5856_0[0]));    relay_conn far_5_5856_0_b(.in(layer_4[657]), .out(far_5_5856_0[1]));
    wire [1:0] far_5_5856_1;    relay_conn far_5_5856_1_a(.in(far_5_5856_0[0]), .out(far_5_5856_1[0]));    relay_conn far_5_5856_1_b(.in(far_5_5856_0[1]), .out(far_5_5856_1[1]));
    wire [1:0] far_5_5856_2;    relay_conn far_5_5856_2_a(.in(far_5_5856_1[0]), .out(far_5_5856_2[0]));    relay_conn far_5_5856_2_b(.in(far_5_5856_1[1]), .out(far_5_5856_2[1]));
    assign layer_5[756] = far_5_5856_2[0] | far_5_5856_2[1]; 
    wire [1:0] far_5_5857_0;    relay_conn far_5_5857_0_a(.in(layer_4[589]), .out(far_5_5857_0[0]));    relay_conn far_5_5857_0_b(.in(layer_4[622]), .out(far_5_5857_0[1]));
    assign layer_5[757] = far_5_5857_0[0] & far_5_5857_0[1]; 
    assign layer_5[758] = layer_4[127]; 
    wire [1:0] far_5_5859_0;    relay_conn far_5_5859_0_a(.in(layer_4[699]), .out(far_5_5859_0[0]));    relay_conn far_5_5859_0_b(.in(layer_4[652]), .out(far_5_5859_0[1]));
    assign layer_5[759] = far_5_5859_0[0] & far_5_5859_0[1]; 
    assign layer_5[760] = ~layer_4[425]; 
    wire [1:0] far_5_5861_0;    relay_conn far_5_5861_0_a(.in(layer_4[731]), .out(far_5_5861_0[0]));    relay_conn far_5_5861_0_b(.in(layer_4[643]), .out(far_5_5861_0[1]));
    wire [1:0] far_5_5861_1;    relay_conn far_5_5861_1_a(.in(far_5_5861_0[0]), .out(far_5_5861_1[0]));    relay_conn far_5_5861_1_b(.in(far_5_5861_0[1]), .out(far_5_5861_1[1]));
    assign layer_5[761] = far_5_5861_1[1]; 
    wire [1:0] far_5_5862_0;    relay_conn far_5_5862_0_a(.in(layer_4[298]), .out(far_5_5862_0[0]));    relay_conn far_5_5862_0_b(.in(layer_4[186]), .out(far_5_5862_0[1]));
    wire [1:0] far_5_5862_1;    relay_conn far_5_5862_1_a(.in(far_5_5862_0[0]), .out(far_5_5862_1[0]));    relay_conn far_5_5862_1_b(.in(far_5_5862_0[1]), .out(far_5_5862_1[1]));
    wire [1:0] far_5_5862_2;    relay_conn far_5_5862_2_a(.in(far_5_5862_1[0]), .out(far_5_5862_2[0]));    relay_conn far_5_5862_2_b(.in(far_5_5862_1[1]), .out(far_5_5862_2[1]));
    assign layer_5[762] = ~(far_5_5862_2[0] & far_5_5862_2[1]); 
    wire [1:0] far_5_5863_0;    relay_conn far_5_5863_0_a(.in(layer_4[674]), .out(far_5_5863_0[0]));    relay_conn far_5_5863_0_b(.in(layer_4[764]), .out(far_5_5863_0[1]));
    wire [1:0] far_5_5863_1;    relay_conn far_5_5863_1_a(.in(far_5_5863_0[0]), .out(far_5_5863_1[0]));    relay_conn far_5_5863_1_b(.in(far_5_5863_0[1]), .out(far_5_5863_1[1]));
    assign layer_5[763] = ~far_5_5863_1[1]; 
    wire [1:0] far_5_5864_0;    relay_conn far_5_5864_0_a(.in(layer_4[185]), .out(far_5_5864_0[0]));    relay_conn far_5_5864_0_b(.in(layer_4[84]), .out(far_5_5864_0[1]));
    wire [1:0] far_5_5864_1;    relay_conn far_5_5864_1_a(.in(far_5_5864_0[0]), .out(far_5_5864_1[0]));    relay_conn far_5_5864_1_b(.in(far_5_5864_0[1]), .out(far_5_5864_1[1]));
    wire [1:0] far_5_5864_2;    relay_conn far_5_5864_2_a(.in(far_5_5864_1[0]), .out(far_5_5864_2[0]));    relay_conn far_5_5864_2_b(.in(far_5_5864_1[1]), .out(far_5_5864_2[1]));
    assign layer_5[764] = ~far_5_5864_2[1]; 
    wire [1:0] far_5_5865_0;    relay_conn far_5_5865_0_a(.in(layer_4[1014]), .out(far_5_5865_0[0]));    relay_conn far_5_5865_0_b(.in(layer_4[905]), .out(far_5_5865_0[1]));
    wire [1:0] far_5_5865_1;    relay_conn far_5_5865_1_a(.in(far_5_5865_0[0]), .out(far_5_5865_1[0]));    relay_conn far_5_5865_1_b(.in(far_5_5865_0[1]), .out(far_5_5865_1[1]));
    wire [1:0] far_5_5865_2;    relay_conn far_5_5865_2_a(.in(far_5_5865_1[0]), .out(far_5_5865_2[0]));    relay_conn far_5_5865_2_b(.in(far_5_5865_1[1]), .out(far_5_5865_2[1]));
    assign layer_5[765] = far_5_5865_2[0] & far_5_5865_2[1]; 
    wire [1:0] far_5_5866_0;    relay_conn far_5_5866_0_a(.in(layer_4[291]), .out(far_5_5866_0[0]));    relay_conn far_5_5866_0_b(.in(layer_4[368]), .out(far_5_5866_0[1]));
    wire [1:0] far_5_5866_1;    relay_conn far_5_5866_1_a(.in(far_5_5866_0[0]), .out(far_5_5866_1[0]));    relay_conn far_5_5866_1_b(.in(far_5_5866_0[1]), .out(far_5_5866_1[1]));
    assign layer_5[766] = far_5_5866_1[0]; 
    assign layer_5[767] = ~(layer_4[167] & layer_4[158]); 
    wire [1:0] far_5_5868_0;    relay_conn far_5_5868_0_a(.in(layer_4[316]), .out(far_5_5868_0[0]));    relay_conn far_5_5868_0_b(.in(layer_4[402]), .out(far_5_5868_0[1]));
    wire [1:0] far_5_5868_1;    relay_conn far_5_5868_1_a(.in(far_5_5868_0[0]), .out(far_5_5868_1[0]));    relay_conn far_5_5868_1_b(.in(far_5_5868_0[1]), .out(far_5_5868_1[1]));
    assign layer_5[768] = ~far_5_5868_1[0]; 
    wire [1:0] far_5_5869_0;    relay_conn far_5_5869_0_a(.in(layer_4[964]), .out(far_5_5869_0[0]));    relay_conn far_5_5869_0_b(.in(layer_4[850]), .out(far_5_5869_0[1]));
    wire [1:0] far_5_5869_1;    relay_conn far_5_5869_1_a(.in(far_5_5869_0[0]), .out(far_5_5869_1[0]));    relay_conn far_5_5869_1_b(.in(far_5_5869_0[1]), .out(far_5_5869_1[1]));
    wire [1:0] far_5_5869_2;    relay_conn far_5_5869_2_a(.in(far_5_5869_1[0]), .out(far_5_5869_2[0]));    relay_conn far_5_5869_2_b(.in(far_5_5869_1[1]), .out(far_5_5869_2[1]));
    assign layer_5[769] = far_5_5869_2[1]; 
    assign layer_5[770] = layer_4[608]; 
    wire [1:0] far_5_5871_0;    relay_conn far_5_5871_0_a(.in(layer_4[832]), .out(far_5_5871_0[0]));    relay_conn far_5_5871_0_b(.in(layer_4[886]), .out(far_5_5871_0[1]));
    assign layer_5[771] = ~far_5_5871_0[0] | (far_5_5871_0[0] & far_5_5871_0[1]); 
    wire [1:0] far_5_5872_0;    relay_conn far_5_5872_0_a(.in(layer_4[291]), .out(far_5_5872_0[0]));    relay_conn far_5_5872_0_b(.in(layer_4[215]), .out(far_5_5872_0[1]));
    wire [1:0] far_5_5872_1;    relay_conn far_5_5872_1_a(.in(far_5_5872_0[0]), .out(far_5_5872_1[0]));    relay_conn far_5_5872_1_b(.in(far_5_5872_0[1]), .out(far_5_5872_1[1]));
    assign layer_5[772] = far_5_5872_1[1]; 
    wire [1:0] far_5_5873_0;    relay_conn far_5_5873_0_a(.in(layer_4[106]), .out(far_5_5873_0[0]));    relay_conn far_5_5873_0_b(.in(layer_4[64]), .out(far_5_5873_0[1]));
    assign layer_5[773] = far_5_5873_0[1] & ~far_5_5873_0[0]; 
    wire [1:0] far_5_5874_0;    relay_conn far_5_5874_0_a(.in(layer_4[428]), .out(far_5_5874_0[0]));    relay_conn far_5_5874_0_b(.in(layer_4[369]), .out(far_5_5874_0[1]));
    assign layer_5[774] = ~far_5_5874_0[0]; 
    wire [1:0] far_5_5875_0;    relay_conn far_5_5875_0_a(.in(layer_4[875]), .out(far_5_5875_0[0]));    relay_conn far_5_5875_0_b(.in(layer_4[958]), .out(far_5_5875_0[1]));
    wire [1:0] far_5_5875_1;    relay_conn far_5_5875_1_a(.in(far_5_5875_0[0]), .out(far_5_5875_1[0]));    relay_conn far_5_5875_1_b(.in(far_5_5875_0[1]), .out(far_5_5875_1[1]));
    assign layer_5[775] = far_5_5875_1[0]; 
    assign layer_5[776] = ~layer_4[604]; 
    assign layer_5[777] = ~(layer_4[299] | layer_4[282]); 
    wire [1:0] far_5_5878_0;    relay_conn far_5_5878_0_a(.in(layer_4[747]), .out(far_5_5878_0[0]));    relay_conn far_5_5878_0_b(.in(layer_4[871]), .out(far_5_5878_0[1]));
    wire [1:0] far_5_5878_1;    relay_conn far_5_5878_1_a(.in(far_5_5878_0[0]), .out(far_5_5878_1[0]));    relay_conn far_5_5878_1_b(.in(far_5_5878_0[1]), .out(far_5_5878_1[1]));
    wire [1:0] far_5_5878_2;    relay_conn far_5_5878_2_a(.in(far_5_5878_1[0]), .out(far_5_5878_2[0]));    relay_conn far_5_5878_2_b(.in(far_5_5878_1[1]), .out(far_5_5878_2[1]));
    assign layer_5[778] = far_5_5878_2[0]; 
    assign layer_5[779] = layer_4[850]; 
    wire [1:0] far_5_5880_0;    relay_conn far_5_5880_0_a(.in(layer_4[767]), .out(far_5_5880_0[0]));    relay_conn far_5_5880_0_b(.in(layer_4[878]), .out(far_5_5880_0[1]));
    wire [1:0] far_5_5880_1;    relay_conn far_5_5880_1_a(.in(far_5_5880_0[0]), .out(far_5_5880_1[0]));    relay_conn far_5_5880_1_b(.in(far_5_5880_0[1]), .out(far_5_5880_1[1]));
    wire [1:0] far_5_5880_2;    relay_conn far_5_5880_2_a(.in(far_5_5880_1[0]), .out(far_5_5880_2[0]));    relay_conn far_5_5880_2_b(.in(far_5_5880_1[1]), .out(far_5_5880_2[1]));
    assign layer_5[780] = far_5_5880_2[0] | far_5_5880_2[1]; 
    assign layer_5[781] = ~(layer_4[875] & layer_4[881]); 
    wire [1:0] far_5_5882_0;    relay_conn far_5_5882_0_a(.in(layer_4[854]), .out(far_5_5882_0[0]));    relay_conn far_5_5882_0_b(.in(layer_4[898]), .out(far_5_5882_0[1]));
    assign layer_5[782] = ~(far_5_5882_0[0] & far_5_5882_0[1]); 
    assign layer_5[783] = layer_4[419] & ~layer_4[437]; 
    assign layer_5[784] = ~layer_4[938] | (layer_4[921] & layer_4[938]); 
    wire [1:0] far_5_5885_0;    relay_conn far_5_5885_0_a(.in(layer_4[576]), .out(far_5_5885_0[0]));    relay_conn far_5_5885_0_b(.in(layer_4[478]), .out(far_5_5885_0[1]));
    wire [1:0] far_5_5885_1;    relay_conn far_5_5885_1_a(.in(far_5_5885_0[0]), .out(far_5_5885_1[0]));    relay_conn far_5_5885_1_b(.in(far_5_5885_0[1]), .out(far_5_5885_1[1]));
    wire [1:0] far_5_5885_2;    relay_conn far_5_5885_2_a(.in(far_5_5885_1[0]), .out(far_5_5885_2[0]));    relay_conn far_5_5885_2_b(.in(far_5_5885_1[1]), .out(far_5_5885_2[1]));
    assign layer_5[785] = far_5_5885_2[0] & far_5_5885_2[1]; 
    wire [1:0] far_5_5886_0;    relay_conn far_5_5886_0_a(.in(layer_4[830]), .out(far_5_5886_0[0]));    relay_conn far_5_5886_0_b(.in(layer_4[884]), .out(far_5_5886_0[1]));
    assign layer_5[786] = far_5_5886_0[1]; 
    wire [1:0] far_5_5887_0;    relay_conn far_5_5887_0_a(.in(layer_4[682]), .out(far_5_5887_0[0]));    relay_conn far_5_5887_0_b(.in(layer_4[639]), .out(far_5_5887_0[1]));
    assign layer_5[787] = far_5_5887_0[0]; 
    wire [1:0] far_5_5888_0;    relay_conn far_5_5888_0_a(.in(layer_4[788]), .out(far_5_5888_0[0]));    relay_conn far_5_5888_0_b(.in(layer_4[914]), .out(far_5_5888_0[1]));
    wire [1:0] far_5_5888_1;    relay_conn far_5_5888_1_a(.in(far_5_5888_0[0]), .out(far_5_5888_1[0]));    relay_conn far_5_5888_1_b(.in(far_5_5888_0[1]), .out(far_5_5888_1[1]));
    wire [1:0] far_5_5888_2;    relay_conn far_5_5888_2_a(.in(far_5_5888_1[0]), .out(far_5_5888_2[0]));    relay_conn far_5_5888_2_b(.in(far_5_5888_1[1]), .out(far_5_5888_2[1]));
    assign layer_5[788] = ~far_5_5888_2[0] | (far_5_5888_2[0] & far_5_5888_2[1]); 
    wire [1:0] far_5_5889_0;    relay_conn far_5_5889_0_a(.in(layer_4[840]), .out(far_5_5889_0[0]));    relay_conn far_5_5889_0_b(.in(layer_4[717]), .out(far_5_5889_0[1]));
    wire [1:0] far_5_5889_1;    relay_conn far_5_5889_1_a(.in(far_5_5889_0[0]), .out(far_5_5889_1[0]));    relay_conn far_5_5889_1_b(.in(far_5_5889_0[1]), .out(far_5_5889_1[1]));
    wire [1:0] far_5_5889_2;    relay_conn far_5_5889_2_a(.in(far_5_5889_1[0]), .out(far_5_5889_2[0]));    relay_conn far_5_5889_2_b(.in(far_5_5889_1[1]), .out(far_5_5889_2[1]));
    assign layer_5[789] = far_5_5889_2[0] | far_5_5889_2[1]; 
    wire [1:0] far_5_5890_0;    relay_conn far_5_5890_0_a(.in(layer_4[15]), .out(far_5_5890_0[0]));    relay_conn far_5_5890_0_b(.in(layer_4[77]), .out(far_5_5890_0[1]));
    assign layer_5[790] = far_5_5890_0[0] ^ far_5_5890_0[1]; 
    wire [1:0] far_5_5891_0;    relay_conn far_5_5891_0_a(.in(layer_4[172]), .out(far_5_5891_0[0]));    relay_conn far_5_5891_0_b(.in(layer_4[300]), .out(far_5_5891_0[1]));
    wire [1:0] far_5_5891_1;    relay_conn far_5_5891_1_a(.in(far_5_5891_0[0]), .out(far_5_5891_1[0]));    relay_conn far_5_5891_1_b(.in(far_5_5891_0[1]), .out(far_5_5891_1[1]));
    wire [1:0] far_5_5891_2;    relay_conn far_5_5891_2_a(.in(far_5_5891_1[0]), .out(far_5_5891_2[0]));    relay_conn far_5_5891_2_b(.in(far_5_5891_1[1]), .out(far_5_5891_2[1]));
    wire [1:0] far_5_5891_3;    relay_conn far_5_5891_3_a(.in(far_5_5891_2[0]), .out(far_5_5891_3[0]));    relay_conn far_5_5891_3_b(.in(far_5_5891_2[1]), .out(far_5_5891_3[1]));
    assign layer_5[791] = far_5_5891_3[1] & ~far_5_5891_3[0]; 
    wire [1:0] far_5_5892_0;    relay_conn far_5_5892_0_a(.in(layer_4[443]), .out(far_5_5892_0[0]));    relay_conn far_5_5892_0_b(.in(layer_4[520]), .out(far_5_5892_0[1]));
    wire [1:0] far_5_5892_1;    relay_conn far_5_5892_1_a(.in(far_5_5892_0[0]), .out(far_5_5892_1[0]));    relay_conn far_5_5892_1_b(.in(far_5_5892_0[1]), .out(far_5_5892_1[1]));
    assign layer_5[792] = far_5_5892_1[0] & far_5_5892_1[1]; 
    assign layer_5[793] = ~layer_4[885]; 
    wire [1:0] far_5_5894_0;    relay_conn far_5_5894_0_a(.in(layer_4[807]), .out(far_5_5894_0[0]));    relay_conn far_5_5894_0_b(.in(layer_4[905]), .out(far_5_5894_0[1]));
    wire [1:0] far_5_5894_1;    relay_conn far_5_5894_1_a(.in(far_5_5894_0[0]), .out(far_5_5894_1[0]));    relay_conn far_5_5894_1_b(.in(far_5_5894_0[1]), .out(far_5_5894_1[1]));
    wire [1:0] far_5_5894_2;    relay_conn far_5_5894_2_a(.in(far_5_5894_1[0]), .out(far_5_5894_2[0]));    relay_conn far_5_5894_2_b(.in(far_5_5894_1[1]), .out(far_5_5894_2[1]));
    assign layer_5[794] = far_5_5894_2[1] & ~far_5_5894_2[0]; 
    wire [1:0] far_5_5895_0;    relay_conn far_5_5895_0_a(.in(layer_4[653]), .out(far_5_5895_0[0]));    relay_conn far_5_5895_0_b(.in(layer_4[620]), .out(far_5_5895_0[1]));
    assign layer_5[795] = ~far_5_5895_0[1]; 
    assign layer_5[796] = ~layer_4[642] | (layer_4[642] & layer_4[665]); 
    wire [1:0] far_5_5897_0;    relay_conn far_5_5897_0_a(.in(layer_4[576]), .out(far_5_5897_0[0]));    relay_conn far_5_5897_0_b(.in(layer_4[630]), .out(far_5_5897_0[1]));
    assign layer_5[797] = ~(far_5_5897_0[0] & far_5_5897_0[1]); 
    assign layer_5[798] = layer_4[1003] & layer_4[1019]; 
    wire [1:0] far_5_5899_0;    relay_conn far_5_5899_0_a(.in(layer_4[1001]), .out(far_5_5899_0[0]));    relay_conn far_5_5899_0_b(.in(layer_4[902]), .out(far_5_5899_0[1]));
    wire [1:0] far_5_5899_1;    relay_conn far_5_5899_1_a(.in(far_5_5899_0[0]), .out(far_5_5899_1[0]));    relay_conn far_5_5899_1_b(.in(far_5_5899_0[1]), .out(far_5_5899_1[1]));
    wire [1:0] far_5_5899_2;    relay_conn far_5_5899_2_a(.in(far_5_5899_1[0]), .out(far_5_5899_2[0]));    relay_conn far_5_5899_2_b(.in(far_5_5899_1[1]), .out(far_5_5899_2[1]));
    assign layer_5[799] = far_5_5899_2[0] & ~far_5_5899_2[1]; 
    wire [1:0] far_5_5900_0;    relay_conn far_5_5900_0_a(.in(layer_4[938]), .out(far_5_5900_0[0]));    relay_conn far_5_5900_0_b(.in(layer_4[876]), .out(far_5_5900_0[1]));
    assign layer_5[800] = far_5_5900_0[0] | far_5_5900_0[1]; 
    wire [1:0] far_5_5901_0;    relay_conn far_5_5901_0_a(.in(layer_4[980]), .out(far_5_5901_0[0]));    relay_conn far_5_5901_0_b(.in(layer_4[875]), .out(far_5_5901_0[1]));
    wire [1:0] far_5_5901_1;    relay_conn far_5_5901_1_a(.in(far_5_5901_0[0]), .out(far_5_5901_1[0]));    relay_conn far_5_5901_1_b(.in(far_5_5901_0[1]), .out(far_5_5901_1[1]));
    wire [1:0] far_5_5901_2;    relay_conn far_5_5901_2_a(.in(far_5_5901_1[0]), .out(far_5_5901_2[0]));    relay_conn far_5_5901_2_b(.in(far_5_5901_1[1]), .out(far_5_5901_2[1]));
    assign layer_5[801] = ~(far_5_5901_2[0] | far_5_5901_2[1]); 
    assign layer_5[802] = ~(layer_4[656] & layer_4[665]); 
    assign layer_5[803] = layer_4[89]; 
    wire [1:0] far_5_5904_0;    relay_conn far_5_5904_0_a(.in(layer_4[397]), .out(far_5_5904_0[0]));    relay_conn far_5_5904_0_b(.in(layer_4[511]), .out(far_5_5904_0[1]));
    wire [1:0] far_5_5904_1;    relay_conn far_5_5904_1_a(.in(far_5_5904_0[0]), .out(far_5_5904_1[0]));    relay_conn far_5_5904_1_b(.in(far_5_5904_0[1]), .out(far_5_5904_1[1]));
    wire [1:0] far_5_5904_2;    relay_conn far_5_5904_2_a(.in(far_5_5904_1[0]), .out(far_5_5904_2[0]));    relay_conn far_5_5904_2_b(.in(far_5_5904_1[1]), .out(far_5_5904_2[1]));
    assign layer_5[804] = ~far_5_5904_2[0] | (far_5_5904_2[0] & far_5_5904_2[1]); 
    wire [1:0] far_5_5905_0;    relay_conn far_5_5905_0_a(.in(layer_4[39]), .out(far_5_5905_0[0]));    relay_conn far_5_5905_0_b(.in(layer_4[158]), .out(far_5_5905_0[1]));
    wire [1:0] far_5_5905_1;    relay_conn far_5_5905_1_a(.in(far_5_5905_0[0]), .out(far_5_5905_1[0]));    relay_conn far_5_5905_1_b(.in(far_5_5905_0[1]), .out(far_5_5905_1[1]));
    wire [1:0] far_5_5905_2;    relay_conn far_5_5905_2_a(.in(far_5_5905_1[0]), .out(far_5_5905_2[0]));    relay_conn far_5_5905_2_b(.in(far_5_5905_1[1]), .out(far_5_5905_2[1]));
    assign layer_5[805] = far_5_5905_2[1]; 
    wire [1:0] far_5_5906_0;    relay_conn far_5_5906_0_a(.in(layer_4[331]), .out(far_5_5906_0[0]));    relay_conn far_5_5906_0_b(.in(layer_4[275]), .out(far_5_5906_0[1]));
    assign layer_5[806] = ~(far_5_5906_0[0] & far_5_5906_0[1]); 
    assign layer_5[807] = ~(layer_4[421] | layer_4[397]); 
    wire [1:0] far_5_5908_0;    relay_conn far_5_5908_0_a(.in(layer_4[15]), .out(far_5_5908_0[0]));    relay_conn far_5_5908_0_b(.in(layer_4[89]), .out(far_5_5908_0[1]));
    wire [1:0] far_5_5908_1;    relay_conn far_5_5908_1_a(.in(far_5_5908_0[0]), .out(far_5_5908_1[0]));    relay_conn far_5_5908_1_b(.in(far_5_5908_0[1]), .out(far_5_5908_1[1]));
    assign layer_5[808] = far_5_5908_1[0] & ~far_5_5908_1[1]; 
    wire [1:0] far_5_5909_0;    relay_conn far_5_5909_0_a(.in(layer_4[768]), .out(far_5_5909_0[0]));    relay_conn far_5_5909_0_b(.in(layer_4[866]), .out(far_5_5909_0[1]));
    wire [1:0] far_5_5909_1;    relay_conn far_5_5909_1_a(.in(far_5_5909_0[0]), .out(far_5_5909_1[0]));    relay_conn far_5_5909_1_b(.in(far_5_5909_0[1]), .out(far_5_5909_1[1]));
    wire [1:0] far_5_5909_2;    relay_conn far_5_5909_2_a(.in(far_5_5909_1[0]), .out(far_5_5909_2[0]));    relay_conn far_5_5909_2_b(.in(far_5_5909_1[1]), .out(far_5_5909_2[1]));
    assign layer_5[809] = ~(far_5_5909_2[0] | far_5_5909_2[1]); 
    assign layer_5[810] = layer_4[593] | layer_4[595]; 
    wire [1:0] far_5_5911_0;    relay_conn far_5_5911_0_a(.in(layer_4[309]), .out(far_5_5911_0[0]));    relay_conn far_5_5911_0_b(.in(layer_4[188]), .out(far_5_5911_0[1]));
    wire [1:0] far_5_5911_1;    relay_conn far_5_5911_1_a(.in(far_5_5911_0[0]), .out(far_5_5911_1[0]));    relay_conn far_5_5911_1_b(.in(far_5_5911_0[1]), .out(far_5_5911_1[1]));
    wire [1:0] far_5_5911_2;    relay_conn far_5_5911_2_a(.in(far_5_5911_1[0]), .out(far_5_5911_2[0]));    relay_conn far_5_5911_2_b(.in(far_5_5911_1[1]), .out(far_5_5911_2[1]));
    assign layer_5[811] = ~far_5_5911_2[1]; 
    wire [1:0] far_5_5912_0;    relay_conn far_5_5912_0_a(.in(layer_4[402]), .out(far_5_5912_0[0]));    relay_conn far_5_5912_0_b(.in(layer_4[443]), .out(far_5_5912_0[1]));
    assign layer_5[812] = ~far_5_5912_0[0] | (far_5_5912_0[0] & far_5_5912_0[1]); 
    assign layer_5[813] = ~(layer_4[16] & layer_4[28]); 
    assign layer_5[814] = layer_4[263]; 
    wire [1:0] far_5_5915_0;    relay_conn far_5_5915_0_a(.in(layer_4[29]), .out(far_5_5915_0[0]));    relay_conn far_5_5915_0_b(.in(layer_4[133]), .out(far_5_5915_0[1]));
    wire [1:0] far_5_5915_1;    relay_conn far_5_5915_1_a(.in(far_5_5915_0[0]), .out(far_5_5915_1[0]));    relay_conn far_5_5915_1_b(.in(far_5_5915_0[1]), .out(far_5_5915_1[1]));
    wire [1:0] far_5_5915_2;    relay_conn far_5_5915_2_a(.in(far_5_5915_1[0]), .out(far_5_5915_2[0]));    relay_conn far_5_5915_2_b(.in(far_5_5915_1[1]), .out(far_5_5915_2[1]));
    assign layer_5[815] = ~(far_5_5915_2[0] & far_5_5915_2[1]); 
    wire [1:0] far_5_5916_0;    relay_conn far_5_5916_0_a(.in(layer_4[253]), .out(far_5_5916_0[0]));    relay_conn far_5_5916_0_b(.in(layer_4[363]), .out(far_5_5916_0[1]));
    wire [1:0] far_5_5916_1;    relay_conn far_5_5916_1_a(.in(far_5_5916_0[0]), .out(far_5_5916_1[0]));    relay_conn far_5_5916_1_b(.in(far_5_5916_0[1]), .out(far_5_5916_1[1]));
    wire [1:0] far_5_5916_2;    relay_conn far_5_5916_2_a(.in(far_5_5916_1[0]), .out(far_5_5916_2[0]));    relay_conn far_5_5916_2_b(.in(far_5_5916_1[1]), .out(far_5_5916_2[1]));
    assign layer_5[816] = far_5_5916_2[0]; 
    wire [1:0] far_5_5917_0;    relay_conn far_5_5917_0_a(.in(layer_4[650]), .out(far_5_5917_0[0]));    relay_conn far_5_5917_0_b(.in(layer_4[553]), .out(far_5_5917_0[1]));
    wire [1:0] far_5_5917_1;    relay_conn far_5_5917_1_a(.in(far_5_5917_0[0]), .out(far_5_5917_1[0]));    relay_conn far_5_5917_1_b(.in(far_5_5917_0[1]), .out(far_5_5917_1[1]));
    wire [1:0] far_5_5917_2;    relay_conn far_5_5917_2_a(.in(far_5_5917_1[0]), .out(far_5_5917_2[0]));    relay_conn far_5_5917_2_b(.in(far_5_5917_1[1]), .out(far_5_5917_2[1]));
    assign layer_5[817] = ~far_5_5917_2[0] | (far_5_5917_2[0] & far_5_5917_2[1]); 
    assign layer_5[818] = layer_4[307] & layer_4[294]; 
    wire [1:0] far_5_5919_0;    relay_conn far_5_5919_0_a(.in(layer_4[904]), .out(far_5_5919_0[0]));    relay_conn far_5_5919_0_b(.in(layer_4[858]), .out(far_5_5919_0[1]));
    assign layer_5[819] = far_5_5919_0[0] ^ far_5_5919_0[1]; 
    wire [1:0] far_5_5920_0;    relay_conn far_5_5920_0_a(.in(layer_4[217]), .out(far_5_5920_0[0]));    relay_conn far_5_5920_0_b(.in(layer_4[289]), .out(far_5_5920_0[1]));
    wire [1:0] far_5_5920_1;    relay_conn far_5_5920_1_a(.in(far_5_5920_0[0]), .out(far_5_5920_1[0]));    relay_conn far_5_5920_1_b(.in(far_5_5920_0[1]), .out(far_5_5920_1[1]));
    assign layer_5[820] = far_5_5920_1[1] & ~far_5_5920_1[0]; 
    wire [1:0] far_5_5921_0;    relay_conn far_5_5921_0_a(.in(layer_4[597]), .out(far_5_5921_0[0]));    relay_conn far_5_5921_0_b(.in(layer_4[719]), .out(far_5_5921_0[1]));
    wire [1:0] far_5_5921_1;    relay_conn far_5_5921_1_a(.in(far_5_5921_0[0]), .out(far_5_5921_1[0]));    relay_conn far_5_5921_1_b(.in(far_5_5921_0[1]), .out(far_5_5921_1[1]));
    wire [1:0] far_5_5921_2;    relay_conn far_5_5921_2_a(.in(far_5_5921_1[0]), .out(far_5_5921_2[0]));    relay_conn far_5_5921_2_b(.in(far_5_5921_1[1]), .out(far_5_5921_2[1]));
    assign layer_5[821] = far_5_5921_2[0] ^ far_5_5921_2[1]; 
    assign layer_5[822] = ~(layer_4[200] | layer_4[171]); 
    assign layer_5[823] = layer_4[656]; 
    wire [1:0] far_5_5924_0;    relay_conn far_5_5924_0_a(.in(layer_4[202]), .out(far_5_5924_0[0]));    relay_conn far_5_5924_0_b(.in(layer_4[94]), .out(far_5_5924_0[1]));
    wire [1:0] far_5_5924_1;    relay_conn far_5_5924_1_a(.in(far_5_5924_0[0]), .out(far_5_5924_1[0]));    relay_conn far_5_5924_1_b(.in(far_5_5924_0[1]), .out(far_5_5924_1[1]));
    wire [1:0] far_5_5924_2;    relay_conn far_5_5924_2_a(.in(far_5_5924_1[0]), .out(far_5_5924_2[0]));    relay_conn far_5_5924_2_b(.in(far_5_5924_1[1]), .out(far_5_5924_2[1]));
    assign layer_5[824] = far_5_5924_2[0] & ~far_5_5924_2[1]; 
    wire [1:0] far_5_5925_0;    relay_conn far_5_5925_0_a(.in(layer_4[238]), .out(far_5_5925_0[0]));    relay_conn far_5_5925_0_b(.in(layer_4[190]), .out(far_5_5925_0[1]));
    assign layer_5[825] = far_5_5925_0[0]; 
    assign layer_5[826] = layer_4[983]; 
    wire [1:0] far_5_5927_0;    relay_conn far_5_5927_0_a(.in(layer_4[605]), .out(far_5_5927_0[0]));    relay_conn far_5_5927_0_b(.in(layer_4[719]), .out(far_5_5927_0[1]));
    wire [1:0] far_5_5927_1;    relay_conn far_5_5927_1_a(.in(far_5_5927_0[0]), .out(far_5_5927_1[0]));    relay_conn far_5_5927_1_b(.in(far_5_5927_0[1]), .out(far_5_5927_1[1]));
    wire [1:0] far_5_5927_2;    relay_conn far_5_5927_2_a(.in(far_5_5927_1[0]), .out(far_5_5927_2[0]));    relay_conn far_5_5927_2_b(.in(far_5_5927_1[1]), .out(far_5_5927_2[1]));
    assign layer_5[827] = far_5_5927_2[0] | far_5_5927_2[1]; 
    wire [1:0] far_5_5928_0;    relay_conn far_5_5928_0_a(.in(layer_4[425]), .out(far_5_5928_0[0]));    relay_conn far_5_5928_0_b(.in(layer_4[389]), .out(far_5_5928_0[1]));
    assign layer_5[828] = far_5_5928_0[0] & far_5_5928_0[1]; 
    wire [1:0] far_5_5929_0;    relay_conn far_5_5929_0_a(.in(layer_4[760]), .out(far_5_5929_0[0]));    relay_conn far_5_5929_0_b(.in(layer_4[860]), .out(far_5_5929_0[1]));
    wire [1:0] far_5_5929_1;    relay_conn far_5_5929_1_a(.in(far_5_5929_0[0]), .out(far_5_5929_1[0]));    relay_conn far_5_5929_1_b(.in(far_5_5929_0[1]), .out(far_5_5929_1[1]));
    wire [1:0] far_5_5929_2;    relay_conn far_5_5929_2_a(.in(far_5_5929_1[0]), .out(far_5_5929_2[0]));    relay_conn far_5_5929_2_b(.in(far_5_5929_1[1]), .out(far_5_5929_2[1]));
    assign layer_5[829] = ~(far_5_5929_2[0] ^ far_5_5929_2[1]); 
    assign layer_5[830] = ~(layer_4[719] | layer_4[704]); 
    assign layer_5[831] = layer_4[150] & layer_4[133]; 
    assign layer_5[832] = ~layer_4[167] | (layer_4[167] & layer_4[198]); 
    wire [1:0] far_5_5933_0;    relay_conn far_5_5933_0_a(.in(layer_4[534]), .out(far_5_5933_0[0]));    relay_conn far_5_5933_0_b(.in(layer_4[416]), .out(far_5_5933_0[1]));
    wire [1:0] far_5_5933_1;    relay_conn far_5_5933_1_a(.in(far_5_5933_0[0]), .out(far_5_5933_1[0]));    relay_conn far_5_5933_1_b(.in(far_5_5933_0[1]), .out(far_5_5933_1[1]));
    wire [1:0] far_5_5933_2;    relay_conn far_5_5933_2_a(.in(far_5_5933_1[0]), .out(far_5_5933_2[0]));    relay_conn far_5_5933_2_b(.in(far_5_5933_1[1]), .out(far_5_5933_2[1]));
    assign layer_5[833] = ~(far_5_5933_2[0] & far_5_5933_2[1]); 
    wire [1:0] far_5_5934_0;    relay_conn far_5_5934_0_a(.in(layer_4[830]), .out(far_5_5934_0[0]));    relay_conn far_5_5934_0_b(.in(layer_4[712]), .out(far_5_5934_0[1]));
    wire [1:0] far_5_5934_1;    relay_conn far_5_5934_1_a(.in(far_5_5934_0[0]), .out(far_5_5934_1[0]));    relay_conn far_5_5934_1_b(.in(far_5_5934_0[1]), .out(far_5_5934_1[1]));
    wire [1:0] far_5_5934_2;    relay_conn far_5_5934_2_a(.in(far_5_5934_1[0]), .out(far_5_5934_2[0]));    relay_conn far_5_5934_2_b(.in(far_5_5934_1[1]), .out(far_5_5934_2[1]));
    assign layer_5[834] = ~(far_5_5934_2[0] | far_5_5934_2[1]); 
    wire [1:0] far_5_5935_0;    relay_conn far_5_5935_0_a(.in(layer_4[571]), .out(far_5_5935_0[0]));    relay_conn far_5_5935_0_b(.in(layer_4[453]), .out(far_5_5935_0[1]));
    wire [1:0] far_5_5935_1;    relay_conn far_5_5935_1_a(.in(far_5_5935_0[0]), .out(far_5_5935_1[0]));    relay_conn far_5_5935_1_b(.in(far_5_5935_0[1]), .out(far_5_5935_1[1]));
    wire [1:0] far_5_5935_2;    relay_conn far_5_5935_2_a(.in(far_5_5935_1[0]), .out(far_5_5935_2[0]));    relay_conn far_5_5935_2_b(.in(far_5_5935_1[1]), .out(far_5_5935_2[1]));
    assign layer_5[835] = ~far_5_5935_2[1]; 
    wire [1:0] far_5_5936_0;    relay_conn far_5_5936_0_a(.in(layer_4[900]), .out(far_5_5936_0[0]));    relay_conn far_5_5936_0_b(.in(layer_4[850]), .out(far_5_5936_0[1]));
    assign layer_5[836] = far_5_5936_0[1] & ~far_5_5936_0[0]; 
    assign layer_5[837] = ~layer_4[970]; 
    wire [1:0] far_5_5938_0;    relay_conn far_5_5938_0_a(.in(layer_4[395]), .out(far_5_5938_0[0]));    relay_conn far_5_5938_0_b(.in(layer_4[429]), .out(far_5_5938_0[1]));
    assign layer_5[838] = far_5_5938_0[0] | far_5_5938_0[1]; 
    wire [1:0] far_5_5939_0;    relay_conn far_5_5939_0_a(.in(layer_4[516]), .out(far_5_5939_0[0]));    relay_conn far_5_5939_0_b(.in(layer_4[638]), .out(far_5_5939_0[1]));
    wire [1:0] far_5_5939_1;    relay_conn far_5_5939_1_a(.in(far_5_5939_0[0]), .out(far_5_5939_1[0]));    relay_conn far_5_5939_1_b(.in(far_5_5939_0[1]), .out(far_5_5939_1[1]));
    wire [1:0] far_5_5939_2;    relay_conn far_5_5939_2_a(.in(far_5_5939_1[0]), .out(far_5_5939_2[0]));    relay_conn far_5_5939_2_b(.in(far_5_5939_1[1]), .out(far_5_5939_2[1]));
    assign layer_5[839] = ~(far_5_5939_2[0] | far_5_5939_2[1]); 
    assign layer_5[840] = ~(layer_4[65] | layer_4[42]); 
    wire [1:0] far_5_5941_0;    relay_conn far_5_5941_0_a(.in(layer_4[576]), .out(far_5_5941_0[0]));    relay_conn far_5_5941_0_b(.in(layer_4[650]), .out(far_5_5941_0[1]));
    wire [1:0] far_5_5941_1;    relay_conn far_5_5941_1_a(.in(far_5_5941_0[0]), .out(far_5_5941_1[0]));    relay_conn far_5_5941_1_b(.in(far_5_5941_0[1]), .out(far_5_5941_1[1]));
    assign layer_5[841] = ~far_5_5941_1[1]; 
    wire [1:0] far_5_5942_0;    relay_conn far_5_5942_0_a(.in(layer_4[268]), .out(far_5_5942_0[0]));    relay_conn far_5_5942_0_b(.in(layer_4[222]), .out(far_5_5942_0[1]));
    assign layer_5[842] = ~far_5_5942_0[1] | (far_5_5942_0[0] & far_5_5942_0[1]); 
    assign layer_5[843] = layer_4[187] | layer_4[199]; 
    wire [1:0] far_5_5944_0;    relay_conn far_5_5944_0_a(.in(layer_4[505]), .out(far_5_5944_0[0]));    relay_conn far_5_5944_0_b(.in(layer_4[423]), .out(far_5_5944_0[1]));
    wire [1:0] far_5_5944_1;    relay_conn far_5_5944_1_a(.in(far_5_5944_0[0]), .out(far_5_5944_1[0]));    relay_conn far_5_5944_1_b(.in(far_5_5944_0[1]), .out(far_5_5944_1[1]));
    assign layer_5[844] = far_5_5944_1[1]; 
    wire [1:0] far_5_5945_0;    relay_conn far_5_5945_0_a(.in(layer_4[620]), .out(far_5_5945_0[0]));    relay_conn far_5_5945_0_b(.in(layer_4[568]), .out(far_5_5945_0[1]));
    assign layer_5[845] = far_5_5945_0[0] & ~far_5_5945_0[1]; 
    wire [1:0] far_5_5946_0;    relay_conn far_5_5946_0_a(.in(layer_4[84]), .out(far_5_5946_0[0]));    relay_conn far_5_5946_0_b(.in(layer_4[9]), .out(far_5_5946_0[1]));
    wire [1:0] far_5_5946_1;    relay_conn far_5_5946_1_a(.in(far_5_5946_0[0]), .out(far_5_5946_1[0]));    relay_conn far_5_5946_1_b(.in(far_5_5946_0[1]), .out(far_5_5946_1[1]));
    assign layer_5[846] = far_5_5946_1[0]; 
    wire [1:0] far_5_5947_0;    relay_conn far_5_5947_0_a(.in(layer_4[995]), .out(far_5_5947_0[0]));    relay_conn far_5_5947_0_b(.in(layer_4[910]), .out(far_5_5947_0[1]));
    wire [1:0] far_5_5947_1;    relay_conn far_5_5947_1_a(.in(far_5_5947_0[0]), .out(far_5_5947_1[0]));    relay_conn far_5_5947_1_b(.in(far_5_5947_0[1]), .out(far_5_5947_1[1]));
    assign layer_5[847] = ~far_5_5947_1[1] | (far_5_5947_1[0] & far_5_5947_1[1]); 
    assign layer_5[848] = layer_4[888] ^ layer_4[904]; 
    wire [1:0] far_5_5949_0;    relay_conn far_5_5949_0_a(.in(layer_4[855]), .out(far_5_5949_0[0]));    relay_conn far_5_5949_0_b(.in(layer_4[970]), .out(far_5_5949_0[1]));
    wire [1:0] far_5_5949_1;    relay_conn far_5_5949_1_a(.in(far_5_5949_0[0]), .out(far_5_5949_1[0]));    relay_conn far_5_5949_1_b(.in(far_5_5949_0[1]), .out(far_5_5949_1[1]));
    wire [1:0] far_5_5949_2;    relay_conn far_5_5949_2_a(.in(far_5_5949_1[0]), .out(far_5_5949_2[0]));    relay_conn far_5_5949_2_b(.in(far_5_5949_1[1]), .out(far_5_5949_2[1]));
    assign layer_5[849] = far_5_5949_2[0]; 
    assign layer_5[850] = ~(layer_4[436] & layer_4[420]); 
    assign layer_5[851] = ~layer_4[466] | (layer_4[439] & layer_4[466]); 
    assign layer_5[852] = layer_4[871] & ~layer_4[898]; 
    wire [1:0] far_5_5953_0;    relay_conn far_5_5953_0_a(.in(layer_4[630]), .out(far_5_5953_0[0]));    relay_conn far_5_5953_0_b(.in(layer_4[692]), .out(far_5_5953_0[1]));
    assign layer_5[853] = far_5_5953_0[1]; 
    wire [1:0] far_5_5954_0;    relay_conn far_5_5954_0_a(.in(layer_4[953]), .out(far_5_5954_0[0]));    relay_conn far_5_5954_0_b(.in(layer_4[827]), .out(far_5_5954_0[1]));
    wire [1:0] far_5_5954_1;    relay_conn far_5_5954_1_a(.in(far_5_5954_0[0]), .out(far_5_5954_1[0]));    relay_conn far_5_5954_1_b(.in(far_5_5954_0[1]), .out(far_5_5954_1[1]));
    wire [1:0] far_5_5954_2;    relay_conn far_5_5954_2_a(.in(far_5_5954_1[0]), .out(far_5_5954_2[0]));    relay_conn far_5_5954_2_b(.in(far_5_5954_1[1]), .out(far_5_5954_2[1]));
    assign layer_5[854] = far_5_5954_2[1]; 
    wire [1:0] far_5_5955_0;    relay_conn far_5_5955_0_a(.in(layer_4[617]), .out(far_5_5955_0[0]));    relay_conn far_5_5955_0_b(.in(layer_4[544]), .out(far_5_5955_0[1]));
    wire [1:0] far_5_5955_1;    relay_conn far_5_5955_1_a(.in(far_5_5955_0[0]), .out(far_5_5955_1[0]));    relay_conn far_5_5955_1_b(.in(far_5_5955_0[1]), .out(far_5_5955_1[1]));
    assign layer_5[855] = far_5_5955_1[0] | far_5_5955_1[1]; 
    wire [1:0] far_5_5956_0;    relay_conn far_5_5956_0_a(.in(layer_4[767]), .out(far_5_5956_0[0]));    relay_conn far_5_5956_0_b(.in(layer_4[826]), .out(far_5_5956_0[1]));
    assign layer_5[856] = ~far_5_5956_0[0]; 
    wire [1:0] far_5_5957_0;    relay_conn far_5_5957_0_a(.in(layer_4[900]), .out(far_5_5957_0[0]));    relay_conn far_5_5957_0_b(.in(layer_4[854]), .out(far_5_5957_0[1]));
    assign layer_5[857] = ~far_5_5957_0[1] | (far_5_5957_0[0] & far_5_5957_0[1]); 
    wire [1:0] far_5_5958_0;    relay_conn far_5_5958_0_a(.in(layer_4[651]), .out(far_5_5958_0[0]));    relay_conn far_5_5958_0_b(.in(layer_4[707]), .out(far_5_5958_0[1]));
    assign layer_5[858] = far_5_5958_0[0] | far_5_5958_0[1]; 
    wire [1:0] far_5_5959_0;    relay_conn far_5_5959_0_a(.in(layer_4[858]), .out(far_5_5959_0[0]));    relay_conn far_5_5959_0_b(.in(layer_4[795]), .out(far_5_5959_0[1]));
    assign layer_5[859] = ~(far_5_5959_0[0] | far_5_5959_0[1]); 
    wire [1:0] far_5_5960_0;    relay_conn far_5_5960_0_a(.in(layer_4[377]), .out(far_5_5960_0[0]));    relay_conn far_5_5960_0_b(.in(layer_4[497]), .out(far_5_5960_0[1]));
    wire [1:0] far_5_5960_1;    relay_conn far_5_5960_1_a(.in(far_5_5960_0[0]), .out(far_5_5960_1[0]));    relay_conn far_5_5960_1_b(.in(far_5_5960_0[1]), .out(far_5_5960_1[1]));
    wire [1:0] far_5_5960_2;    relay_conn far_5_5960_2_a(.in(far_5_5960_1[0]), .out(far_5_5960_2[0]));    relay_conn far_5_5960_2_b(.in(far_5_5960_1[1]), .out(far_5_5960_2[1]));
    assign layer_5[860] = ~far_5_5960_2[1]; 
    wire [1:0] far_5_5961_0;    relay_conn far_5_5961_0_a(.in(layer_4[217]), .out(far_5_5961_0[0]));    relay_conn far_5_5961_0_b(.in(layer_4[271]), .out(far_5_5961_0[1]));
    assign layer_5[861] = ~far_5_5961_0[1]; 
    wire [1:0] far_5_5962_0;    relay_conn far_5_5962_0_a(.in(layer_4[1015]), .out(far_5_5962_0[0]));    relay_conn far_5_5962_0_b(.in(layer_4[947]), .out(far_5_5962_0[1]));
    wire [1:0] far_5_5962_1;    relay_conn far_5_5962_1_a(.in(far_5_5962_0[0]), .out(far_5_5962_1[0]));    relay_conn far_5_5962_1_b(.in(far_5_5962_0[1]), .out(far_5_5962_1[1]));
    assign layer_5[862] = ~(far_5_5962_1[0] ^ far_5_5962_1[1]); 
    wire [1:0] far_5_5963_0;    relay_conn far_5_5963_0_a(.in(layer_4[23]), .out(far_5_5963_0[0]));    relay_conn far_5_5963_0_b(.in(layer_4[133]), .out(far_5_5963_0[1]));
    wire [1:0] far_5_5963_1;    relay_conn far_5_5963_1_a(.in(far_5_5963_0[0]), .out(far_5_5963_1[0]));    relay_conn far_5_5963_1_b(.in(far_5_5963_0[1]), .out(far_5_5963_1[1]));
    wire [1:0] far_5_5963_2;    relay_conn far_5_5963_2_a(.in(far_5_5963_1[0]), .out(far_5_5963_2[0]));    relay_conn far_5_5963_2_b(.in(far_5_5963_1[1]), .out(far_5_5963_2[1]));
    assign layer_5[863] = ~far_5_5963_2[0]; 
    wire [1:0] far_5_5964_0;    relay_conn far_5_5964_0_a(.in(layer_4[153]), .out(far_5_5964_0[0]));    relay_conn far_5_5964_0_b(.in(layer_4[66]), .out(far_5_5964_0[1]));
    wire [1:0] far_5_5964_1;    relay_conn far_5_5964_1_a(.in(far_5_5964_0[0]), .out(far_5_5964_1[0]));    relay_conn far_5_5964_1_b(.in(far_5_5964_0[1]), .out(far_5_5964_1[1]));
    assign layer_5[864] = far_5_5964_1[1] & ~far_5_5964_1[0]; 
    wire [1:0] far_5_5965_0;    relay_conn far_5_5965_0_a(.in(layer_4[127]), .out(far_5_5965_0[0]));    relay_conn far_5_5965_0_b(.in(layer_4[232]), .out(far_5_5965_0[1]));
    wire [1:0] far_5_5965_1;    relay_conn far_5_5965_1_a(.in(far_5_5965_0[0]), .out(far_5_5965_1[0]));    relay_conn far_5_5965_1_b(.in(far_5_5965_0[1]), .out(far_5_5965_1[1]));
    wire [1:0] far_5_5965_2;    relay_conn far_5_5965_2_a(.in(far_5_5965_1[0]), .out(far_5_5965_2[0]));    relay_conn far_5_5965_2_b(.in(far_5_5965_1[1]), .out(far_5_5965_2[1]));
    assign layer_5[865] = ~far_5_5965_2[1]; 
    wire [1:0] far_5_5966_0;    relay_conn far_5_5966_0_a(.in(layer_4[190]), .out(far_5_5966_0[0]));    relay_conn far_5_5966_0_b(.in(layer_4[103]), .out(far_5_5966_0[1]));
    wire [1:0] far_5_5966_1;    relay_conn far_5_5966_1_a(.in(far_5_5966_0[0]), .out(far_5_5966_1[0]));    relay_conn far_5_5966_1_b(.in(far_5_5966_0[1]), .out(far_5_5966_1[1]));
    assign layer_5[866] = ~far_5_5966_1[0] | (far_5_5966_1[0] & far_5_5966_1[1]); 
    wire [1:0] far_5_5967_0;    relay_conn far_5_5967_0_a(.in(layer_4[307]), .out(far_5_5967_0[0]));    relay_conn far_5_5967_0_b(.in(layer_4[392]), .out(far_5_5967_0[1]));
    wire [1:0] far_5_5967_1;    relay_conn far_5_5967_1_a(.in(far_5_5967_0[0]), .out(far_5_5967_1[0]));    relay_conn far_5_5967_1_b(.in(far_5_5967_0[1]), .out(far_5_5967_1[1]));
    assign layer_5[867] = far_5_5967_1[0]; 
    wire [1:0] far_5_5968_0;    relay_conn far_5_5968_0_a(.in(layer_4[423]), .out(far_5_5968_0[0]));    relay_conn far_5_5968_0_b(.in(layer_4[545]), .out(far_5_5968_0[1]));
    wire [1:0] far_5_5968_1;    relay_conn far_5_5968_1_a(.in(far_5_5968_0[0]), .out(far_5_5968_1[0]));    relay_conn far_5_5968_1_b(.in(far_5_5968_0[1]), .out(far_5_5968_1[1]));
    wire [1:0] far_5_5968_2;    relay_conn far_5_5968_2_a(.in(far_5_5968_1[0]), .out(far_5_5968_2[0]));    relay_conn far_5_5968_2_b(.in(far_5_5968_1[1]), .out(far_5_5968_2[1]));
    assign layer_5[868] = ~far_5_5968_2[1] | (far_5_5968_2[0] & far_5_5968_2[1]); 
    wire [1:0] far_5_5969_0;    relay_conn far_5_5969_0_a(.in(layer_4[617]), .out(far_5_5969_0[0]));    relay_conn far_5_5969_0_b(.in(layer_4[656]), .out(far_5_5969_0[1]));
    assign layer_5[869] = far_5_5969_0[0] & ~far_5_5969_0[1]; 
    wire [1:0] far_5_5970_0;    relay_conn far_5_5970_0_a(.in(layer_4[177]), .out(far_5_5970_0[0]));    relay_conn far_5_5970_0_b(.in(layer_4[295]), .out(far_5_5970_0[1]));
    wire [1:0] far_5_5970_1;    relay_conn far_5_5970_1_a(.in(far_5_5970_0[0]), .out(far_5_5970_1[0]));    relay_conn far_5_5970_1_b(.in(far_5_5970_0[1]), .out(far_5_5970_1[1]));
    wire [1:0] far_5_5970_2;    relay_conn far_5_5970_2_a(.in(far_5_5970_1[0]), .out(far_5_5970_2[0]));    relay_conn far_5_5970_2_b(.in(far_5_5970_1[1]), .out(far_5_5970_2[1]));
    assign layer_5[870] = ~far_5_5970_2[0] | (far_5_5970_2[0] & far_5_5970_2[1]); 
    wire [1:0] far_5_5971_0;    relay_conn far_5_5971_0_a(.in(layer_4[224]), .out(far_5_5971_0[0]));    relay_conn far_5_5971_0_b(.in(layer_4[118]), .out(far_5_5971_0[1]));
    wire [1:0] far_5_5971_1;    relay_conn far_5_5971_1_a(.in(far_5_5971_0[0]), .out(far_5_5971_1[0]));    relay_conn far_5_5971_1_b(.in(far_5_5971_0[1]), .out(far_5_5971_1[1]));
    wire [1:0] far_5_5971_2;    relay_conn far_5_5971_2_a(.in(far_5_5971_1[0]), .out(far_5_5971_2[0]));    relay_conn far_5_5971_2_b(.in(far_5_5971_1[1]), .out(far_5_5971_2[1]));
    assign layer_5[871] = ~far_5_5971_2[0]; 
    wire [1:0] far_5_5972_0;    relay_conn far_5_5972_0_a(.in(layer_4[711]), .out(far_5_5972_0[0]));    relay_conn far_5_5972_0_b(.in(layer_4[630]), .out(far_5_5972_0[1]));
    wire [1:0] far_5_5972_1;    relay_conn far_5_5972_1_a(.in(far_5_5972_0[0]), .out(far_5_5972_1[0]));    relay_conn far_5_5972_1_b(.in(far_5_5972_0[1]), .out(far_5_5972_1[1]));
    assign layer_5[872] = ~far_5_5972_1[1]; 
    wire [1:0] far_5_5973_0;    relay_conn far_5_5973_0_a(.in(layer_4[223]), .out(far_5_5973_0[0]));    relay_conn far_5_5973_0_b(.in(layer_4[291]), .out(far_5_5973_0[1]));
    wire [1:0] far_5_5973_1;    relay_conn far_5_5973_1_a(.in(far_5_5973_0[0]), .out(far_5_5973_1[0]));    relay_conn far_5_5973_1_b(.in(far_5_5973_0[1]), .out(far_5_5973_1[1]));
    assign layer_5[873] = ~(far_5_5973_1[0] | far_5_5973_1[1]); 
    wire [1:0] far_5_5974_0;    relay_conn far_5_5974_0_a(.in(layer_4[135]), .out(far_5_5974_0[0]));    relay_conn far_5_5974_0_b(.in(layer_4[90]), .out(far_5_5974_0[1]));
    assign layer_5[874] = far_5_5974_0[1]; 
    wire [1:0] far_5_5975_0;    relay_conn far_5_5975_0_a(.in(layer_4[322]), .out(far_5_5975_0[0]));    relay_conn far_5_5975_0_b(.in(layer_4[420]), .out(far_5_5975_0[1]));
    wire [1:0] far_5_5975_1;    relay_conn far_5_5975_1_a(.in(far_5_5975_0[0]), .out(far_5_5975_1[0]));    relay_conn far_5_5975_1_b(.in(far_5_5975_0[1]), .out(far_5_5975_1[1]));
    wire [1:0] far_5_5975_2;    relay_conn far_5_5975_2_a(.in(far_5_5975_1[0]), .out(far_5_5975_2[0]));    relay_conn far_5_5975_2_b(.in(far_5_5975_1[1]), .out(far_5_5975_2[1]));
    assign layer_5[875] = ~far_5_5975_2[0] | (far_5_5975_2[0] & far_5_5975_2[1]); 
    wire [1:0] far_5_5976_0;    relay_conn far_5_5976_0_a(.in(layer_4[778]), .out(far_5_5976_0[0]));    relay_conn far_5_5976_0_b(.in(layer_4[680]), .out(far_5_5976_0[1]));
    wire [1:0] far_5_5976_1;    relay_conn far_5_5976_1_a(.in(far_5_5976_0[0]), .out(far_5_5976_1[0]));    relay_conn far_5_5976_1_b(.in(far_5_5976_0[1]), .out(far_5_5976_1[1]));
    wire [1:0] far_5_5976_2;    relay_conn far_5_5976_2_a(.in(far_5_5976_1[0]), .out(far_5_5976_2[0]));    relay_conn far_5_5976_2_b(.in(far_5_5976_1[1]), .out(far_5_5976_2[1]));
    assign layer_5[876] = far_5_5976_2[0] & far_5_5976_2[1]; 
    wire [1:0] far_5_5977_0;    relay_conn far_5_5977_0_a(.in(layer_4[97]), .out(far_5_5977_0[0]));    relay_conn far_5_5977_0_b(.in(layer_4[156]), .out(far_5_5977_0[1]));
    assign layer_5[877] = far_5_5977_0[0]; 
    wire [1:0] far_5_5978_0;    relay_conn far_5_5978_0_a(.in(layer_4[360]), .out(far_5_5978_0[0]));    relay_conn far_5_5978_0_b(.in(layer_4[442]), .out(far_5_5978_0[1]));
    wire [1:0] far_5_5978_1;    relay_conn far_5_5978_1_a(.in(far_5_5978_0[0]), .out(far_5_5978_1[0]));    relay_conn far_5_5978_1_b(.in(far_5_5978_0[1]), .out(far_5_5978_1[1]));
    assign layer_5[878] = ~(far_5_5978_1[0] | far_5_5978_1[1]); 
    assign layer_5[879] = layer_4[665]; 
    assign layer_5[880] = ~(layer_4[190] ^ layer_4[163]); 
    assign layer_5[881] = ~(layer_4[869] | layer_4[852]); 
    wire [1:0] far_5_5982_0;    relay_conn far_5_5982_0_a(.in(layer_4[181]), .out(far_5_5982_0[0]));    relay_conn far_5_5982_0_b(.in(layer_4[279]), .out(far_5_5982_0[1]));
    wire [1:0] far_5_5982_1;    relay_conn far_5_5982_1_a(.in(far_5_5982_0[0]), .out(far_5_5982_1[0]));    relay_conn far_5_5982_1_b(.in(far_5_5982_0[1]), .out(far_5_5982_1[1]));
    wire [1:0] far_5_5982_2;    relay_conn far_5_5982_2_a(.in(far_5_5982_1[0]), .out(far_5_5982_2[0]));    relay_conn far_5_5982_2_b(.in(far_5_5982_1[1]), .out(far_5_5982_2[1]));
    assign layer_5[882] = ~far_5_5982_2[0] | (far_5_5982_2[0] & far_5_5982_2[1]); 
    wire [1:0] far_5_5983_0;    relay_conn far_5_5983_0_a(.in(layer_4[516]), .out(far_5_5983_0[0]));    relay_conn far_5_5983_0_b(.in(layer_4[389]), .out(far_5_5983_0[1]));
    wire [1:0] far_5_5983_1;    relay_conn far_5_5983_1_a(.in(far_5_5983_0[0]), .out(far_5_5983_1[0]));    relay_conn far_5_5983_1_b(.in(far_5_5983_0[1]), .out(far_5_5983_1[1]));
    wire [1:0] far_5_5983_2;    relay_conn far_5_5983_2_a(.in(far_5_5983_1[0]), .out(far_5_5983_2[0]));    relay_conn far_5_5983_2_b(.in(far_5_5983_1[1]), .out(far_5_5983_2[1]));
    assign layer_5[883] = far_5_5983_2[0]; 
    wire [1:0] far_5_5984_0;    relay_conn far_5_5984_0_a(.in(layer_4[84]), .out(far_5_5984_0[0]));    relay_conn far_5_5984_0_b(.in(layer_4[12]), .out(far_5_5984_0[1]));
    wire [1:0] far_5_5984_1;    relay_conn far_5_5984_1_a(.in(far_5_5984_0[0]), .out(far_5_5984_1[0]));    relay_conn far_5_5984_1_b(.in(far_5_5984_0[1]), .out(far_5_5984_1[1]));
    assign layer_5[884] = far_5_5984_1[0]; 
    assign layer_5[885] = ~(layer_4[875] ^ layer_4[879]); 
    wire [1:0] far_5_5986_0;    relay_conn far_5_5986_0_a(.in(layer_4[249]), .out(far_5_5986_0[0]));    relay_conn far_5_5986_0_b(.in(layer_4[122]), .out(far_5_5986_0[1]));
    wire [1:0] far_5_5986_1;    relay_conn far_5_5986_1_a(.in(far_5_5986_0[0]), .out(far_5_5986_1[0]));    relay_conn far_5_5986_1_b(.in(far_5_5986_0[1]), .out(far_5_5986_1[1]));
    wire [1:0] far_5_5986_2;    relay_conn far_5_5986_2_a(.in(far_5_5986_1[0]), .out(far_5_5986_2[0]));    relay_conn far_5_5986_2_b(.in(far_5_5986_1[1]), .out(far_5_5986_2[1]));
    assign layer_5[886] = far_5_5986_2[1]; 
    wire [1:0] far_5_5987_0;    relay_conn far_5_5987_0_a(.in(layer_4[136]), .out(far_5_5987_0[0]));    relay_conn far_5_5987_0_b(.in(layer_4[185]), .out(far_5_5987_0[1]));
    assign layer_5[887] = far_5_5987_0[1] & ~far_5_5987_0[0]; 
    wire [1:0] far_5_5988_0;    relay_conn far_5_5988_0_a(.in(layer_4[766]), .out(far_5_5988_0[0]));    relay_conn far_5_5988_0_b(.in(layer_4[657]), .out(far_5_5988_0[1]));
    wire [1:0] far_5_5988_1;    relay_conn far_5_5988_1_a(.in(far_5_5988_0[0]), .out(far_5_5988_1[0]));    relay_conn far_5_5988_1_b(.in(far_5_5988_0[1]), .out(far_5_5988_1[1]));
    wire [1:0] far_5_5988_2;    relay_conn far_5_5988_2_a(.in(far_5_5988_1[0]), .out(far_5_5988_2[0]));    relay_conn far_5_5988_2_b(.in(far_5_5988_1[1]), .out(far_5_5988_2[1]));
    assign layer_5[888] = far_5_5988_2[0]; 
    wire [1:0] far_5_5989_0;    relay_conn far_5_5989_0_a(.in(layer_4[593]), .out(far_5_5989_0[0]));    relay_conn far_5_5989_0_b(.in(layer_4[658]), .out(far_5_5989_0[1]));
    wire [1:0] far_5_5989_1;    relay_conn far_5_5989_1_a(.in(far_5_5989_0[0]), .out(far_5_5989_1[0]));    relay_conn far_5_5989_1_b(.in(far_5_5989_0[1]), .out(far_5_5989_1[1]));
    assign layer_5[889] = ~far_5_5989_1[0] | (far_5_5989_1[0] & far_5_5989_1[1]); 
    assign layer_5[890] = layer_4[381] & ~layer_4[361]; 
    assign layer_5[891] = layer_4[833]; 
    wire [1:0] far_5_5992_0;    relay_conn far_5_5992_0_a(.in(layer_4[899]), .out(far_5_5992_0[0]));    relay_conn far_5_5992_0_b(.in(layer_4[980]), .out(far_5_5992_0[1]));
    wire [1:0] far_5_5992_1;    relay_conn far_5_5992_1_a(.in(far_5_5992_0[0]), .out(far_5_5992_1[0]));    relay_conn far_5_5992_1_b(.in(far_5_5992_0[1]), .out(far_5_5992_1[1]));
    assign layer_5[892] = far_5_5992_1[1] & ~far_5_5992_1[0]; 
    wire [1:0] far_5_5993_0;    relay_conn far_5_5993_0_a(.in(layer_4[520]), .out(far_5_5993_0[0]));    relay_conn far_5_5993_0_b(.in(layer_4[468]), .out(far_5_5993_0[1]));
    assign layer_5[893] = far_5_5993_0[1]; 
    wire [1:0] far_5_5994_0;    relay_conn far_5_5994_0_a(.in(layer_4[1015]), .out(far_5_5994_0[0]));    relay_conn far_5_5994_0_b(.in(layer_4[910]), .out(far_5_5994_0[1]));
    wire [1:0] far_5_5994_1;    relay_conn far_5_5994_1_a(.in(far_5_5994_0[0]), .out(far_5_5994_1[0]));    relay_conn far_5_5994_1_b(.in(far_5_5994_0[1]), .out(far_5_5994_1[1]));
    wire [1:0] far_5_5994_2;    relay_conn far_5_5994_2_a(.in(far_5_5994_1[0]), .out(far_5_5994_2[0]));    relay_conn far_5_5994_2_b(.in(far_5_5994_1[1]), .out(far_5_5994_2[1]));
    assign layer_5[894] = ~(far_5_5994_2[0] ^ far_5_5994_2[1]); 
    wire [1:0] far_5_5995_0;    relay_conn far_5_5995_0_a(.in(layer_4[806]), .out(far_5_5995_0[0]));    relay_conn far_5_5995_0_b(.in(layer_4[921]), .out(far_5_5995_0[1]));
    wire [1:0] far_5_5995_1;    relay_conn far_5_5995_1_a(.in(far_5_5995_0[0]), .out(far_5_5995_1[0]));    relay_conn far_5_5995_1_b(.in(far_5_5995_0[1]), .out(far_5_5995_1[1]));
    wire [1:0] far_5_5995_2;    relay_conn far_5_5995_2_a(.in(far_5_5995_1[0]), .out(far_5_5995_2[0]));    relay_conn far_5_5995_2_b(.in(far_5_5995_1[1]), .out(far_5_5995_2[1]));
    assign layer_5[895] = far_5_5995_2[0]; 
    wire [1:0] far_5_5996_0;    relay_conn far_5_5996_0_a(.in(layer_4[538]), .out(far_5_5996_0[0]));    relay_conn far_5_5996_0_b(.in(layer_4[443]), .out(far_5_5996_0[1]));
    wire [1:0] far_5_5996_1;    relay_conn far_5_5996_1_a(.in(far_5_5996_0[0]), .out(far_5_5996_1[0]));    relay_conn far_5_5996_1_b(.in(far_5_5996_0[1]), .out(far_5_5996_1[1]));
    assign layer_5[896] = far_5_5996_1[1] & ~far_5_5996_1[0]; 
    assign layer_5[897] = layer_4[369]; 
    wire [1:0] far_5_5998_0;    relay_conn far_5_5998_0_a(.in(layer_4[665]), .out(far_5_5998_0[0]));    relay_conn far_5_5998_0_b(.in(layer_4[538]), .out(far_5_5998_0[1]));
    wire [1:0] far_5_5998_1;    relay_conn far_5_5998_1_a(.in(far_5_5998_0[0]), .out(far_5_5998_1[0]));    relay_conn far_5_5998_1_b(.in(far_5_5998_0[1]), .out(far_5_5998_1[1]));
    wire [1:0] far_5_5998_2;    relay_conn far_5_5998_2_a(.in(far_5_5998_1[0]), .out(far_5_5998_2[0]));    relay_conn far_5_5998_2_b(.in(far_5_5998_1[1]), .out(far_5_5998_2[1]));
    assign layer_5[898] = far_5_5998_2[0]; 
    assign layer_5[899] = layer_4[337] | layer_4[318]; 
    wire [1:0] far_5_6000_0;    relay_conn far_5_6000_0_a(.in(layer_4[300]), .out(far_5_6000_0[0]));    relay_conn far_5_6000_0_b(.in(layer_4[217]), .out(far_5_6000_0[1]));
    wire [1:0] far_5_6000_1;    relay_conn far_5_6000_1_a(.in(far_5_6000_0[0]), .out(far_5_6000_1[0]));    relay_conn far_5_6000_1_b(.in(far_5_6000_0[1]), .out(far_5_6000_1[1]));
    assign layer_5[900] = far_5_6000_1[0] & ~far_5_6000_1[1]; 
    wire [1:0] far_5_6001_0;    relay_conn far_5_6001_0_a(.in(layer_4[569]), .out(far_5_6001_0[0]));    relay_conn far_5_6001_0_b(.in(layer_4[654]), .out(far_5_6001_0[1]));
    wire [1:0] far_5_6001_1;    relay_conn far_5_6001_1_a(.in(far_5_6001_0[0]), .out(far_5_6001_1[0]));    relay_conn far_5_6001_1_b(.in(far_5_6001_0[1]), .out(far_5_6001_1[1]));
    assign layer_5[901] = ~far_5_6001_1[1]; 
    wire [1:0] far_5_6002_0;    relay_conn far_5_6002_0_a(.in(layer_4[833]), .out(far_5_6002_0[0]));    relay_conn far_5_6002_0_b(.in(layer_4[711]), .out(far_5_6002_0[1]));
    wire [1:0] far_5_6002_1;    relay_conn far_5_6002_1_a(.in(far_5_6002_0[0]), .out(far_5_6002_1[0]));    relay_conn far_5_6002_1_b(.in(far_5_6002_0[1]), .out(far_5_6002_1[1]));
    wire [1:0] far_5_6002_2;    relay_conn far_5_6002_2_a(.in(far_5_6002_1[0]), .out(far_5_6002_2[0]));    relay_conn far_5_6002_2_b(.in(far_5_6002_1[1]), .out(far_5_6002_2[1]));
    assign layer_5[902] = far_5_6002_2[0] | far_5_6002_2[1]; 
    wire [1:0] far_5_6003_0;    relay_conn far_5_6003_0_a(.in(layer_4[713]), .out(far_5_6003_0[0]));    relay_conn far_5_6003_0_b(.in(layer_4[597]), .out(far_5_6003_0[1]));
    wire [1:0] far_5_6003_1;    relay_conn far_5_6003_1_a(.in(far_5_6003_0[0]), .out(far_5_6003_1[0]));    relay_conn far_5_6003_1_b(.in(far_5_6003_0[1]), .out(far_5_6003_1[1]));
    wire [1:0] far_5_6003_2;    relay_conn far_5_6003_2_a(.in(far_5_6003_1[0]), .out(far_5_6003_2[0]));    relay_conn far_5_6003_2_b(.in(far_5_6003_1[1]), .out(far_5_6003_2[1]));
    assign layer_5[903] = ~far_5_6003_2[1] | (far_5_6003_2[0] & far_5_6003_2[1]); 
    wire [1:0] far_5_6004_0;    relay_conn far_5_6004_0_a(.in(layer_4[337]), .out(far_5_6004_0[0]));    relay_conn far_5_6004_0_b(.in(layer_4[381]), .out(far_5_6004_0[1]));
    assign layer_5[904] = far_5_6004_0[0] ^ far_5_6004_0[1]; 
    assign layer_5[905] = ~layer_4[857]; 
    assign layer_5[906] = layer_4[685]; 
    wire [1:0] far_5_6007_0;    relay_conn far_5_6007_0_a(.in(layer_4[911]), .out(far_5_6007_0[0]));    relay_conn far_5_6007_0_b(.in(layer_4[797]), .out(far_5_6007_0[1]));
    wire [1:0] far_5_6007_1;    relay_conn far_5_6007_1_a(.in(far_5_6007_0[0]), .out(far_5_6007_1[0]));    relay_conn far_5_6007_1_b(.in(far_5_6007_0[1]), .out(far_5_6007_1[1]));
    wire [1:0] far_5_6007_2;    relay_conn far_5_6007_2_a(.in(far_5_6007_1[0]), .out(far_5_6007_2[0]));    relay_conn far_5_6007_2_b(.in(far_5_6007_1[1]), .out(far_5_6007_2[1]));
    assign layer_5[907] = ~far_5_6007_2[0] | (far_5_6007_2[0] & far_5_6007_2[1]); 
    wire [1:0] far_5_6008_0;    relay_conn far_5_6008_0_a(.in(layer_4[333]), .out(far_5_6008_0[0]));    relay_conn far_5_6008_0_b(.in(layer_4[394]), .out(far_5_6008_0[1]));
    assign layer_5[908] = ~(far_5_6008_0[0] & far_5_6008_0[1]); 
    wire [1:0] far_5_6009_0;    relay_conn far_5_6009_0_a(.in(layer_4[596]), .out(far_5_6009_0[0]));    relay_conn far_5_6009_0_b(.in(layer_4[469]), .out(far_5_6009_0[1]));
    wire [1:0] far_5_6009_1;    relay_conn far_5_6009_1_a(.in(far_5_6009_0[0]), .out(far_5_6009_1[0]));    relay_conn far_5_6009_1_b(.in(far_5_6009_0[1]), .out(far_5_6009_1[1]));
    wire [1:0] far_5_6009_2;    relay_conn far_5_6009_2_a(.in(far_5_6009_1[0]), .out(far_5_6009_2[0]));    relay_conn far_5_6009_2_b(.in(far_5_6009_1[1]), .out(far_5_6009_2[1]));
    assign layer_5[909] = ~far_5_6009_2[1] | (far_5_6009_2[0] & far_5_6009_2[1]); 
    wire [1:0] far_5_6010_0;    relay_conn far_5_6010_0_a(.in(layer_4[597]), .out(far_5_6010_0[0]));    relay_conn far_5_6010_0_b(.in(layer_4[673]), .out(far_5_6010_0[1]));
    wire [1:0] far_5_6010_1;    relay_conn far_5_6010_1_a(.in(far_5_6010_0[0]), .out(far_5_6010_1[0]));    relay_conn far_5_6010_1_b(.in(far_5_6010_0[1]), .out(far_5_6010_1[1]));
    assign layer_5[910] = far_5_6010_1[0] & far_5_6010_1[1]; 
    wire [1:0] far_5_6011_0;    relay_conn far_5_6011_0_a(.in(layer_4[304]), .out(far_5_6011_0[0]));    relay_conn far_5_6011_0_b(.in(layer_4[360]), .out(far_5_6011_0[1]));
    assign layer_5[911] = far_5_6011_0[0] | far_5_6011_0[1]; 
    assign layer_5[912] = ~layer_4[402] | (layer_4[402] & layer_4[398]); 
    wire [1:0] far_5_6013_0;    relay_conn far_5_6013_0_a(.in(layer_4[785]), .out(far_5_6013_0[0]));    relay_conn far_5_6013_0_b(.in(layer_4[709]), .out(far_5_6013_0[1]));
    wire [1:0] far_5_6013_1;    relay_conn far_5_6013_1_a(.in(far_5_6013_0[0]), .out(far_5_6013_1[0]));    relay_conn far_5_6013_1_b(.in(far_5_6013_0[1]), .out(far_5_6013_1[1]));
    assign layer_5[913] = ~far_5_6013_1[0]; 
    wire [1:0] far_5_6014_0;    relay_conn far_5_6014_0_a(.in(layer_4[248]), .out(far_5_6014_0[0]));    relay_conn far_5_6014_0_b(.in(layer_4[142]), .out(far_5_6014_0[1]));
    wire [1:0] far_5_6014_1;    relay_conn far_5_6014_1_a(.in(far_5_6014_0[0]), .out(far_5_6014_1[0]));    relay_conn far_5_6014_1_b(.in(far_5_6014_0[1]), .out(far_5_6014_1[1]));
    wire [1:0] far_5_6014_2;    relay_conn far_5_6014_2_a(.in(far_5_6014_1[0]), .out(far_5_6014_2[0]));    relay_conn far_5_6014_2_b(.in(far_5_6014_1[1]), .out(far_5_6014_2[1]));
    assign layer_5[914] = ~far_5_6014_2[0]; 
    wire [1:0] far_5_6015_0;    relay_conn far_5_6015_0_a(.in(layer_4[357]), .out(far_5_6015_0[0]));    relay_conn far_5_6015_0_b(.in(layer_4[443]), .out(far_5_6015_0[1]));
    wire [1:0] far_5_6015_1;    relay_conn far_5_6015_1_a(.in(far_5_6015_0[0]), .out(far_5_6015_1[0]));    relay_conn far_5_6015_1_b(.in(far_5_6015_0[1]), .out(far_5_6015_1[1]));
    assign layer_5[915] = far_5_6015_1[0]; 
    assign layer_5[916] = layer_4[787] & ~layer_4[789]; 
    wire [1:0] far_5_6017_0;    relay_conn far_5_6017_0_a(.in(layer_4[938]), .out(far_5_6017_0[0]));    relay_conn far_5_6017_0_b(.in(layer_4[850]), .out(far_5_6017_0[1]));
    wire [1:0] far_5_6017_1;    relay_conn far_5_6017_1_a(.in(far_5_6017_0[0]), .out(far_5_6017_1[0]));    relay_conn far_5_6017_1_b(.in(far_5_6017_0[1]), .out(far_5_6017_1[1]));
    assign layer_5[917] = far_5_6017_1[1]; 
    assign layer_5[918] = ~layer_4[282] | (layer_4[305] & layer_4[282]); 
    wire [1:0] far_5_6019_0;    relay_conn far_5_6019_0_a(.in(layer_4[499]), .out(far_5_6019_0[0]));    relay_conn far_5_6019_0_b(.in(layer_4[583]), .out(far_5_6019_0[1]));
    wire [1:0] far_5_6019_1;    relay_conn far_5_6019_1_a(.in(far_5_6019_0[0]), .out(far_5_6019_1[0]));    relay_conn far_5_6019_1_b(.in(far_5_6019_0[1]), .out(far_5_6019_1[1]));
    assign layer_5[919] = far_5_6019_1[1]; 
    wire [1:0] far_5_6020_0;    relay_conn far_5_6020_0_a(.in(layer_4[660]), .out(far_5_6020_0[0]));    relay_conn far_5_6020_0_b(.in(layer_4[718]), .out(far_5_6020_0[1]));
    assign layer_5[920] = ~(far_5_6020_0[0] | far_5_6020_0[1]); 
    assign layer_5[921] = ~layer_4[631] | (layer_4[631] & layer_4[636]); 
    wire [1:0] far_5_6022_0;    relay_conn far_5_6022_0_a(.in(layer_4[200]), .out(far_5_6022_0[0]));    relay_conn far_5_6022_0_b(.in(layer_4[300]), .out(far_5_6022_0[1]));
    wire [1:0] far_5_6022_1;    relay_conn far_5_6022_1_a(.in(far_5_6022_0[0]), .out(far_5_6022_1[0]));    relay_conn far_5_6022_1_b(.in(far_5_6022_0[1]), .out(far_5_6022_1[1]));
    wire [1:0] far_5_6022_2;    relay_conn far_5_6022_2_a(.in(far_5_6022_1[0]), .out(far_5_6022_2[0]));    relay_conn far_5_6022_2_b(.in(far_5_6022_1[1]), .out(far_5_6022_2[1]));
    assign layer_5[922] = ~far_5_6022_2[0]; 
    wire [1:0] far_5_6023_0;    relay_conn far_5_6023_0_a(.in(layer_4[507]), .out(far_5_6023_0[0]));    relay_conn far_5_6023_0_b(.in(layer_4[428]), .out(far_5_6023_0[1]));
    wire [1:0] far_5_6023_1;    relay_conn far_5_6023_1_a(.in(far_5_6023_0[0]), .out(far_5_6023_1[0]));    relay_conn far_5_6023_1_b(.in(far_5_6023_0[1]), .out(far_5_6023_1[1]));
    assign layer_5[923] = ~far_5_6023_1[0] | (far_5_6023_1[0] & far_5_6023_1[1]); 
    wire [1:0] far_5_6024_0;    relay_conn far_5_6024_0_a(.in(layer_4[703]), .out(far_5_6024_0[0]));    relay_conn far_5_6024_0_b(.in(layer_4[745]), .out(far_5_6024_0[1]));
    assign layer_5[924] = ~far_5_6024_0[0] | (far_5_6024_0[0] & far_5_6024_0[1]); 
    assign layer_5[925] = ~layer_4[567]; 
    wire [1:0] far_5_6026_0;    relay_conn far_5_6026_0_a(.in(layer_4[970]), .out(far_5_6026_0[0]));    relay_conn far_5_6026_0_b(.in(layer_4[872]), .out(far_5_6026_0[1]));
    wire [1:0] far_5_6026_1;    relay_conn far_5_6026_1_a(.in(far_5_6026_0[0]), .out(far_5_6026_1[0]));    relay_conn far_5_6026_1_b(.in(far_5_6026_0[1]), .out(far_5_6026_1[1]));
    wire [1:0] far_5_6026_2;    relay_conn far_5_6026_2_a(.in(far_5_6026_1[0]), .out(far_5_6026_2[0]));    relay_conn far_5_6026_2_b(.in(far_5_6026_1[1]), .out(far_5_6026_2[1]));
    assign layer_5[926] = ~far_5_6026_2[1]; 
    wire [1:0] far_5_6027_0;    relay_conn far_5_6027_0_a(.in(layer_4[325]), .out(far_5_6027_0[0]));    relay_conn far_5_6027_0_b(.in(layer_4[242]), .out(far_5_6027_0[1]));
    wire [1:0] far_5_6027_1;    relay_conn far_5_6027_1_a(.in(far_5_6027_0[0]), .out(far_5_6027_1[0]));    relay_conn far_5_6027_1_b(.in(far_5_6027_0[1]), .out(far_5_6027_1[1]));
    assign layer_5[927] = far_5_6027_1[0]; 
    wire [1:0] far_5_6028_0;    relay_conn far_5_6028_0_a(.in(layer_4[283]), .out(far_5_6028_0[0]));    relay_conn far_5_6028_0_b(.in(layer_4[387]), .out(far_5_6028_0[1]));
    wire [1:0] far_5_6028_1;    relay_conn far_5_6028_1_a(.in(far_5_6028_0[0]), .out(far_5_6028_1[0]));    relay_conn far_5_6028_1_b(.in(far_5_6028_0[1]), .out(far_5_6028_1[1]));
    wire [1:0] far_5_6028_2;    relay_conn far_5_6028_2_a(.in(far_5_6028_1[0]), .out(far_5_6028_2[0]));    relay_conn far_5_6028_2_b(.in(far_5_6028_1[1]), .out(far_5_6028_2[1]));
    assign layer_5[928] = far_5_6028_2[0] ^ far_5_6028_2[1]; 
    wire [1:0] far_5_6029_0;    relay_conn far_5_6029_0_a(.in(layer_4[997]), .out(far_5_6029_0[0]));    relay_conn far_5_6029_0_b(.in(layer_4[947]), .out(far_5_6029_0[1]));
    assign layer_5[929] = far_5_6029_0[0] ^ far_5_6029_0[1]; 
    wire [1:0] far_5_6030_0;    relay_conn far_5_6030_0_a(.in(layer_4[370]), .out(far_5_6030_0[0]));    relay_conn far_5_6030_0_b(.in(layer_4[423]), .out(far_5_6030_0[1]));
    assign layer_5[930] = ~(far_5_6030_0[0] | far_5_6030_0[1]); 
    assign layer_5[931] = layer_4[888] & ~layer_4[893]; 
    wire [1:0] far_5_6032_0;    relay_conn far_5_6032_0_a(.in(layer_4[867]), .out(far_5_6032_0[0]));    relay_conn far_5_6032_0_b(.in(layer_4[933]), .out(far_5_6032_0[1]));
    wire [1:0] far_5_6032_1;    relay_conn far_5_6032_1_a(.in(far_5_6032_0[0]), .out(far_5_6032_1[0]));    relay_conn far_5_6032_1_b(.in(far_5_6032_0[1]), .out(far_5_6032_1[1]));
    assign layer_5[932] = far_5_6032_1[0] & far_5_6032_1[1]; 
    wire [1:0] far_5_6033_0;    relay_conn far_5_6033_0_a(.in(layer_4[467]), .out(far_5_6033_0[0]));    relay_conn far_5_6033_0_b(.in(layer_4[415]), .out(far_5_6033_0[1]));
    assign layer_5[933] = far_5_6033_0[1]; 
    wire [1:0] far_5_6034_0;    relay_conn far_5_6034_0_a(.in(layer_4[443]), .out(far_5_6034_0[0]));    relay_conn far_5_6034_0_b(.in(layer_4[559]), .out(far_5_6034_0[1]));
    wire [1:0] far_5_6034_1;    relay_conn far_5_6034_1_a(.in(far_5_6034_0[0]), .out(far_5_6034_1[0]));    relay_conn far_5_6034_1_b(.in(far_5_6034_0[1]), .out(far_5_6034_1[1]));
    wire [1:0] far_5_6034_2;    relay_conn far_5_6034_2_a(.in(far_5_6034_1[0]), .out(far_5_6034_2[0]));    relay_conn far_5_6034_2_b(.in(far_5_6034_1[1]), .out(far_5_6034_2[1]));
    assign layer_5[934] = far_5_6034_2[1]; 
    wire [1:0] far_5_6035_0;    relay_conn far_5_6035_0_a(.in(layer_4[644]), .out(far_5_6035_0[0]));    relay_conn far_5_6035_0_b(.in(layer_4[683]), .out(far_5_6035_0[1]));
    assign layer_5[935] = far_5_6035_0[1] & ~far_5_6035_0[0]; 
    wire [1:0] far_5_6036_0;    relay_conn far_5_6036_0_a(.in(layer_4[167]), .out(far_5_6036_0[0]));    relay_conn far_5_6036_0_b(.in(layer_4[217]), .out(far_5_6036_0[1]));
    assign layer_5[936] = ~far_5_6036_0[0] | (far_5_6036_0[0] & far_5_6036_0[1]); 
    wire [1:0] far_5_6037_0;    relay_conn far_5_6037_0_a(.in(layer_4[520]), .out(far_5_6037_0[0]));    relay_conn far_5_6037_0_b(.in(layer_4[424]), .out(far_5_6037_0[1]));
    wire [1:0] far_5_6037_1;    relay_conn far_5_6037_1_a(.in(far_5_6037_0[0]), .out(far_5_6037_1[0]));    relay_conn far_5_6037_1_b(.in(far_5_6037_0[1]), .out(far_5_6037_1[1]));
    wire [1:0] far_5_6037_2;    relay_conn far_5_6037_2_a(.in(far_5_6037_1[0]), .out(far_5_6037_2[0]));    relay_conn far_5_6037_2_b(.in(far_5_6037_1[1]), .out(far_5_6037_2[1]));
    assign layer_5[937] = far_5_6037_2[0] ^ far_5_6037_2[1]; 
    wire [1:0] far_5_6038_0;    relay_conn far_5_6038_0_a(.in(layer_4[896]), .out(far_5_6038_0[0]));    relay_conn far_5_6038_0_b(.in(layer_4[999]), .out(far_5_6038_0[1]));
    wire [1:0] far_5_6038_1;    relay_conn far_5_6038_1_a(.in(far_5_6038_0[0]), .out(far_5_6038_1[0]));    relay_conn far_5_6038_1_b(.in(far_5_6038_0[1]), .out(far_5_6038_1[1]));
    wire [1:0] far_5_6038_2;    relay_conn far_5_6038_2_a(.in(far_5_6038_1[0]), .out(far_5_6038_2[0]));    relay_conn far_5_6038_2_b(.in(far_5_6038_1[1]), .out(far_5_6038_2[1]));
    assign layer_5[938] = far_5_6038_2[0] & ~far_5_6038_2[1]; 
    assign layer_5[939] = layer_4[622] & layer_4[644]; 
    wire [1:0] far_5_6040_0;    relay_conn far_5_6040_0_a(.in(layer_4[294]), .out(far_5_6040_0[0]));    relay_conn far_5_6040_0_b(.in(layer_4[361]), .out(far_5_6040_0[1]));
    wire [1:0] far_5_6040_1;    relay_conn far_5_6040_1_a(.in(far_5_6040_0[0]), .out(far_5_6040_1[0]));    relay_conn far_5_6040_1_b(.in(far_5_6040_0[1]), .out(far_5_6040_1[1]));
    assign layer_5[940] = far_5_6040_1[0] | far_5_6040_1[1]; 
    wire [1:0] far_5_6041_0;    relay_conn far_5_6041_0_a(.in(layer_4[22]), .out(far_5_6041_0[0]));    relay_conn far_5_6041_0_b(.in(layer_4[63]), .out(far_5_6041_0[1]));
    assign layer_5[941] = ~(far_5_6041_0[0] ^ far_5_6041_0[1]); 
    assign layer_5[942] = layer_4[790] | layer_4[800]; 
    assign layer_5[943] = layer_4[164] & ~layer_4[181]; 
    wire [1:0] far_5_6044_0;    relay_conn far_5_6044_0_a(.in(layer_4[921]), .out(far_5_6044_0[0]));    relay_conn far_5_6044_0_b(.in(layer_4[986]), .out(far_5_6044_0[1]));
    wire [1:0] far_5_6044_1;    relay_conn far_5_6044_1_a(.in(far_5_6044_0[0]), .out(far_5_6044_1[0]));    relay_conn far_5_6044_1_b(.in(far_5_6044_0[1]), .out(far_5_6044_1[1]));
    assign layer_5[944] = ~far_5_6044_1[1]; 
    wire [1:0] far_5_6045_0;    relay_conn far_5_6045_0_a(.in(layer_4[525]), .out(far_5_6045_0[0]));    relay_conn far_5_6045_0_b(.in(layer_4[597]), .out(far_5_6045_0[1]));
    wire [1:0] far_5_6045_1;    relay_conn far_5_6045_1_a(.in(far_5_6045_0[0]), .out(far_5_6045_1[0]));    relay_conn far_5_6045_1_b(.in(far_5_6045_0[1]), .out(far_5_6045_1[1]));
    assign layer_5[945] = ~(far_5_6045_1[0] & far_5_6045_1[1]); 
    wire [1:0] far_5_6046_0;    relay_conn far_5_6046_0_a(.in(layer_4[999]), .out(far_5_6046_0[0]));    relay_conn far_5_6046_0_b(.in(layer_4[910]), .out(far_5_6046_0[1]));
    wire [1:0] far_5_6046_1;    relay_conn far_5_6046_1_a(.in(far_5_6046_0[0]), .out(far_5_6046_1[0]));    relay_conn far_5_6046_1_b(.in(far_5_6046_0[1]), .out(far_5_6046_1[1]));
    assign layer_5[946] = far_5_6046_1[0]; 
    wire [1:0] far_5_6047_0;    relay_conn far_5_6047_0_a(.in(layer_4[773]), .out(far_5_6047_0[0]));    relay_conn far_5_6047_0_b(.in(layer_4[658]), .out(far_5_6047_0[1]));
    wire [1:0] far_5_6047_1;    relay_conn far_5_6047_1_a(.in(far_5_6047_0[0]), .out(far_5_6047_1[0]));    relay_conn far_5_6047_1_b(.in(far_5_6047_0[1]), .out(far_5_6047_1[1]));
    wire [1:0] far_5_6047_2;    relay_conn far_5_6047_2_a(.in(far_5_6047_1[0]), .out(far_5_6047_2[0]));    relay_conn far_5_6047_2_b(.in(far_5_6047_1[1]), .out(far_5_6047_2[1]));
    assign layer_5[947] = ~far_5_6047_2[0]; 
    wire [1:0] far_5_6048_0;    relay_conn far_5_6048_0_a(.in(layer_4[499]), .out(far_5_6048_0[0]));    relay_conn far_5_6048_0_b(.in(layer_4[602]), .out(far_5_6048_0[1]));
    wire [1:0] far_5_6048_1;    relay_conn far_5_6048_1_a(.in(far_5_6048_0[0]), .out(far_5_6048_1[0]));    relay_conn far_5_6048_1_b(.in(far_5_6048_0[1]), .out(far_5_6048_1[1]));
    wire [1:0] far_5_6048_2;    relay_conn far_5_6048_2_a(.in(far_5_6048_1[0]), .out(far_5_6048_2[0]));    relay_conn far_5_6048_2_b(.in(far_5_6048_1[1]), .out(far_5_6048_2[1]));
    assign layer_5[948] = ~far_5_6048_2[0]; 
    wire [1:0] far_5_6049_0;    relay_conn far_5_6049_0_a(.in(layer_4[650]), .out(far_5_6049_0[0]));    relay_conn far_5_6049_0_b(.in(layer_4[745]), .out(far_5_6049_0[1]));
    wire [1:0] far_5_6049_1;    relay_conn far_5_6049_1_a(.in(far_5_6049_0[0]), .out(far_5_6049_1[0]));    relay_conn far_5_6049_1_b(.in(far_5_6049_0[1]), .out(far_5_6049_1[1]));
    assign layer_5[949] = ~far_5_6049_1[0]; 
    wire [1:0] far_5_6050_0;    relay_conn far_5_6050_0_a(.in(layer_4[478]), .out(far_5_6050_0[0]));    relay_conn far_5_6050_0_b(.in(layer_4[386]), .out(far_5_6050_0[1]));
    wire [1:0] far_5_6050_1;    relay_conn far_5_6050_1_a(.in(far_5_6050_0[0]), .out(far_5_6050_1[0]));    relay_conn far_5_6050_1_b(.in(far_5_6050_0[1]), .out(far_5_6050_1[1]));
    assign layer_5[950] = far_5_6050_1[0]; 
    wire [1:0] far_5_6051_0;    relay_conn far_5_6051_0_a(.in(layer_4[197]), .out(far_5_6051_0[0]));    relay_conn far_5_6051_0_b(.in(layer_4[89]), .out(far_5_6051_0[1]));
    wire [1:0] far_5_6051_1;    relay_conn far_5_6051_1_a(.in(far_5_6051_0[0]), .out(far_5_6051_1[0]));    relay_conn far_5_6051_1_b(.in(far_5_6051_0[1]), .out(far_5_6051_1[1]));
    wire [1:0] far_5_6051_2;    relay_conn far_5_6051_2_a(.in(far_5_6051_1[0]), .out(far_5_6051_2[0]));    relay_conn far_5_6051_2_b(.in(far_5_6051_1[1]), .out(far_5_6051_2[1]));
    assign layer_5[951] = far_5_6051_2[1]; 
    wire [1:0] far_5_6052_0;    relay_conn far_5_6052_0_a(.in(layer_4[269]), .out(far_5_6052_0[0]));    relay_conn far_5_6052_0_b(.in(layer_4[215]), .out(far_5_6052_0[1]));
    assign layer_5[952] = far_5_6052_0[0] & ~far_5_6052_0[1]; 
    wire [1:0] far_5_6053_0;    relay_conn far_5_6053_0_a(.in(layer_4[386]), .out(far_5_6053_0[0]));    relay_conn far_5_6053_0_b(.in(layer_4[475]), .out(far_5_6053_0[1]));
    wire [1:0] far_5_6053_1;    relay_conn far_5_6053_1_a(.in(far_5_6053_0[0]), .out(far_5_6053_1[0]));    relay_conn far_5_6053_1_b(.in(far_5_6053_0[1]), .out(far_5_6053_1[1]));
    assign layer_5[953] = ~far_5_6053_1[0]; 
    wire [1:0] far_5_6054_0;    relay_conn far_5_6054_0_a(.in(layer_4[16]), .out(far_5_6054_0[0]));    relay_conn far_5_6054_0_b(.in(layer_4[59]), .out(far_5_6054_0[1]));
    assign layer_5[954] = ~far_5_6054_0[0]; 
    wire [1:0] far_5_6055_0;    relay_conn far_5_6055_0_a(.in(layer_4[718]), .out(far_5_6055_0[0]));    relay_conn far_5_6055_0_b(.in(layer_4[806]), .out(far_5_6055_0[1]));
    wire [1:0] far_5_6055_1;    relay_conn far_5_6055_1_a(.in(far_5_6055_0[0]), .out(far_5_6055_1[0]));    relay_conn far_5_6055_1_b(.in(far_5_6055_0[1]), .out(far_5_6055_1[1]));
    assign layer_5[955] = ~(far_5_6055_1[0] | far_5_6055_1[1]); 
    wire [1:0] far_5_6056_0;    relay_conn far_5_6056_0_a(.in(layer_4[123]), .out(far_5_6056_0[0]));    relay_conn far_5_6056_0_b(.in(layer_4[207]), .out(far_5_6056_0[1]));
    wire [1:0] far_5_6056_1;    relay_conn far_5_6056_1_a(.in(far_5_6056_0[0]), .out(far_5_6056_1[0]));    relay_conn far_5_6056_1_b(.in(far_5_6056_0[1]), .out(far_5_6056_1[1]));
    assign layer_5[956] = ~far_5_6056_1[0]; 
    wire [1:0] far_5_6057_0;    relay_conn far_5_6057_0_a(.in(layer_4[881]), .out(far_5_6057_0[0]));    relay_conn far_5_6057_0_b(.in(layer_4[830]), .out(far_5_6057_0[1]));
    assign layer_5[957] = ~(far_5_6057_0[0] | far_5_6057_0[1]); 
    wire [1:0] far_5_6058_0;    relay_conn far_5_6058_0_a(.in(layer_4[298]), .out(far_5_6058_0[0]));    relay_conn far_5_6058_0_b(.in(layer_4[176]), .out(far_5_6058_0[1]));
    wire [1:0] far_5_6058_1;    relay_conn far_5_6058_1_a(.in(far_5_6058_0[0]), .out(far_5_6058_1[0]));    relay_conn far_5_6058_1_b(.in(far_5_6058_0[1]), .out(far_5_6058_1[1]));
    wire [1:0] far_5_6058_2;    relay_conn far_5_6058_2_a(.in(far_5_6058_1[0]), .out(far_5_6058_2[0]));    relay_conn far_5_6058_2_b(.in(far_5_6058_1[1]), .out(far_5_6058_2[1]));
    assign layer_5[958] = far_5_6058_2[1] & ~far_5_6058_2[0]; 
    wire [1:0] far_5_6059_0;    relay_conn far_5_6059_0_a(.in(layer_4[711]), .out(far_5_6059_0[0]));    relay_conn far_5_6059_0_b(.in(layer_4[595]), .out(far_5_6059_0[1]));
    wire [1:0] far_5_6059_1;    relay_conn far_5_6059_1_a(.in(far_5_6059_0[0]), .out(far_5_6059_1[0]));    relay_conn far_5_6059_1_b(.in(far_5_6059_0[1]), .out(far_5_6059_1[1]));
    wire [1:0] far_5_6059_2;    relay_conn far_5_6059_2_a(.in(far_5_6059_1[0]), .out(far_5_6059_2[0]));    relay_conn far_5_6059_2_b(.in(far_5_6059_1[1]), .out(far_5_6059_2[1]));
    assign layer_5[959] = ~(far_5_6059_2[0] | far_5_6059_2[1]); 
    wire [1:0] far_5_6060_0;    relay_conn far_5_6060_0_a(.in(layer_4[970]), .out(far_5_6060_0[0]));    relay_conn far_5_6060_0_b(.in(layer_4[888]), .out(far_5_6060_0[1]));
    wire [1:0] far_5_6060_1;    relay_conn far_5_6060_1_a(.in(far_5_6060_0[0]), .out(far_5_6060_1[0]));    relay_conn far_5_6060_1_b(.in(far_5_6060_0[1]), .out(far_5_6060_1[1]));
    assign layer_5[960] = far_5_6060_1[0] | far_5_6060_1[1]; 
    wire [1:0] far_5_6061_0;    relay_conn far_5_6061_0_a(.in(layer_4[697]), .out(far_5_6061_0[0]));    relay_conn far_5_6061_0_b(.in(layer_4[589]), .out(far_5_6061_0[1]));
    wire [1:0] far_5_6061_1;    relay_conn far_5_6061_1_a(.in(far_5_6061_0[0]), .out(far_5_6061_1[0]));    relay_conn far_5_6061_1_b(.in(far_5_6061_0[1]), .out(far_5_6061_1[1]));
    wire [1:0] far_5_6061_2;    relay_conn far_5_6061_2_a(.in(far_5_6061_1[0]), .out(far_5_6061_2[0]));    relay_conn far_5_6061_2_b(.in(far_5_6061_1[1]), .out(far_5_6061_2[1]));
    assign layer_5[961] = far_5_6061_2[0] & far_5_6061_2[1]; 
    wire [1:0] far_5_6062_0;    relay_conn far_5_6062_0_a(.in(layer_4[650]), .out(far_5_6062_0[0]));    relay_conn far_5_6062_0_b(.in(layer_4[601]), .out(far_5_6062_0[1]));
    assign layer_5[962] = far_5_6062_0[0]; 
    wire [1:0] far_5_6063_0;    relay_conn far_5_6063_0_a(.in(layer_4[176]), .out(far_5_6063_0[0]));    relay_conn far_5_6063_0_b(.in(layer_4[69]), .out(far_5_6063_0[1]));
    wire [1:0] far_5_6063_1;    relay_conn far_5_6063_1_a(.in(far_5_6063_0[0]), .out(far_5_6063_1[0]));    relay_conn far_5_6063_1_b(.in(far_5_6063_0[1]), .out(far_5_6063_1[1]));
    wire [1:0] far_5_6063_2;    relay_conn far_5_6063_2_a(.in(far_5_6063_1[0]), .out(far_5_6063_2[0]));    relay_conn far_5_6063_2_b(.in(far_5_6063_1[1]), .out(far_5_6063_2[1]));
    assign layer_5[963] = ~(far_5_6063_2[0] & far_5_6063_2[1]); 
    wire [1:0] far_5_6064_0;    relay_conn far_5_6064_0_a(.in(layer_4[425]), .out(far_5_6064_0[0]));    relay_conn far_5_6064_0_b(.in(layer_4[333]), .out(far_5_6064_0[1]));
    wire [1:0] far_5_6064_1;    relay_conn far_5_6064_1_a(.in(far_5_6064_0[0]), .out(far_5_6064_1[0]));    relay_conn far_5_6064_1_b(.in(far_5_6064_0[1]), .out(far_5_6064_1[1]));
    assign layer_5[964] = far_5_6064_1[0] & ~far_5_6064_1[1]; 
    wire [1:0] far_5_6065_0;    relay_conn far_5_6065_0_a(.in(layer_4[499]), .out(far_5_6065_0[0]));    relay_conn far_5_6065_0_b(.in(layer_4[608]), .out(far_5_6065_0[1]));
    wire [1:0] far_5_6065_1;    relay_conn far_5_6065_1_a(.in(far_5_6065_0[0]), .out(far_5_6065_1[0]));    relay_conn far_5_6065_1_b(.in(far_5_6065_0[1]), .out(far_5_6065_1[1]));
    wire [1:0] far_5_6065_2;    relay_conn far_5_6065_2_a(.in(far_5_6065_1[0]), .out(far_5_6065_2[0]));    relay_conn far_5_6065_2_b(.in(far_5_6065_1[1]), .out(far_5_6065_2[1]));
    assign layer_5[965] = far_5_6065_2[1] & ~far_5_6065_2[0]; 
    wire [1:0] far_5_6066_0;    relay_conn far_5_6066_0_a(.in(layer_4[898]), .out(far_5_6066_0[0]));    relay_conn far_5_6066_0_b(.in(layer_4[852]), .out(far_5_6066_0[1]));
    assign layer_5[966] = far_5_6066_0[0] & ~far_5_6066_0[1]; 
    assign layer_5[967] = layer_4[562] & ~layer_4[580]; 
    wire [1:0] far_5_6068_0;    relay_conn far_5_6068_0_a(.in(layer_4[955]), .out(far_5_6068_0[0]));    relay_conn far_5_6068_0_b(.in(layer_4[878]), .out(far_5_6068_0[1]));
    wire [1:0] far_5_6068_1;    relay_conn far_5_6068_1_a(.in(far_5_6068_0[0]), .out(far_5_6068_1[0]));    relay_conn far_5_6068_1_b(.in(far_5_6068_0[1]), .out(far_5_6068_1[1]));
    assign layer_5[968] = ~far_5_6068_1[1]; 
    wire [1:0] far_5_6069_0;    relay_conn far_5_6069_0_a(.in(layer_4[13]), .out(far_5_6069_0[0]));    relay_conn far_5_6069_0_b(.in(layer_4[89]), .out(far_5_6069_0[1]));
    wire [1:0] far_5_6069_1;    relay_conn far_5_6069_1_a(.in(far_5_6069_0[0]), .out(far_5_6069_1[0]));    relay_conn far_5_6069_1_b(.in(far_5_6069_0[1]), .out(far_5_6069_1[1]));
    assign layer_5[969] = far_5_6069_1[0] ^ far_5_6069_1[1]; 
    wire [1:0] far_5_6070_0;    relay_conn far_5_6070_0_a(.in(layer_4[186]), .out(far_5_6070_0[0]));    relay_conn far_5_6070_0_b(.in(layer_4[133]), .out(far_5_6070_0[1]));
    assign layer_5[970] = far_5_6070_0[0] & far_5_6070_0[1]; 
    assign layer_5[971] = layer_4[275] & ~layer_4[267]; 
    wire [1:0] far_5_6072_0;    relay_conn far_5_6072_0_a(.in(layer_4[422]), .out(far_5_6072_0[0]));    relay_conn far_5_6072_0_b(.in(layer_4[517]), .out(far_5_6072_0[1]));
    wire [1:0] far_5_6072_1;    relay_conn far_5_6072_1_a(.in(far_5_6072_0[0]), .out(far_5_6072_1[0]));    relay_conn far_5_6072_1_b(.in(far_5_6072_0[1]), .out(far_5_6072_1[1]));
    assign layer_5[972] = ~(far_5_6072_1[0] & far_5_6072_1[1]); 
    wire [1:0] far_5_6073_0;    relay_conn far_5_6073_0_a(.in(layer_4[794]), .out(far_5_6073_0[0]));    relay_conn far_5_6073_0_b(.in(layer_4[759]), .out(far_5_6073_0[1]));
    assign layer_5[973] = ~(far_5_6073_0[0] | far_5_6073_0[1]); 
    wire [1:0] far_5_6074_0;    relay_conn far_5_6074_0_a(.in(layer_4[142]), .out(far_5_6074_0[0]));    relay_conn far_5_6074_0_b(.in(layer_4[43]), .out(far_5_6074_0[1]));
    wire [1:0] far_5_6074_1;    relay_conn far_5_6074_1_a(.in(far_5_6074_0[0]), .out(far_5_6074_1[0]));    relay_conn far_5_6074_1_b(.in(far_5_6074_0[1]), .out(far_5_6074_1[1]));
    wire [1:0] far_5_6074_2;    relay_conn far_5_6074_2_a(.in(far_5_6074_1[0]), .out(far_5_6074_2[0]));    relay_conn far_5_6074_2_b(.in(far_5_6074_1[1]), .out(far_5_6074_2[1]));
    assign layer_5[974] = far_5_6074_2[1] & ~far_5_6074_2[0]; 
    wire [1:0] far_5_6075_0;    relay_conn far_5_6075_0_a(.in(layer_4[653]), .out(far_5_6075_0[0]));    relay_conn far_5_6075_0_b(.in(layer_4[736]), .out(far_5_6075_0[1]));
    wire [1:0] far_5_6075_1;    relay_conn far_5_6075_1_a(.in(far_5_6075_0[0]), .out(far_5_6075_1[0]));    relay_conn far_5_6075_1_b(.in(far_5_6075_0[1]), .out(far_5_6075_1[1]));
    assign layer_5[975] = far_5_6075_1[1] & ~far_5_6075_1[0]; 
    wire [1:0] far_5_6076_0;    relay_conn far_5_6076_0_a(.in(layer_4[489]), .out(far_5_6076_0[0]));    relay_conn far_5_6076_0_b(.in(layer_4[375]), .out(far_5_6076_0[1]));
    wire [1:0] far_5_6076_1;    relay_conn far_5_6076_1_a(.in(far_5_6076_0[0]), .out(far_5_6076_1[0]));    relay_conn far_5_6076_1_b(.in(far_5_6076_0[1]), .out(far_5_6076_1[1]));
    wire [1:0] far_5_6076_2;    relay_conn far_5_6076_2_a(.in(far_5_6076_1[0]), .out(far_5_6076_2[0]));    relay_conn far_5_6076_2_b(.in(far_5_6076_1[1]), .out(far_5_6076_2[1]));
    assign layer_5[976] = far_5_6076_2[0]; 
    assign layer_5[977] = ~layer_4[163]; 
    wire [1:0] far_5_6078_0;    relay_conn far_5_6078_0_a(.in(layer_4[42]), .out(far_5_6078_0[0]));    relay_conn far_5_6078_0_b(.in(layer_4[81]), .out(far_5_6078_0[1]));
    assign layer_5[978] = far_5_6078_0[1]; 
    wire [1:0] far_5_6079_0;    relay_conn far_5_6079_0_a(.in(layer_4[424]), .out(far_5_6079_0[0]));    relay_conn far_5_6079_0_b(.in(layer_4[517]), .out(far_5_6079_0[1]));
    wire [1:0] far_5_6079_1;    relay_conn far_5_6079_1_a(.in(far_5_6079_0[0]), .out(far_5_6079_1[0]));    relay_conn far_5_6079_1_b(.in(far_5_6079_0[1]), .out(far_5_6079_1[1]));
    assign layer_5[979] = far_5_6079_1[1] & ~far_5_6079_1[0]; 
    wire [1:0] far_5_6080_0;    relay_conn far_5_6080_0_a(.in(layer_4[931]), .out(far_5_6080_0[0]));    relay_conn far_5_6080_0_b(.in(layer_4[824]), .out(far_5_6080_0[1]));
    wire [1:0] far_5_6080_1;    relay_conn far_5_6080_1_a(.in(far_5_6080_0[0]), .out(far_5_6080_1[0]));    relay_conn far_5_6080_1_b(.in(far_5_6080_0[1]), .out(far_5_6080_1[1]));
    wire [1:0] far_5_6080_2;    relay_conn far_5_6080_2_a(.in(far_5_6080_1[0]), .out(far_5_6080_2[0]));    relay_conn far_5_6080_2_b(.in(far_5_6080_1[1]), .out(far_5_6080_2[1]));
    assign layer_5[980] = ~far_5_6080_2[1]; 
    wire [1:0] far_5_6081_0;    relay_conn far_5_6081_0_a(.in(layer_4[858]), .out(far_5_6081_0[0]));    relay_conn far_5_6081_0_b(.in(layer_4[775]), .out(far_5_6081_0[1]));
    wire [1:0] far_5_6081_1;    relay_conn far_5_6081_1_a(.in(far_5_6081_0[0]), .out(far_5_6081_1[0]));    relay_conn far_5_6081_1_b(.in(far_5_6081_0[1]), .out(far_5_6081_1[1]));
    assign layer_5[981] = far_5_6081_1[0] & far_5_6081_1[1]; 
    wire [1:0] far_5_6082_0;    relay_conn far_5_6082_0_a(.in(layer_4[354]), .out(far_5_6082_0[0]));    relay_conn far_5_6082_0_b(.in(layer_4[436]), .out(far_5_6082_0[1]));
    wire [1:0] far_5_6082_1;    relay_conn far_5_6082_1_a(.in(far_5_6082_0[0]), .out(far_5_6082_1[0]));    relay_conn far_5_6082_1_b(.in(far_5_6082_0[1]), .out(far_5_6082_1[1]));
    assign layer_5[982] = ~(far_5_6082_1[0] & far_5_6082_1[1]); 
    wire [1:0] far_5_6083_0;    relay_conn far_5_6083_0_a(.in(layer_4[947]), .out(far_5_6083_0[0]));    relay_conn far_5_6083_0_b(.in(layer_4[998]), .out(far_5_6083_0[1]));
    assign layer_5[983] = ~far_5_6083_0[1] | (far_5_6083_0[0] & far_5_6083_0[1]); 
    wire [1:0] far_5_6084_0;    relay_conn far_5_6084_0_a(.in(layer_4[130]), .out(far_5_6084_0[0]));    relay_conn far_5_6084_0_b(.in(layer_4[28]), .out(far_5_6084_0[1]));
    wire [1:0] far_5_6084_1;    relay_conn far_5_6084_1_a(.in(far_5_6084_0[0]), .out(far_5_6084_1[0]));    relay_conn far_5_6084_1_b(.in(far_5_6084_0[1]), .out(far_5_6084_1[1]));
    wire [1:0] far_5_6084_2;    relay_conn far_5_6084_2_a(.in(far_5_6084_1[0]), .out(far_5_6084_2[0]));    relay_conn far_5_6084_2_b(.in(far_5_6084_1[1]), .out(far_5_6084_2[1]));
    assign layer_5[984] = ~(far_5_6084_2[0] & far_5_6084_2[1]); 
    assign layer_5[985] = ~layer_4[499]; 
    wire [1:0] far_5_6086_0;    relay_conn far_5_6086_0_a(.in(layer_4[104]), .out(far_5_6086_0[0]));    relay_conn far_5_6086_0_b(.in(layer_4[224]), .out(far_5_6086_0[1]));
    wire [1:0] far_5_6086_1;    relay_conn far_5_6086_1_a(.in(far_5_6086_0[0]), .out(far_5_6086_1[0]));    relay_conn far_5_6086_1_b(.in(far_5_6086_0[1]), .out(far_5_6086_1[1]));
    wire [1:0] far_5_6086_2;    relay_conn far_5_6086_2_a(.in(far_5_6086_1[0]), .out(far_5_6086_2[0]));    relay_conn far_5_6086_2_b(.in(far_5_6086_1[1]), .out(far_5_6086_2[1]));
    assign layer_5[986] = far_5_6086_2[1] & ~far_5_6086_2[0]; 
    wire [1:0] far_5_6087_0;    relay_conn far_5_6087_0_a(.in(layer_4[454]), .out(far_5_6087_0[0]));    relay_conn far_5_6087_0_b(.in(layer_4[415]), .out(far_5_6087_0[1]));
    assign layer_5[987] = far_5_6087_0[1]; 
    assign layer_5[988] = layer_4[721] ^ layer_4[747]; 
    wire [1:0] far_5_6089_0;    relay_conn far_5_6089_0_a(.in(layer_4[876]), .out(far_5_6089_0[0]));    relay_conn far_5_6089_0_b(.in(layer_4[910]), .out(far_5_6089_0[1]));
    assign layer_5[989] = far_5_6089_0[1]; 
    wire [1:0] far_5_6090_0;    relay_conn far_5_6090_0_a(.in(layer_4[122]), .out(far_5_6090_0[0]));    relay_conn far_5_6090_0_b(.in(layer_4[168]), .out(far_5_6090_0[1]));
    assign layer_5[990] = ~(far_5_6090_0[0] | far_5_6090_0[1]); 
    wire [1:0] far_5_6091_0;    relay_conn far_5_6091_0_a(.in(layer_4[69]), .out(far_5_6091_0[0]));    relay_conn far_5_6091_0_b(.in(layer_4[107]), .out(far_5_6091_0[1]));
    assign layer_5[991] = far_5_6091_0[1]; 
    wire [1:0] far_5_6092_0;    relay_conn far_5_6092_0_a(.in(layer_4[605]), .out(far_5_6092_0[0]));    relay_conn far_5_6092_0_b(.in(layer_4[511]), .out(far_5_6092_0[1]));
    wire [1:0] far_5_6092_1;    relay_conn far_5_6092_1_a(.in(far_5_6092_0[0]), .out(far_5_6092_1[0]));    relay_conn far_5_6092_1_b(.in(far_5_6092_0[1]), .out(far_5_6092_1[1]));
    assign layer_5[992] = far_5_6092_1[0] | far_5_6092_1[1]; 
    assign layer_5[993] = layer_4[508] | layer_4[516]; 
    wire [1:0] far_5_6094_0;    relay_conn far_5_6094_0_a(.in(layer_4[684]), .out(far_5_6094_0[0]));    relay_conn far_5_6094_0_b(.in(layer_4[740]), .out(far_5_6094_0[1]));
    assign layer_5[994] = far_5_6094_0[0] ^ far_5_6094_0[1]; 
    wire [1:0] far_5_6095_0;    relay_conn far_5_6095_0_a(.in(layer_4[1004]), .out(far_5_6095_0[0]));    relay_conn far_5_6095_0_b(.in(layer_4[902]), .out(far_5_6095_0[1]));
    wire [1:0] far_5_6095_1;    relay_conn far_5_6095_1_a(.in(far_5_6095_0[0]), .out(far_5_6095_1[0]));    relay_conn far_5_6095_1_b(.in(far_5_6095_0[1]), .out(far_5_6095_1[1]));
    wire [1:0] far_5_6095_2;    relay_conn far_5_6095_2_a(.in(far_5_6095_1[0]), .out(far_5_6095_2[0]));    relay_conn far_5_6095_2_b(.in(far_5_6095_1[1]), .out(far_5_6095_2[1]));
    assign layer_5[995] = far_5_6095_2[0]; 
    wire [1:0] far_5_6096_0;    relay_conn far_5_6096_0_a(.in(layer_4[499]), .out(far_5_6096_0[0]));    relay_conn far_5_6096_0_b(.in(layer_4[558]), .out(far_5_6096_0[1]));
    assign layer_5[996] = far_5_6096_0[0] & ~far_5_6096_0[1]; 
    assign layer_5[997] = ~(layer_4[603] | layer_4[589]); 
    wire [1:0] far_5_6098_0;    relay_conn far_5_6098_0_a(.in(layer_4[266]), .out(far_5_6098_0[0]));    relay_conn far_5_6098_0_b(.in(layer_4[369]), .out(far_5_6098_0[1]));
    wire [1:0] far_5_6098_1;    relay_conn far_5_6098_1_a(.in(far_5_6098_0[0]), .out(far_5_6098_1[0]));    relay_conn far_5_6098_1_b(.in(far_5_6098_0[1]), .out(far_5_6098_1[1]));
    wire [1:0] far_5_6098_2;    relay_conn far_5_6098_2_a(.in(far_5_6098_1[0]), .out(far_5_6098_2[0]));    relay_conn far_5_6098_2_b(.in(far_5_6098_1[1]), .out(far_5_6098_2[1]));
    assign layer_5[998] = ~far_5_6098_2[1] | (far_5_6098_2[0] & far_5_6098_2[1]); 
    wire [1:0] far_5_6099_0;    relay_conn far_5_6099_0_a(.in(layer_4[795]), .out(far_5_6099_0[0]));    relay_conn far_5_6099_0_b(.in(layer_4[872]), .out(far_5_6099_0[1]));
    wire [1:0] far_5_6099_1;    relay_conn far_5_6099_1_a(.in(far_5_6099_0[0]), .out(far_5_6099_1[0]));    relay_conn far_5_6099_1_b(.in(far_5_6099_0[1]), .out(far_5_6099_1[1]));
    assign layer_5[999] = ~far_5_6099_1[0] | (far_5_6099_1[0] & far_5_6099_1[1]); 
    wire [1:0] far_5_6100_0;    relay_conn far_5_6100_0_a(.in(layer_4[136]), .out(far_5_6100_0[0]));    relay_conn far_5_6100_0_b(.in(layer_4[172]), .out(far_5_6100_0[1]));
    assign layer_5[1000] = ~far_5_6100_0[0] | (far_5_6100_0[0] & far_5_6100_0[1]); 
    assign layer_5[1001] = ~(layer_4[978] | layer_4[947]); 
    assign layer_5[1002] = ~layer_4[182]; 
    wire [1:0] far_5_6103_0;    relay_conn far_5_6103_0_a(.in(layer_4[650]), .out(far_5_6103_0[0]));    relay_conn far_5_6103_0_b(.in(layer_4[605]), .out(far_5_6103_0[1]));
    assign layer_5[1003] = far_5_6103_0[0]; 
    assign layer_5[1004] = layer_4[295] & layer_4[285]; 
    assign layer_5[1005] = layer_4[538] | layer_4[516]; 
    wire [1:0] far_5_6106_0;    relay_conn far_5_6106_0_a(.in(layer_4[580]), .out(far_5_6106_0[0]));    relay_conn far_5_6106_0_b(.in(layer_4[614]), .out(far_5_6106_0[1]));
    assign layer_5[1006] = far_5_6106_0[0] ^ far_5_6106_0[1]; 
    assign layer_5[1007] = layer_4[559]; 
    wire [1:0] far_5_6108_0;    relay_conn far_5_6108_0_a(.in(layer_4[365]), .out(far_5_6108_0[0]));    relay_conn far_5_6108_0_b(.in(layer_4[473]), .out(far_5_6108_0[1]));
    wire [1:0] far_5_6108_1;    relay_conn far_5_6108_1_a(.in(far_5_6108_0[0]), .out(far_5_6108_1[0]));    relay_conn far_5_6108_1_b(.in(far_5_6108_0[1]), .out(far_5_6108_1[1]));
    wire [1:0] far_5_6108_2;    relay_conn far_5_6108_2_a(.in(far_5_6108_1[0]), .out(far_5_6108_2[0]));    relay_conn far_5_6108_2_b(.in(far_5_6108_1[1]), .out(far_5_6108_2[1]));
    assign layer_5[1008] = far_5_6108_2[0] | far_5_6108_2[1]; 
    assign layer_5[1009] = layer_4[314] & layer_4[306]; 
    wire [1:0] far_5_6110_0;    relay_conn far_5_6110_0_a(.in(layer_4[296]), .out(far_5_6110_0[0]));    relay_conn far_5_6110_0_b(.in(layer_4[384]), .out(far_5_6110_0[1]));
    wire [1:0] far_5_6110_1;    relay_conn far_5_6110_1_a(.in(far_5_6110_0[0]), .out(far_5_6110_1[0]));    relay_conn far_5_6110_1_b(.in(far_5_6110_0[1]), .out(far_5_6110_1[1]));
    assign layer_5[1010] = ~far_5_6110_1[1]; 
    wire [1:0] far_5_6111_0;    relay_conn far_5_6111_0_a(.in(layer_4[916]), .out(far_5_6111_0[0]));    relay_conn far_5_6111_0_b(.in(layer_4[815]), .out(far_5_6111_0[1]));
    wire [1:0] far_5_6111_1;    relay_conn far_5_6111_1_a(.in(far_5_6111_0[0]), .out(far_5_6111_1[0]));    relay_conn far_5_6111_1_b(.in(far_5_6111_0[1]), .out(far_5_6111_1[1]));
    wire [1:0] far_5_6111_2;    relay_conn far_5_6111_2_a(.in(far_5_6111_1[0]), .out(far_5_6111_2[0]));    relay_conn far_5_6111_2_b(.in(far_5_6111_1[1]), .out(far_5_6111_2[1]));
    assign layer_5[1011] = ~(far_5_6111_2[0] | far_5_6111_2[1]); 
    wire [1:0] far_5_6112_0;    relay_conn far_5_6112_0_a(.in(layer_4[401]), .out(far_5_6112_0[0]));    relay_conn far_5_6112_0_b(.in(layer_4[517]), .out(far_5_6112_0[1]));
    wire [1:0] far_5_6112_1;    relay_conn far_5_6112_1_a(.in(far_5_6112_0[0]), .out(far_5_6112_1[0]));    relay_conn far_5_6112_1_b(.in(far_5_6112_0[1]), .out(far_5_6112_1[1]));
    wire [1:0] far_5_6112_2;    relay_conn far_5_6112_2_a(.in(far_5_6112_1[0]), .out(far_5_6112_2[0]));    relay_conn far_5_6112_2_b(.in(far_5_6112_1[1]), .out(far_5_6112_2[1]));
    assign layer_5[1012] = ~far_5_6112_2[1] | (far_5_6112_2[0] & far_5_6112_2[1]); 
    wire [1:0] far_5_6113_0;    relay_conn far_5_6113_0_a(.in(layer_4[366]), .out(far_5_6113_0[0]));    relay_conn far_5_6113_0_b(.in(layer_4[422]), .out(far_5_6113_0[1]));
    assign layer_5[1013] = ~far_5_6113_0[0] | (far_5_6113_0[0] & far_5_6113_0[1]); 
    wire [1:0] far_5_6114_0;    relay_conn far_5_6114_0_a(.in(layer_4[869]), .out(far_5_6114_0[0]));    relay_conn far_5_6114_0_b(.in(layer_4[806]), .out(far_5_6114_0[1]));
    assign layer_5[1014] = far_5_6114_0[0] & ~far_5_6114_0[1]; 
    wire [1:0] far_5_6115_0;    relay_conn far_5_6115_0_a(.in(layer_4[175]), .out(far_5_6115_0[0]));    relay_conn far_5_6115_0_b(.in(layer_4[215]), .out(far_5_6115_0[1]));
    assign layer_5[1015] = far_5_6115_0[1]; 
    wire [1:0] far_5_6116_0;    relay_conn far_5_6116_0_a(.in(layer_4[983]), .out(far_5_6116_0[0]));    relay_conn far_5_6116_0_b(.in(layer_4[906]), .out(far_5_6116_0[1]));
    wire [1:0] far_5_6116_1;    relay_conn far_5_6116_1_a(.in(far_5_6116_0[0]), .out(far_5_6116_1[0]));    relay_conn far_5_6116_1_b(.in(far_5_6116_0[1]), .out(far_5_6116_1[1]));
    assign layer_5[1016] = ~far_5_6116_1[0]; 
    wire [1:0] far_5_6117_0;    relay_conn far_5_6117_0_a(.in(layer_4[913]), .out(far_5_6117_0[0]));    relay_conn far_5_6117_0_b(.in(layer_4[954]), .out(far_5_6117_0[1]));
    assign layer_5[1017] = ~far_5_6117_0[0] | (far_5_6117_0[0] & far_5_6117_0[1]); 
    wire [1:0] far_5_6118_0;    relay_conn far_5_6118_0_a(.in(layer_4[542]), .out(far_5_6118_0[0]));    relay_conn far_5_6118_0_b(.in(layer_4[632]), .out(far_5_6118_0[1]));
    wire [1:0] far_5_6118_1;    relay_conn far_5_6118_1_a(.in(far_5_6118_0[0]), .out(far_5_6118_1[0]));    relay_conn far_5_6118_1_b(.in(far_5_6118_0[1]), .out(far_5_6118_1[1]));
    assign layer_5[1018] = far_5_6118_1[0] | far_5_6118_1[1]; 
    assign layer_5[1019] = ~layer_4[619]; 
    // Layer 6 ============================================================
    assign layer_6[0] = ~(layer_5[983] ^ layer_5[960]); 
    wire [1:0] far_6_6121_0;    relay_conn far_6_6121_0_a(.in(layer_5[273]), .out(far_6_6121_0[0]));    relay_conn far_6_6121_0_b(.in(layer_5[180]), .out(far_6_6121_0[1]));
    wire [1:0] far_6_6121_1;    relay_conn far_6_6121_1_a(.in(far_6_6121_0[0]), .out(far_6_6121_1[0]));    relay_conn far_6_6121_1_b(.in(far_6_6121_0[1]), .out(far_6_6121_1[1]));
    assign layer_6[1] = ~far_6_6121_1[0]; 
    wire [1:0] far_6_6122_0;    relay_conn far_6_6122_0_a(.in(layer_5[477]), .out(far_6_6122_0[0]));    relay_conn far_6_6122_0_b(.in(layer_5[599]), .out(far_6_6122_0[1]));
    wire [1:0] far_6_6122_1;    relay_conn far_6_6122_1_a(.in(far_6_6122_0[0]), .out(far_6_6122_1[0]));    relay_conn far_6_6122_1_b(.in(far_6_6122_0[1]), .out(far_6_6122_1[1]));
    wire [1:0] far_6_6122_2;    relay_conn far_6_6122_2_a(.in(far_6_6122_1[0]), .out(far_6_6122_2[0]));    relay_conn far_6_6122_2_b(.in(far_6_6122_1[1]), .out(far_6_6122_2[1]));
    assign layer_6[2] = far_6_6122_2[0] | far_6_6122_2[1]; 
    wire [1:0] far_6_6123_0;    relay_conn far_6_6123_0_a(.in(layer_5[269]), .out(far_6_6123_0[0]));    relay_conn far_6_6123_0_b(.in(layer_5[158]), .out(far_6_6123_0[1]));
    wire [1:0] far_6_6123_1;    relay_conn far_6_6123_1_a(.in(far_6_6123_0[0]), .out(far_6_6123_1[0]));    relay_conn far_6_6123_1_b(.in(far_6_6123_0[1]), .out(far_6_6123_1[1]));
    wire [1:0] far_6_6123_2;    relay_conn far_6_6123_2_a(.in(far_6_6123_1[0]), .out(far_6_6123_2[0]));    relay_conn far_6_6123_2_b(.in(far_6_6123_1[1]), .out(far_6_6123_2[1]));
    assign layer_6[3] = far_6_6123_2[0] | far_6_6123_2[1]; 
    wire [1:0] far_6_6124_0;    relay_conn far_6_6124_0_a(.in(layer_5[734]), .out(far_6_6124_0[0]));    relay_conn far_6_6124_0_b(.in(layer_5[617]), .out(far_6_6124_0[1]));
    wire [1:0] far_6_6124_1;    relay_conn far_6_6124_1_a(.in(far_6_6124_0[0]), .out(far_6_6124_1[0]));    relay_conn far_6_6124_1_b(.in(far_6_6124_0[1]), .out(far_6_6124_1[1]));
    wire [1:0] far_6_6124_2;    relay_conn far_6_6124_2_a(.in(far_6_6124_1[0]), .out(far_6_6124_2[0]));    relay_conn far_6_6124_2_b(.in(far_6_6124_1[1]), .out(far_6_6124_2[1]));
    assign layer_6[4] = far_6_6124_2[1] & ~far_6_6124_2[0]; 
    wire [1:0] far_6_6125_0;    relay_conn far_6_6125_0_a(.in(layer_5[720]), .out(far_6_6125_0[0]));    relay_conn far_6_6125_0_b(.in(layer_5[604]), .out(far_6_6125_0[1]));
    wire [1:0] far_6_6125_1;    relay_conn far_6_6125_1_a(.in(far_6_6125_0[0]), .out(far_6_6125_1[0]));    relay_conn far_6_6125_1_b(.in(far_6_6125_0[1]), .out(far_6_6125_1[1]));
    wire [1:0] far_6_6125_2;    relay_conn far_6_6125_2_a(.in(far_6_6125_1[0]), .out(far_6_6125_2[0]));    relay_conn far_6_6125_2_b(.in(far_6_6125_1[1]), .out(far_6_6125_2[1]));
    assign layer_6[5] = far_6_6125_2[0] & far_6_6125_2[1]; 
    wire [1:0] far_6_6126_0;    relay_conn far_6_6126_0_a(.in(layer_5[698]), .out(far_6_6126_0[0]));    relay_conn far_6_6126_0_b(.in(layer_5[665]), .out(far_6_6126_0[1]));
    assign layer_6[6] = ~far_6_6126_0[0] | (far_6_6126_0[0] & far_6_6126_0[1]); 
    wire [1:0] far_6_6127_0;    relay_conn far_6_6127_0_a(.in(layer_5[325]), .out(far_6_6127_0[0]));    relay_conn far_6_6127_0_b(.in(layer_5[415]), .out(far_6_6127_0[1]));
    wire [1:0] far_6_6127_1;    relay_conn far_6_6127_1_a(.in(far_6_6127_0[0]), .out(far_6_6127_1[0]));    relay_conn far_6_6127_1_b(.in(far_6_6127_0[1]), .out(far_6_6127_1[1]));
    assign layer_6[7] = ~far_6_6127_1[1]; 
    wire [1:0] far_6_6128_0;    relay_conn far_6_6128_0_a(.in(layer_5[313]), .out(far_6_6128_0[0]));    relay_conn far_6_6128_0_b(.in(layer_5[219]), .out(far_6_6128_0[1]));
    wire [1:0] far_6_6128_1;    relay_conn far_6_6128_1_a(.in(far_6_6128_0[0]), .out(far_6_6128_1[0]));    relay_conn far_6_6128_1_b(.in(far_6_6128_0[1]), .out(far_6_6128_1[1]));
    assign layer_6[8] = far_6_6128_1[0] ^ far_6_6128_1[1]; 
    wire [1:0] far_6_6129_0;    relay_conn far_6_6129_0_a(.in(layer_5[218]), .out(far_6_6129_0[0]));    relay_conn far_6_6129_0_b(.in(layer_5[150]), .out(far_6_6129_0[1]));
    wire [1:0] far_6_6129_1;    relay_conn far_6_6129_1_a(.in(far_6_6129_0[0]), .out(far_6_6129_1[0]));    relay_conn far_6_6129_1_b(.in(far_6_6129_0[1]), .out(far_6_6129_1[1]));
    assign layer_6[9] = ~far_6_6129_1[1]; 
    wire [1:0] far_6_6130_0;    relay_conn far_6_6130_0_a(.in(layer_5[777]), .out(far_6_6130_0[0]));    relay_conn far_6_6130_0_b(.in(layer_5[855]), .out(far_6_6130_0[1]));
    wire [1:0] far_6_6130_1;    relay_conn far_6_6130_1_a(.in(far_6_6130_0[0]), .out(far_6_6130_1[0]));    relay_conn far_6_6130_1_b(.in(far_6_6130_0[1]), .out(far_6_6130_1[1]));
    assign layer_6[10] = far_6_6130_1[0] & far_6_6130_1[1]; 
    wire [1:0] far_6_6131_0;    relay_conn far_6_6131_0_a(.in(layer_5[666]), .out(far_6_6131_0[0]));    relay_conn far_6_6131_0_b(.in(layer_5[613]), .out(far_6_6131_0[1]));
    assign layer_6[11] = ~far_6_6131_0[0]; 
    wire [1:0] far_6_6132_0;    relay_conn far_6_6132_0_a(.in(layer_5[330]), .out(far_6_6132_0[0]));    relay_conn far_6_6132_0_b(.in(layer_5[445]), .out(far_6_6132_0[1]));
    wire [1:0] far_6_6132_1;    relay_conn far_6_6132_1_a(.in(far_6_6132_0[0]), .out(far_6_6132_1[0]));    relay_conn far_6_6132_1_b(.in(far_6_6132_0[1]), .out(far_6_6132_1[1]));
    wire [1:0] far_6_6132_2;    relay_conn far_6_6132_2_a(.in(far_6_6132_1[0]), .out(far_6_6132_2[0]));    relay_conn far_6_6132_2_b(.in(far_6_6132_1[1]), .out(far_6_6132_2[1]));
    assign layer_6[12] = far_6_6132_2[0] | far_6_6132_2[1]; 
    assign layer_6[13] = layer_5[996]; 
    wire [1:0] far_6_6134_0;    relay_conn far_6_6134_0_a(.in(layer_5[634]), .out(far_6_6134_0[0]));    relay_conn far_6_6134_0_b(.in(layer_5[584]), .out(far_6_6134_0[1]));
    assign layer_6[14] = far_6_6134_0[0] & far_6_6134_0[1]; 
    assign layer_6[15] = layer_5[77]; 
    assign layer_6[16] = ~(layer_5[894] ^ layer_5[919]); 
    assign layer_6[17] = ~layer_5[67] | (layer_5[52] & layer_5[67]); 
    wire [1:0] far_6_6138_0;    relay_conn far_6_6138_0_a(.in(layer_5[860]), .out(far_6_6138_0[0]));    relay_conn far_6_6138_0_b(.in(layer_5[763]), .out(far_6_6138_0[1]));
    wire [1:0] far_6_6138_1;    relay_conn far_6_6138_1_a(.in(far_6_6138_0[0]), .out(far_6_6138_1[0]));    relay_conn far_6_6138_1_b(.in(far_6_6138_0[1]), .out(far_6_6138_1[1]));
    wire [1:0] far_6_6138_2;    relay_conn far_6_6138_2_a(.in(far_6_6138_1[0]), .out(far_6_6138_2[0]));    relay_conn far_6_6138_2_b(.in(far_6_6138_1[1]), .out(far_6_6138_2[1]));
    assign layer_6[18] = ~far_6_6138_2[1] | (far_6_6138_2[0] & far_6_6138_2[1]); 
    wire [1:0] far_6_6139_0;    relay_conn far_6_6139_0_a(.in(layer_5[944]), .out(far_6_6139_0[0]));    relay_conn far_6_6139_0_b(.in(layer_5[857]), .out(far_6_6139_0[1]));
    wire [1:0] far_6_6139_1;    relay_conn far_6_6139_1_a(.in(far_6_6139_0[0]), .out(far_6_6139_1[0]));    relay_conn far_6_6139_1_b(.in(far_6_6139_0[1]), .out(far_6_6139_1[1]));
    assign layer_6[19] = ~far_6_6139_1[1] | (far_6_6139_1[0] & far_6_6139_1[1]); 
    wire [1:0] far_6_6140_0;    relay_conn far_6_6140_0_a(.in(layer_5[849]), .out(far_6_6140_0[0]));    relay_conn far_6_6140_0_b(.in(layer_5[891]), .out(far_6_6140_0[1]));
    assign layer_6[20] = ~far_6_6140_0[1] | (far_6_6140_0[0] & far_6_6140_0[1]); 
    assign layer_6[21] = ~layer_5[464]; 
    assign layer_6[22] = ~(layer_5[563] | layer_5[552]); 
    wire [1:0] far_6_6143_0;    relay_conn far_6_6143_0_a(.in(layer_5[660]), .out(far_6_6143_0[0]));    relay_conn far_6_6143_0_b(.in(layer_5[776]), .out(far_6_6143_0[1]));
    wire [1:0] far_6_6143_1;    relay_conn far_6_6143_1_a(.in(far_6_6143_0[0]), .out(far_6_6143_1[0]));    relay_conn far_6_6143_1_b(.in(far_6_6143_0[1]), .out(far_6_6143_1[1]));
    wire [1:0] far_6_6143_2;    relay_conn far_6_6143_2_a(.in(far_6_6143_1[0]), .out(far_6_6143_2[0]));    relay_conn far_6_6143_2_b(.in(far_6_6143_1[1]), .out(far_6_6143_2[1]));
    assign layer_6[23] = ~(far_6_6143_2[0] ^ far_6_6143_2[1]); 
    wire [1:0] far_6_6144_0;    relay_conn far_6_6144_0_a(.in(layer_5[360]), .out(far_6_6144_0[0]));    relay_conn far_6_6144_0_b(.in(layer_5[396]), .out(far_6_6144_0[1]));
    assign layer_6[24] = far_6_6144_0[0]; 
    wire [1:0] far_6_6145_0;    relay_conn far_6_6145_0_a(.in(layer_5[234]), .out(far_6_6145_0[0]));    relay_conn far_6_6145_0_b(.in(layer_5[178]), .out(far_6_6145_0[1]));
    assign layer_6[25] = ~far_6_6145_0[1]; 
    wire [1:0] far_6_6146_0;    relay_conn far_6_6146_0_a(.in(layer_5[189]), .out(far_6_6146_0[0]));    relay_conn far_6_6146_0_b(.in(layer_5[283]), .out(far_6_6146_0[1]));
    wire [1:0] far_6_6146_1;    relay_conn far_6_6146_1_a(.in(far_6_6146_0[0]), .out(far_6_6146_1[0]));    relay_conn far_6_6146_1_b(.in(far_6_6146_0[1]), .out(far_6_6146_1[1]));
    assign layer_6[26] = far_6_6146_1[0] & far_6_6146_1[1]; 
    wire [1:0] far_6_6147_0;    relay_conn far_6_6147_0_a(.in(layer_5[544]), .out(far_6_6147_0[0]));    relay_conn far_6_6147_0_b(.in(layer_5[598]), .out(far_6_6147_0[1]));
    assign layer_6[27] = ~far_6_6147_0[1]; 
    assign layer_6[28] = ~layer_5[761]; 
    assign layer_6[29] = layer_5[922] & layer_5[952]; 
    wire [1:0] far_6_6150_0;    relay_conn far_6_6150_0_a(.in(layer_5[636]), .out(far_6_6150_0[0]));    relay_conn far_6_6150_0_b(.in(layer_5[562]), .out(far_6_6150_0[1]));
    wire [1:0] far_6_6150_1;    relay_conn far_6_6150_1_a(.in(far_6_6150_0[0]), .out(far_6_6150_1[0]));    relay_conn far_6_6150_1_b(.in(far_6_6150_0[1]), .out(far_6_6150_1[1]));
    assign layer_6[30] = far_6_6150_1[0] | far_6_6150_1[1]; 
    wire [1:0] far_6_6151_0;    relay_conn far_6_6151_0_a(.in(layer_5[348]), .out(far_6_6151_0[0]));    relay_conn far_6_6151_0_b(.in(layer_5[222]), .out(far_6_6151_0[1]));
    wire [1:0] far_6_6151_1;    relay_conn far_6_6151_1_a(.in(far_6_6151_0[0]), .out(far_6_6151_1[0]));    relay_conn far_6_6151_1_b(.in(far_6_6151_0[1]), .out(far_6_6151_1[1]));
    wire [1:0] far_6_6151_2;    relay_conn far_6_6151_2_a(.in(far_6_6151_1[0]), .out(far_6_6151_2[0]));    relay_conn far_6_6151_2_b(.in(far_6_6151_1[1]), .out(far_6_6151_2[1]));
    assign layer_6[31] = ~(far_6_6151_2[0] | far_6_6151_2[1]); 
    wire [1:0] far_6_6152_0;    relay_conn far_6_6152_0_a(.in(layer_5[607]), .out(far_6_6152_0[0]));    relay_conn far_6_6152_0_b(.in(layer_5[668]), .out(far_6_6152_0[1]));
    assign layer_6[32] = far_6_6152_0[0]; 
    wire [1:0] far_6_6153_0;    relay_conn far_6_6153_0_a(.in(layer_5[282]), .out(far_6_6153_0[0]));    relay_conn far_6_6153_0_b(.in(layer_5[158]), .out(far_6_6153_0[1]));
    wire [1:0] far_6_6153_1;    relay_conn far_6_6153_1_a(.in(far_6_6153_0[0]), .out(far_6_6153_1[0]));    relay_conn far_6_6153_1_b(.in(far_6_6153_0[1]), .out(far_6_6153_1[1]));
    wire [1:0] far_6_6153_2;    relay_conn far_6_6153_2_a(.in(far_6_6153_1[0]), .out(far_6_6153_2[0]));    relay_conn far_6_6153_2_b(.in(far_6_6153_1[1]), .out(far_6_6153_2[1]));
    assign layer_6[33] = ~far_6_6153_2[0] | (far_6_6153_2[0] & far_6_6153_2[1]); 
    assign layer_6[34] = ~layer_5[944] | (layer_5[944] & layer_5[967]); 
    assign layer_6[35] = layer_5[956] & ~layer_5[981]; 
    wire [1:0] far_6_6156_0;    relay_conn far_6_6156_0_a(.in(layer_5[364]), .out(far_6_6156_0[0]));    relay_conn far_6_6156_0_b(.in(layer_5[489]), .out(far_6_6156_0[1]));
    wire [1:0] far_6_6156_1;    relay_conn far_6_6156_1_a(.in(far_6_6156_0[0]), .out(far_6_6156_1[0]));    relay_conn far_6_6156_1_b(.in(far_6_6156_0[1]), .out(far_6_6156_1[1]));
    wire [1:0] far_6_6156_2;    relay_conn far_6_6156_2_a(.in(far_6_6156_1[0]), .out(far_6_6156_2[0]));    relay_conn far_6_6156_2_b(.in(far_6_6156_1[1]), .out(far_6_6156_2[1]));
    assign layer_6[36] = far_6_6156_2[0] ^ far_6_6156_2[1]; 
    assign layer_6[37] = layer_5[130] & ~layer_5[128]; 
    wire [1:0] far_6_6158_0;    relay_conn far_6_6158_0_a(.in(layer_5[576]), .out(far_6_6158_0[0]));    relay_conn far_6_6158_0_b(.in(layer_5[675]), .out(far_6_6158_0[1]));
    wire [1:0] far_6_6158_1;    relay_conn far_6_6158_1_a(.in(far_6_6158_0[0]), .out(far_6_6158_1[0]));    relay_conn far_6_6158_1_b(.in(far_6_6158_0[1]), .out(far_6_6158_1[1]));
    wire [1:0] far_6_6158_2;    relay_conn far_6_6158_2_a(.in(far_6_6158_1[0]), .out(far_6_6158_2[0]));    relay_conn far_6_6158_2_b(.in(far_6_6158_1[1]), .out(far_6_6158_2[1]));
    assign layer_6[38] = ~far_6_6158_2[1]; 
    assign layer_6[39] = ~layer_5[772]; 
    wire [1:0] far_6_6160_0;    relay_conn far_6_6160_0_a(.in(layer_5[284]), .out(far_6_6160_0[0]));    relay_conn far_6_6160_0_b(.in(layer_5[231]), .out(far_6_6160_0[1]));
    assign layer_6[40] = ~far_6_6160_0[1]; 
    assign layer_6[41] = ~layer_5[932] | (layer_5[932] & layer_5[956]); 
    wire [1:0] far_6_6162_0;    relay_conn far_6_6162_0_a(.in(layer_5[216]), .out(far_6_6162_0[0]));    relay_conn far_6_6162_0_b(.in(layer_5[125]), .out(far_6_6162_0[1]));
    wire [1:0] far_6_6162_1;    relay_conn far_6_6162_1_a(.in(far_6_6162_0[0]), .out(far_6_6162_1[0]));    relay_conn far_6_6162_1_b(.in(far_6_6162_0[1]), .out(far_6_6162_1[1]));
    assign layer_6[42] = ~(far_6_6162_1[0] | far_6_6162_1[1]); 
    wire [1:0] far_6_6163_0;    relay_conn far_6_6163_0_a(.in(layer_5[366]), .out(far_6_6163_0[0]));    relay_conn far_6_6163_0_b(.in(layer_5[423]), .out(far_6_6163_0[1]));
    assign layer_6[43] = ~far_6_6163_0[1] | (far_6_6163_0[0] & far_6_6163_0[1]); 
    wire [1:0] far_6_6164_0;    relay_conn far_6_6164_0_a(.in(layer_5[746]), .out(far_6_6164_0[0]));    relay_conn far_6_6164_0_b(.in(layer_5[706]), .out(far_6_6164_0[1]));
    assign layer_6[44] = far_6_6164_0[0] & ~far_6_6164_0[1]; 
    wire [1:0] far_6_6165_0;    relay_conn far_6_6165_0_a(.in(layer_5[124]), .out(far_6_6165_0[0]));    relay_conn far_6_6165_0_b(.in(layer_5[22]), .out(far_6_6165_0[1]));
    wire [1:0] far_6_6165_1;    relay_conn far_6_6165_1_a(.in(far_6_6165_0[0]), .out(far_6_6165_1[0]));    relay_conn far_6_6165_1_b(.in(far_6_6165_0[1]), .out(far_6_6165_1[1]));
    wire [1:0] far_6_6165_2;    relay_conn far_6_6165_2_a(.in(far_6_6165_1[0]), .out(far_6_6165_2[0]));    relay_conn far_6_6165_2_b(.in(far_6_6165_1[1]), .out(far_6_6165_2[1]));
    assign layer_6[45] = far_6_6165_2[0] & far_6_6165_2[1]; 
    wire [1:0] far_6_6166_0;    relay_conn far_6_6166_0_a(.in(layer_5[91]), .out(far_6_6166_0[0]));    relay_conn far_6_6166_0_b(.in(layer_5[194]), .out(far_6_6166_0[1]));
    wire [1:0] far_6_6166_1;    relay_conn far_6_6166_1_a(.in(far_6_6166_0[0]), .out(far_6_6166_1[0]));    relay_conn far_6_6166_1_b(.in(far_6_6166_0[1]), .out(far_6_6166_1[1]));
    wire [1:0] far_6_6166_2;    relay_conn far_6_6166_2_a(.in(far_6_6166_1[0]), .out(far_6_6166_2[0]));    relay_conn far_6_6166_2_b(.in(far_6_6166_1[1]), .out(far_6_6166_2[1]));
    assign layer_6[46] = far_6_6166_2[0] | far_6_6166_2[1]; 
    wire [1:0] far_6_6167_0;    relay_conn far_6_6167_0_a(.in(layer_5[845]), .out(far_6_6167_0[0]));    relay_conn far_6_6167_0_b(.in(layer_5[772]), .out(far_6_6167_0[1]));
    wire [1:0] far_6_6167_1;    relay_conn far_6_6167_1_a(.in(far_6_6167_0[0]), .out(far_6_6167_1[0]));    relay_conn far_6_6167_1_b(.in(far_6_6167_0[1]), .out(far_6_6167_1[1]));
    assign layer_6[47] = far_6_6167_1[0]; 
    assign layer_6[48] = ~layer_5[44]; 
    wire [1:0] far_6_6169_0;    relay_conn far_6_6169_0_a(.in(layer_5[436]), .out(far_6_6169_0[0]));    relay_conn far_6_6169_0_b(.in(layer_5[473]), .out(far_6_6169_0[1]));
    assign layer_6[49] = ~(far_6_6169_0[0] & far_6_6169_0[1]); 
    wire [1:0] far_6_6170_0;    relay_conn far_6_6170_0_a(.in(layer_5[31]), .out(far_6_6170_0[0]));    relay_conn far_6_6170_0_b(.in(layer_5[63]), .out(far_6_6170_0[1]));
    assign layer_6[50] = far_6_6170_0[0] | far_6_6170_0[1]; 
    wire [1:0] far_6_6171_0;    relay_conn far_6_6171_0_a(.in(layer_5[748]), .out(far_6_6171_0[0]));    relay_conn far_6_6171_0_b(.in(layer_5[837]), .out(far_6_6171_0[1]));
    wire [1:0] far_6_6171_1;    relay_conn far_6_6171_1_a(.in(far_6_6171_0[0]), .out(far_6_6171_1[0]));    relay_conn far_6_6171_1_b(.in(far_6_6171_0[1]), .out(far_6_6171_1[1]));
    assign layer_6[51] = ~far_6_6171_1[0]; 
    wire [1:0] far_6_6172_0;    relay_conn far_6_6172_0_a(.in(layer_5[44]), .out(far_6_6172_0[0]));    relay_conn far_6_6172_0_b(.in(layer_5[150]), .out(far_6_6172_0[1]));
    wire [1:0] far_6_6172_1;    relay_conn far_6_6172_1_a(.in(far_6_6172_0[0]), .out(far_6_6172_1[0]));    relay_conn far_6_6172_1_b(.in(far_6_6172_0[1]), .out(far_6_6172_1[1]));
    wire [1:0] far_6_6172_2;    relay_conn far_6_6172_2_a(.in(far_6_6172_1[0]), .out(far_6_6172_2[0]));    relay_conn far_6_6172_2_b(.in(far_6_6172_1[1]), .out(far_6_6172_2[1]));
    assign layer_6[52] = far_6_6172_2[0] ^ far_6_6172_2[1]; 
    wire [1:0] far_6_6173_0;    relay_conn far_6_6173_0_a(.in(layer_5[751]), .out(far_6_6173_0[0]));    relay_conn far_6_6173_0_b(.in(layer_5[689]), .out(far_6_6173_0[1]));
    assign layer_6[53] = ~far_6_6173_0[1]; 
    assign layer_6[54] = ~layer_5[917]; 
    wire [1:0] far_6_6175_0;    relay_conn far_6_6175_0_a(.in(layer_5[974]), .out(far_6_6175_0[0]));    relay_conn far_6_6175_0_b(.in(layer_5[886]), .out(far_6_6175_0[1]));
    wire [1:0] far_6_6175_1;    relay_conn far_6_6175_1_a(.in(far_6_6175_0[0]), .out(far_6_6175_1[0]));    relay_conn far_6_6175_1_b(.in(far_6_6175_0[1]), .out(far_6_6175_1[1]));
    assign layer_6[55] = ~(far_6_6175_1[0] & far_6_6175_1[1]); 
    wire [1:0] far_6_6176_0;    relay_conn far_6_6176_0_a(.in(layer_5[236]), .out(far_6_6176_0[0]));    relay_conn far_6_6176_0_b(.in(layer_5[355]), .out(far_6_6176_0[1]));
    wire [1:0] far_6_6176_1;    relay_conn far_6_6176_1_a(.in(far_6_6176_0[0]), .out(far_6_6176_1[0]));    relay_conn far_6_6176_1_b(.in(far_6_6176_0[1]), .out(far_6_6176_1[1]));
    wire [1:0] far_6_6176_2;    relay_conn far_6_6176_2_a(.in(far_6_6176_1[0]), .out(far_6_6176_2[0]));    relay_conn far_6_6176_2_b(.in(far_6_6176_1[1]), .out(far_6_6176_2[1]));
    assign layer_6[56] = ~far_6_6176_2[0] | (far_6_6176_2[0] & far_6_6176_2[1]); 
    wire [1:0] far_6_6177_0;    relay_conn far_6_6177_0_a(.in(layer_5[282]), .out(far_6_6177_0[0]));    relay_conn far_6_6177_0_b(.in(layer_5[348]), .out(far_6_6177_0[1]));
    wire [1:0] far_6_6177_1;    relay_conn far_6_6177_1_a(.in(far_6_6177_0[0]), .out(far_6_6177_1[0]));    relay_conn far_6_6177_1_b(.in(far_6_6177_0[1]), .out(far_6_6177_1[1]));
    assign layer_6[57] = far_6_6177_1[1] & ~far_6_6177_1[0]; 
    wire [1:0] far_6_6178_0;    relay_conn far_6_6178_0_a(.in(layer_5[576]), .out(far_6_6178_0[0]));    relay_conn far_6_6178_0_b(.in(layer_5[629]), .out(far_6_6178_0[1]));
    assign layer_6[58] = ~far_6_6178_0[0] | (far_6_6178_0[0] & far_6_6178_0[1]); 
    wire [1:0] far_6_6179_0;    relay_conn far_6_6179_0_a(.in(layer_5[388]), .out(far_6_6179_0[0]));    relay_conn far_6_6179_0_b(.in(layer_5[439]), .out(far_6_6179_0[1]));
    assign layer_6[59] = far_6_6179_0[1] & ~far_6_6179_0[0]; 
    wire [1:0] far_6_6180_0;    relay_conn far_6_6180_0_a(.in(layer_5[411]), .out(far_6_6180_0[0]));    relay_conn far_6_6180_0_b(.in(layer_5[315]), .out(far_6_6180_0[1]));
    wire [1:0] far_6_6180_1;    relay_conn far_6_6180_1_a(.in(far_6_6180_0[0]), .out(far_6_6180_1[0]));    relay_conn far_6_6180_1_b(.in(far_6_6180_0[1]), .out(far_6_6180_1[1]));
    wire [1:0] far_6_6180_2;    relay_conn far_6_6180_2_a(.in(far_6_6180_1[0]), .out(far_6_6180_2[0]));    relay_conn far_6_6180_2_b(.in(far_6_6180_1[1]), .out(far_6_6180_2[1]));
    assign layer_6[60] = far_6_6180_2[1]; 
    wire [1:0] far_6_6181_0;    relay_conn far_6_6181_0_a(.in(layer_5[165]), .out(far_6_6181_0[0]));    relay_conn far_6_6181_0_b(.in(layer_5[117]), .out(far_6_6181_0[1]));
    assign layer_6[61] = far_6_6181_0[0] ^ far_6_6181_0[1]; 
    wire [1:0] far_6_6182_0;    relay_conn far_6_6182_0_a(.in(layer_5[152]), .out(far_6_6182_0[0]));    relay_conn far_6_6182_0_b(.in(layer_5[58]), .out(far_6_6182_0[1]));
    wire [1:0] far_6_6182_1;    relay_conn far_6_6182_1_a(.in(far_6_6182_0[0]), .out(far_6_6182_1[0]));    relay_conn far_6_6182_1_b(.in(far_6_6182_0[1]), .out(far_6_6182_1[1]));
    assign layer_6[62] = ~(far_6_6182_1[0] | far_6_6182_1[1]); 
    assign layer_6[63] = layer_5[412]; 
    assign layer_6[64] = ~(layer_5[925] | layer_5[913]); 
    assign layer_6[65] = layer_5[464] | layer_5[474]; 
    wire [1:0] far_6_6186_0;    relay_conn far_6_6186_0_a(.in(layer_5[802]), .out(far_6_6186_0[0]));    relay_conn far_6_6186_0_b(.in(layer_5[748]), .out(far_6_6186_0[1]));
    assign layer_6[66] = ~far_6_6186_0[1] | (far_6_6186_0[0] & far_6_6186_0[1]); 
    wire [1:0] far_6_6187_0;    relay_conn far_6_6187_0_a(.in(layer_5[774]), .out(far_6_6187_0[0]));    relay_conn far_6_6187_0_b(.in(layer_5[845]), .out(far_6_6187_0[1]));
    wire [1:0] far_6_6187_1;    relay_conn far_6_6187_1_a(.in(far_6_6187_0[0]), .out(far_6_6187_1[0]));    relay_conn far_6_6187_1_b(.in(far_6_6187_0[1]), .out(far_6_6187_1[1]));
    assign layer_6[67] = ~far_6_6187_1[0] | (far_6_6187_1[0] & far_6_6187_1[1]); 
    assign layer_6[68] = ~layer_5[19]; 
    assign layer_6[69] = layer_5[777] ^ layer_5[769]; 
    assign layer_6[70] = layer_5[319] & ~layer_5[290]; 
    wire [1:0] far_6_6191_0;    relay_conn far_6_6191_0_a(.in(layer_5[668]), .out(far_6_6191_0[0]));    relay_conn far_6_6191_0_b(.in(layer_5[620]), .out(far_6_6191_0[1]));
    assign layer_6[71] = ~far_6_6191_0[1]; 
    wire [1:0] far_6_6192_0;    relay_conn far_6_6192_0_a(.in(layer_5[406]), .out(far_6_6192_0[0]));    relay_conn far_6_6192_0_b(.in(layer_5[473]), .out(far_6_6192_0[1]));
    wire [1:0] far_6_6192_1;    relay_conn far_6_6192_1_a(.in(far_6_6192_0[0]), .out(far_6_6192_1[0]));    relay_conn far_6_6192_1_b(.in(far_6_6192_0[1]), .out(far_6_6192_1[1]));
    assign layer_6[72] = ~far_6_6192_1[0]; 
    wire [1:0] far_6_6193_0;    relay_conn far_6_6193_0_a(.in(layer_5[487]), .out(far_6_6193_0[0]));    relay_conn far_6_6193_0_b(.in(layer_5[454]), .out(far_6_6193_0[1]));
    assign layer_6[73] = far_6_6193_0[0]; 
    wire [1:0] far_6_6194_0;    relay_conn far_6_6194_0_a(.in(layer_5[224]), .out(far_6_6194_0[0]));    relay_conn far_6_6194_0_b(.in(layer_5[185]), .out(far_6_6194_0[1]));
    assign layer_6[74] = ~far_6_6194_0[1] | (far_6_6194_0[0] & far_6_6194_0[1]); 
    wire [1:0] far_6_6195_0;    relay_conn far_6_6195_0_a(.in(layer_5[759]), .out(far_6_6195_0[0]));    relay_conn far_6_6195_0_b(.in(layer_5[817]), .out(far_6_6195_0[1]));
    assign layer_6[75] = ~(far_6_6195_0[0] | far_6_6195_0[1]); 
    wire [1:0] far_6_6196_0;    relay_conn far_6_6196_0_a(.in(layer_5[795]), .out(far_6_6196_0[0]));    relay_conn far_6_6196_0_b(.in(layer_5[827]), .out(far_6_6196_0[1]));
    assign layer_6[76] = far_6_6196_0[0]; 
    wire [1:0] far_6_6197_0;    relay_conn far_6_6197_0_a(.in(layer_5[735]), .out(far_6_6197_0[0]));    relay_conn far_6_6197_0_b(.in(layer_5[657]), .out(far_6_6197_0[1]));
    wire [1:0] far_6_6197_1;    relay_conn far_6_6197_1_a(.in(far_6_6197_0[0]), .out(far_6_6197_1[0]));    relay_conn far_6_6197_1_b(.in(far_6_6197_0[1]), .out(far_6_6197_1[1]));
    assign layer_6[77] = ~far_6_6197_1[0] | (far_6_6197_1[0] & far_6_6197_1[1]); 
    wire [1:0] far_6_6198_0;    relay_conn far_6_6198_0_a(.in(layer_5[827]), .out(far_6_6198_0[0]));    relay_conn far_6_6198_0_b(.in(layer_5[752]), .out(far_6_6198_0[1]));
    wire [1:0] far_6_6198_1;    relay_conn far_6_6198_1_a(.in(far_6_6198_0[0]), .out(far_6_6198_1[0]));    relay_conn far_6_6198_1_b(.in(far_6_6198_0[1]), .out(far_6_6198_1[1]));
    assign layer_6[78] = far_6_6198_1[0] & ~far_6_6198_1[1]; 
    assign layer_6[79] = layer_5[748] | layer_5[765]; 
    wire [1:0] far_6_6200_0;    relay_conn far_6_6200_0_a(.in(layer_5[743]), .out(far_6_6200_0[0]));    relay_conn far_6_6200_0_b(.in(layer_5[688]), .out(far_6_6200_0[1]));
    assign layer_6[80] = ~far_6_6200_0[1] | (far_6_6200_0[0] & far_6_6200_0[1]); 
    wire [1:0] far_6_6201_0;    relay_conn far_6_6201_0_a(.in(layer_5[729]), .out(far_6_6201_0[0]));    relay_conn far_6_6201_0_b(.in(layer_5[683]), .out(far_6_6201_0[1]));
    assign layer_6[81] = ~(far_6_6201_0[0] | far_6_6201_0[1]); 
    wire [1:0] far_6_6202_0;    relay_conn far_6_6202_0_a(.in(layer_5[328]), .out(far_6_6202_0[0]));    relay_conn far_6_6202_0_b(.in(layer_5[260]), .out(far_6_6202_0[1]));
    wire [1:0] far_6_6202_1;    relay_conn far_6_6202_1_a(.in(far_6_6202_0[0]), .out(far_6_6202_1[0]));    relay_conn far_6_6202_1_b(.in(far_6_6202_0[1]), .out(far_6_6202_1[1]));
    assign layer_6[82] = ~far_6_6202_1[0] | (far_6_6202_1[0] & far_6_6202_1[1]); 
    assign layer_6[83] = layer_5[640] & ~layer_5[616]; 
    assign layer_6[84] = ~layer_5[492]; 
    assign layer_6[85] = layer_5[51] | layer_5[26]; 
    wire [1:0] far_6_6206_0;    relay_conn far_6_6206_0_a(.in(layer_5[837]), .out(far_6_6206_0[0]));    relay_conn far_6_6206_0_b(.in(layer_5[870]), .out(far_6_6206_0[1]));
    assign layer_6[86] = ~far_6_6206_0[1]; 
    wire [1:0] far_6_6207_0;    relay_conn far_6_6207_0_a(.in(layer_5[772]), .out(far_6_6207_0[0]));    relay_conn far_6_6207_0_b(.in(layer_5[729]), .out(far_6_6207_0[1]));
    assign layer_6[87] = ~far_6_6207_0[1] | (far_6_6207_0[0] & far_6_6207_0[1]); 
    wire [1:0] far_6_6208_0;    relay_conn far_6_6208_0_a(.in(layer_5[886]), .out(far_6_6208_0[0]));    relay_conn far_6_6208_0_b(.in(layer_5[939]), .out(far_6_6208_0[1]));
    assign layer_6[88] = far_6_6208_0[1] & ~far_6_6208_0[0]; 
    assign layer_6[89] = ~layer_5[95]; 
    wire [1:0] far_6_6210_0;    relay_conn far_6_6210_0_a(.in(layer_5[457]), .out(far_6_6210_0[0]));    relay_conn far_6_6210_0_b(.in(layer_5[527]), .out(far_6_6210_0[1]));
    wire [1:0] far_6_6210_1;    relay_conn far_6_6210_1_a(.in(far_6_6210_0[0]), .out(far_6_6210_1[0]));    relay_conn far_6_6210_1_b(.in(far_6_6210_0[1]), .out(far_6_6210_1[1]));
    assign layer_6[90] = far_6_6210_1[0] & far_6_6210_1[1]; 
    wire [1:0] far_6_6211_0;    relay_conn far_6_6211_0_a(.in(layer_5[717]), .out(far_6_6211_0[0]));    relay_conn far_6_6211_0_b(.in(layer_5[840]), .out(far_6_6211_0[1]));
    wire [1:0] far_6_6211_1;    relay_conn far_6_6211_1_a(.in(far_6_6211_0[0]), .out(far_6_6211_1[0]));    relay_conn far_6_6211_1_b(.in(far_6_6211_0[1]), .out(far_6_6211_1[1]));
    wire [1:0] far_6_6211_2;    relay_conn far_6_6211_2_a(.in(far_6_6211_1[0]), .out(far_6_6211_2[0]));    relay_conn far_6_6211_2_b(.in(far_6_6211_1[1]), .out(far_6_6211_2[1]));
    assign layer_6[91] = far_6_6211_2[1]; 
    assign layer_6[92] = layer_5[258]; 
    assign layer_6[93] = ~layer_5[108] | (layer_5[127] & layer_5[108]); 
    wire [1:0] far_6_6214_0;    relay_conn far_6_6214_0_a(.in(layer_5[148]), .out(far_6_6214_0[0]));    relay_conn far_6_6214_0_b(.in(layer_5[78]), .out(far_6_6214_0[1]));
    wire [1:0] far_6_6214_1;    relay_conn far_6_6214_1_a(.in(far_6_6214_0[0]), .out(far_6_6214_1[0]));    relay_conn far_6_6214_1_b(.in(far_6_6214_0[1]), .out(far_6_6214_1[1]));
    assign layer_6[94] = far_6_6214_1[0]; 
    assign layer_6[95] = ~layer_5[95]; 
    wire [1:0] far_6_6216_0;    relay_conn far_6_6216_0_a(.in(layer_5[869]), .out(far_6_6216_0[0]));    relay_conn far_6_6216_0_b(.in(layer_5[939]), .out(far_6_6216_0[1]));
    wire [1:0] far_6_6216_1;    relay_conn far_6_6216_1_a(.in(far_6_6216_0[0]), .out(far_6_6216_1[0]));    relay_conn far_6_6216_1_b(.in(far_6_6216_0[1]), .out(far_6_6216_1[1]));
    assign layer_6[96] = far_6_6216_1[0]; 
    assign layer_6[97] = layer_5[791] & ~layer_5[805]; 
    wire [1:0] far_6_6218_0;    relay_conn far_6_6218_0_a(.in(layer_5[791]), .out(far_6_6218_0[0]));    relay_conn far_6_6218_0_b(.in(layer_5[886]), .out(far_6_6218_0[1]));
    wire [1:0] far_6_6218_1;    relay_conn far_6_6218_1_a(.in(far_6_6218_0[0]), .out(far_6_6218_1[0]));    relay_conn far_6_6218_1_b(.in(far_6_6218_0[1]), .out(far_6_6218_1[1]));
    assign layer_6[98] = ~far_6_6218_1[0]; 
    assign layer_6[99] = ~(layer_5[655] ^ layer_5[668]); 
    wire [1:0] far_6_6220_0;    relay_conn far_6_6220_0_a(.in(layer_5[111]), .out(far_6_6220_0[0]));    relay_conn far_6_6220_0_b(.in(layer_5[205]), .out(far_6_6220_0[1]));
    wire [1:0] far_6_6220_1;    relay_conn far_6_6220_1_a(.in(far_6_6220_0[0]), .out(far_6_6220_1[0]));    relay_conn far_6_6220_1_b(.in(far_6_6220_0[1]), .out(far_6_6220_1[1]));
    assign layer_6[100] = far_6_6220_1[1]; 
    wire [1:0] far_6_6221_0;    relay_conn far_6_6221_0_a(.in(layer_5[688]), .out(far_6_6221_0[0]));    relay_conn far_6_6221_0_b(.in(layer_5[629]), .out(far_6_6221_0[1]));
    assign layer_6[101] = far_6_6221_0[0] | far_6_6221_0[1]; 
    wire [1:0] far_6_6222_0;    relay_conn far_6_6222_0_a(.in(layer_5[190]), .out(far_6_6222_0[0]));    relay_conn far_6_6222_0_b(.in(layer_5[247]), .out(far_6_6222_0[1]));
    assign layer_6[102] = far_6_6222_0[1] & ~far_6_6222_0[0]; 
    wire [1:0] far_6_6223_0;    relay_conn far_6_6223_0_a(.in(layer_5[423]), .out(far_6_6223_0[0]));    relay_conn far_6_6223_0_b(.in(layer_5[470]), .out(far_6_6223_0[1]));
    assign layer_6[103] = far_6_6223_0[1] & ~far_6_6223_0[0]; 
    assign layer_6[104] = ~layer_5[333] | (layer_5[333] & layer_5[330]); 
    wire [1:0] far_6_6225_0;    relay_conn far_6_6225_0_a(.in(layer_5[797]), .out(far_6_6225_0[0]));    relay_conn far_6_6225_0_b(.in(layer_5[704]), .out(far_6_6225_0[1]));
    wire [1:0] far_6_6225_1;    relay_conn far_6_6225_1_a(.in(far_6_6225_0[0]), .out(far_6_6225_1[0]));    relay_conn far_6_6225_1_b(.in(far_6_6225_0[1]), .out(far_6_6225_1[1]));
    assign layer_6[105] = ~far_6_6225_1[0]; 
    assign layer_6[106] = layer_5[190] ^ layer_5[194]; 
    wire [1:0] far_6_6227_0;    relay_conn far_6_6227_0_a(.in(layer_5[408]), .out(far_6_6227_0[0]));    relay_conn far_6_6227_0_b(.in(layer_5[477]), .out(far_6_6227_0[1]));
    wire [1:0] far_6_6227_1;    relay_conn far_6_6227_1_a(.in(far_6_6227_0[0]), .out(far_6_6227_1[0]));    relay_conn far_6_6227_1_b(.in(far_6_6227_0[1]), .out(far_6_6227_1[1]));
    assign layer_6[107] = ~(far_6_6227_1[0] | far_6_6227_1[1]); 
    wire [1:0] far_6_6228_0;    relay_conn far_6_6228_0_a(.in(layer_5[952]), .out(far_6_6228_0[0]));    relay_conn far_6_6228_0_b(.in(layer_5[875]), .out(far_6_6228_0[1]));
    wire [1:0] far_6_6228_1;    relay_conn far_6_6228_1_a(.in(far_6_6228_0[0]), .out(far_6_6228_1[0]));    relay_conn far_6_6228_1_b(.in(far_6_6228_0[1]), .out(far_6_6228_1[1]));
    assign layer_6[108] = ~(far_6_6228_1[0] | far_6_6228_1[1]); 
    wire [1:0] far_6_6229_0;    relay_conn far_6_6229_0_a(.in(layer_5[337]), .out(far_6_6229_0[0]));    relay_conn far_6_6229_0_b(.in(layer_5[418]), .out(far_6_6229_0[1]));
    wire [1:0] far_6_6229_1;    relay_conn far_6_6229_1_a(.in(far_6_6229_0[0]), .out(far_6_6229_1[0]));    relay_conn far_6_6229_1_b(.in(far_6_6229_0[1]), .out(far_6_6229_1[1]));
    assign layer_6[109] = ~far_6_6229_1[1]; 
    wire [1:0] far_6_6230_0;    relay_conn far_6_6230_0_a(.in(layer_5[22]), .out(far_6_6230_0[0]));    relay_conn far_6_6230_0_b(.in(layer_5[128]), .out(far_6_6230_0[1]));
    wire [1:0] far_6_6230_1;    relay_conn far_6_6230_1_a(.in(far_6_6230_0[0]), .out(far_6_6230_1[0]));    relay_conn far_6_6230_1_b(.in(far_6_6230_0[1]), .out(far_6_6230_1[1]));
    wire [1:0] far_6_6230_2;    relay_conn far_6_6230_2_a(.in(far_6_6230_1[0]), .out(far_6_6230_2[0]));    relay_conn far_6_6230_2_b(.in(far_6_6230_1[1]), .out(far_6_6230_2[1]));
    assign layer_6[110] = ~far_6_6230_2[0] | (far_6_6230_2[0] & far_6_6230_2[1]); 
    wire [1:0] far_6_6231_0;    relay_conn far_6_6231_0_a(.in(layer_5[746]), .out(far_6_6231_0[0]));    relay_conn far_6_6231_0_b(.in(layer_5[670]), .out(far_6_6231_0[1]));
    wire [1:0] far_6_6231_1;    relay_conn far_6_6231_1_a(.in(far_6_6231_0[0]), .out(far_6_6231_1[0]));    relay_conn far_6_6231_1_b(.in(far_6_6231_0[1]), .out(far_6_6231_1[1]));
    assign layer_6[111] = ~far_6_6231_1[0] | (far_6_6231_1[0] & far_6_6231_1[1]); 
    assign layer_6[112] = layer_5[355] & ~layer_5[376]; 
    wire [1:0] far_6_6233_0;    relay_conn far_6_6233_0_a(.in(layer_5[147]), .out(far_6_6233_0[0]));    relay_conn far_6_6233_0_b(.in(layer_5[45]), .out(far_6_6233_0[1]));
    wire [1:0] far_6_6233_1;    relay_conn far_6_6233_1_a(.in(far_6_6233_0[0]), .out(far_6_6233_1[0]));    relay_conn far_6_6233_1_b(.in(far_6_6233_0[1]), .out(far_6_6233_1[1]));
    wire [1:0] far_6_6233_2;    relay_conn far_6_6233_2_a(.in(far_6_6233_1[0]), .out(far_6_6233_2[0]));    relay_conn far_6_6233_2_b(.in(far_6_6233_1[1]), .out(far_6_6233_2[1]));
    assign layer_6[113] = ~far_6_6233_2[1]; 
    wire [1:0] far_6_6234_0;    relay_conn far_6_6234_0_a(.in(layer_5[513]), .out(far_6_6234_0[0]));    relay_conn far_6_6234_0_b(.in(layer_5[637]), .out(far_6_6234_0[1]));
    wire [1:0] far_6_6234_1;    relay_conn far_6_6234_1_a(.in(far_6_6234_0[0]), .out(far_6_6234_1[0]));    relay_conn far_6_6234_1_b(.in(far_6_6234_0[1]), .out(far_6_6234_1[1]));
    wire [1:0] far_6_6234_2;    relay_conn far_6_6234_2_a(.in(far_6_6234_1[0]), .out(far_6_6234_2[0]));    relay_conn far_6_6234_2_b(.in(far_6_6234_1[1]), .out(far_6_6234_2[1]));
    assign layer_6[114] = far_6_6234_2[0]; 
    wire [1:0] far_6_6235_0;    relay_conn far_6_6235_0_a(.in(layer_5[351]), .out(far_6_6235_0[0]));    relay_conn far_6_6235_0_b(.in(layer_5[415]), .out(far_6_6235_0[1]));
    wire [1:0] far_6_6235_1;    relay_conn far_6_6235_1_a(.in(far_6_6235_0[0]), .out(far_6_6235_1[0]));    relay_conn far_6_6235_1_b(.in(far_6_6235_0[1]), .out(far_6_6235_1[1]));
    assign layer_6[115] = ~(far_6_6235_1[0] ^ far_6_6235_1[1]); 
    wire [1:0] far_6_6236_0;    relay_conn far_6_6236_0_a(.in(layer_5[457]), .out(far_6_6236_0[0]));    relay_conn far_6_6236_0_b(.in(layer_5[415]), .out(far_6_6236_0[1]));
    assign layer_6[116] = far_6_6236_0[1] & ~far_6_6236_0[0]; 
    assign layer_6[117] = layer_5[727]; 
    wire [1:0] far_6_6238_0;    relay_conn far_6_6238_0_a(.in(layer_5[667]), .out(far_6_6238_0[0]));    relay_conn far_6_6238_0_b(.in(layer_5[752]), .out(far_6_6238_0[1]));
    wire [1:0] far_6_6238_1;    relay_conn far_6_6238_1_a(.in(far_6_6238_0[0]), .out(far_6_6238_1[0]));    relay_conn far_6_6238_1_b(.in(far_6_6238_0[1]), .out(far_6_6238_1[1]));
    assign layer_6[118] = ~(far_6_6238_1[0] | far_6_6238_1[1]); 
    wire [1:0] far_6_6239_0;    relay_conn far_6_6239_0_a(.in(layer_5[276]), .out(far_6_6239_0[0]));    relay_conn far_6_6239_0_b(.in(layer_5[375]), .out(far_6_6239_0[1]));
    wire [1:0] far_6_6239_1;    relay_conn far_6_6239_1_a(.in(far_6_6239_0[0]), .out(far_6_6239_1[0]));    relay_conn far_6_6239_1_b(.in(far_6_6239_0[1]), .out(far_6_6239_1[1]));
    wire [1:0] far_6_6239_2;    relay_conn far_6_6239_2_a(.in(far_6_6239_1[0]), .out(far_6_6239_2[0]));    relay_conn far_6_6239_2_b(.in(far_6_6239_1[1]), .out(far_6_6239_2[1]));
    assign layer_6[119] = far_6_6239_2[0] & far_6_6239_2[1]; 
    wire [1:0] far_6_6240_0;    relay_conn far_6_6240_0_a(.in(layer_5[925]), .out(far_6_6240_0[0]));    relay_conn far_6_6240_0_b(.in(layer_5[968]), .out(far_6_6240_0[1]));
    assign layer_6[120] = far_6_6240_0[1] & ~far_6_6240_0[0]; 
    assign layer_6[121] = ~layer_5[780]; 
    wire [1:0] far_6_6242_0;    relay_conn far_6_6242_0_a(.in(layer_5[325]), .out(far_6_6242_0[0]));    relay_conn far_6_6242_0_b(.in(layer_5[359]), .out(far_6_6242_0[1]));
    assign layer_6[122] = ~far_6_6242_0[1]; 
    wire [1:0] far_6_6243_0;    relay_conn far_6_6243_0_a(.in(layer_5[276]), .out(far_6_6243_0[0]));    relay_conn far_6_6243_0_b(.in(layer_5[308]), .out(far_6_6243_0[1]));
    assign layer_6[123] = ~(far_6_6243_0[0] ^ far_6_6243_0[1]); 
    wire [1:0] far_6_6244_0;    relay_conn far_6_6244_0_a(.in(layer_5[432]), .out(far_6_6244_0[0]));    relay_conn far_6_6244_0_b(.in(layer_5[532]), .out(far_6_6244_0[1]));
    wire [1:0] far_6_6244_1;    relay_conn far_6_6244_1_a(.in(far_6_6244_0[0]), .out(far_6_6244_1[0]));    relay_conn far_6_6244_1_b(.in(far_6_6244_0[1]), .out(far_6_6244_1[1]));
    wire [1:0] far_6_6244_2;    relay_conn far_6_6244_2_a(.in(far_6_6244_1[0]), .out(far_6_6244_2[0]));    relay_conn far_6_6244_2_b(.in(far_6_6244_1[1]), .out(far_6_6244_2[1]));
    assign layer_6[124] = far_6_6244_2[0] | far_6_6244_2[1]; 
    assign layer_6[125] = ~layer_5[487] | (layer_5[487] & layer_5[467]); 
    wire [1:0] far_6_6246_0;    relay_conn far_6_6246_0_a(.in(layer_5[690]), .out(far_6_6246_0[0]));    relay_conn far_6_6246_0_b(.in(layer_5[568]), .out(far_6_6246_0[1]));
    wire [1:0] far_6_6246_1;    relay_conn far_6_6246_1_a(.in(far_6_6246_0[0]), .out(far_6_6246_1[0]));    relay_conn far_6_6246_1_b(.in(far_6_6246_0[1]), .out(far_6_6246_1[1]));
    wire [1:0] far_6_6246_2;    relay_conn far_6_6246_2_a(.in(far_6_6246_1[0]), .out(far_6_6246_2[0]));    relay_conn far_6_6246_2_b(.in(far_6_6246_1[1]), .out(far_6_6246_2[1]));
    assign layer_6[126] = far_6_6246_2[0] & ~far_6_6246_2[1]; 
    wire [1:0] far_6_6247_0;    relay_conn far_6_6247_0_a(.in(layer_5[58]), .out(far_6_6247_0[0]));    relay_conn far_6_6247_0_b(.in(layer_5[6]), .out(far_6_6247_0[1]));
    assign layer_6[127] = far_6_6247_0[0] | far_6_6247_0[1]; 
    wire [1:0] far_6_6248_0;    relay_conn far_6_6248_0_a(.in(layer_5[637]), .out(far_6_6248_0[0]));    relay_conn far_6_6248_0_b(.in(layer_5[758]), .out(far_6_6248_0[1]));
    wire [1:0] far_6_6248_1;    relay_conn far_6_6248_1_a(.in(far_6_6248_0[0]), .out(far_6_6248_1[0]));    relay_conn far_6_6248_1_b(.in(far_6_6248_0[1]), .out(far_6_6248_1[1]));
    wire [1:0] far_6_6248_2;    relay_conn far_6_6248_2_a(.in(far_6_6248_1[0]), .out(far_6_6248_2[0]));    relay_conn far_6_6248_2_b(.in(far_6_6248_1[1]), .out(far_6_6248_2[1]));
    assign layer_6[128] = far_6_6248_2[0]; 
    wire [1:0] far_6_6249_0;    relay_conn far_6_6249_0_a(.in(layer_5[860]), .out(far_6_6249_0[0]));    relay_conn far_6_6249_0_b(.in(layer_5[753]), .out(far_6_6249_0[1]));
    wire [1:0] far_6_6249_1;    relay_conn far_6_6249_1_a(.in(far_6_6249_0[0]), .out(far_6_6249_1[0]));    relay_conn far_6_6249_1_b(.in(far_6_6249_0[1]), .out(far_6_6249_1[1]));
    wire [1:0] far_6_6249_2;    relay_conn far_6_6249_2_a(.in(far_6_6249_1[0]), .out(far_6_6249_2[0]));    relay_conn far_6_6249_2_b(.in(far_6_6249_1[1]), .out(far_6_6249_2[1]));
    assign layer_6[129] = ~(far_6_6249_2[0] | far_6_6249_2[1]); 
    assign layer_6[130] = layer_5[110]; 
    wire [1:0] far_6_6251_0;    relay_conn far_6_6251_0_a(.in(layer_5[489]), .out(far_6_6251_0[0]));    relay_conn far_6_6251_0_b(.in(layer_5[613]), .out(far_6_6251_0[1]));
    wire [1:0] far_6_6251_1;    relay_conn far_6_6251_1_a(.in(far_6_6251_0[0]), .out(far_6_6251_1[0]));    relay_conn far_6_6251_1_b(.in(far_6_6251_0[1]), .out(far_6_6251_1[1]));
    wire [1:0] far_6_6251_2;    relay_conn far_6_6251_2_a(.in(far_6_6251_1[0]), .out(far_6_6251_2[0]));    relay_conn far_6_6251_2_b(.in(far_6_6251_1[1]), .out(far_6_6251_2[1]));
    assign layer_6[131] = far_6_6251_2[0] & far_6_6251_2[1]; 
    assign layer_6[132] = layer_5[877] & layer_5[872]; 
    assign layer_6[133] = layer_5[463] & layer_5[494]; 
    assign layer_6[134] = layer_5[400] & ~layer_5[396]; 
    assign layer_6[135] = layer_5[956] | layer_5[949]; 
    wire [1:0] far_6_6256_0;    relay_conn far_6_6256_0_a(.in(layer_5[870]), .out(far_6_6256_0[0]));    relay_conn far_6_6256_0_b(.in(layer_5[952]), .out(far_6_6256_0[1]));
    wire [1:0] far_6_6256_1;    relay_conn far_6_6256_1_a(.in(far_6_6256_0[0]), .out(far_6_6256_1[0]));    relay_conn far_6_6256_1_b(.in(far_6_6256_0[1]), .out(far_6_6256_1[1]));
    assign layer_6[136] = far_6_6256_1[1]; 
    wire [1:0] far_6_6257_0;    relay_conn far_6_6257_0_a(.in(layer_5[996]), .out(far_6_6257_0[0]));    relay_conn far_6_6257_0_b(.in(layer_5[875]), .out(far_6_6257_0[1]));
    wire [1:0] far_6_6257_1;    relay_conn far_6_6257_1_a(.in(far_6_6257_0[0]), .out(far_6_6257_1[0]));    relay_conn far_6_6257_1_b(.in(far_6_6257_0[1]), .out(far_6_6257_1[1]));
    wire [1:0] far_6_6257_2;    relay_conn far_6_6257_2_a(.in(far_6_6257_1[0]), .out(far_6_6257_2[0]));    relay_conn far_6_6257_2_b(.in(far_6_6257_1[1]), .out(far_6_6257_2[1]));
    assign layer_6[137] = far_6_6257_2[0] ^ far_6_6257_2[1]; 
    wire [1:0] far_6_6258_0;    relay_conn far_6_6258_0_a(.in(layer_5[651]), .out(far_6_6258_0[0]));    relay_conn far_6_6258_0_b(.in(layer_5[689]), .out(far_6_6258_0[1]));
    assign layer_6[138] = ~far_6_6258_0[1] | (far_6_6258_0[0] & far_6_6258_0[1]); 
    assign layer_6[139] = ~layer_5[126]; 
    wire [1:0] far_6_6260_0;    relay_conn far_6_6260_0_a(.in(layer_5[980]), .out(far_6_6260_0[0]));    relay_conn far_6_6260_0_b(.in(layer_5[928]), .out(far_6_6260_0[1]));
    assign layer_6[140] = far_6_6260_0[0] | far_6_6260_0[1]; 
    wire [1:0] far_6_6261_0;    relay_conn far_6_6261_0_a(.in(layer_5[80]), .out(far_6_6261_0[0]));    relay_conn far_6_6261_0_b(.in(layer_5[152]), .out(far_6_6261_0[1]));
    wire [1:0] far_6_6261_1;    relay_conn far_6_6261_1_a(.in(far_6_6261_0[0]), .out(far_6_6261_1[0]));    relay_conn far_6_6261_1_b(.in(far_6_6261_0[1]), .out(far_6_6261_1[1]));
    assign layer_6[141] = far_6_6261_1[1]; 
    wire [1:0] far_6_6262_0;    relay_conn far_6_6262_0_a(.in(layer_5[792]), .out(far_6_6262_0[0]));    relay_conn far_6_6262_0_b(.in(layer_5[845]), .out(far_6_6262_0[1]));
    assign layer_6[142] = ~far_6_6262_0[0]; 
    wire [1:0] far_6_6263_0;    relay_conn far_6_6263_0_a(.in(layer_5[612]), .out(far_6_6263_0[0]));    relay_conn far_6_6263_0_b(.in(layer_5[648]), .out(far_6_6263_0[1]));
    assign layer_6[143] = ~far_6_6263_0[0] | (far_6_6263_0[0] & far_6_6263_0[1]); 
    assign layer_6[144] = ~(layer_5[70] & layer_5[47]); 
    wire [1:0] far_6_6265_0;    relay_conn far_6_6265_0_a(.in(layer_5[793]), .out(far_6_6265_0[0]));    relay_conn far_6_6265_0_b(.in(layer_5[740]), .out(far_6_6265_0[1]));
    assign layer_6[145] = far_6_6265_0[1]; 
    assign layer_6[146] = layer_5[1010] & layer_5[996]; 
    wire [1:0] far_6_6267_0;    relay_conn far_6_6267_0_a(.in(layer_5[732]), .out(far_6_6267_0[0]));    relay_conn far_6_6267_0_b(.in(layer_5[688]), .out(far_6_6267_0[1]));
    assign layer_6[147] = far_6_6267_0[0] ^ far_6_6267_0[1]; 
    wire [1:0] far_6_6268_0;    relay_conn far_6_6268_0_a(.in(layer_5[1018]), .out(far_6_6268_0[0]));    relay_conn far_6_6268_0_b(.in(layer_5[972]), .out(far_6_6268_0[1]));
    assign layer_6[148] = far_6_6268_0[0]; 
    wire [1:0] far_6_6269_0;    relay_conn far_6_6269_0_a(.in(layer_5[930]), .out(far_6_6269_0[0]));    relay_conn far_6_6269_0_b(.in(layer_5[839]), .out(far_6_6269_0[1]));
    wire [1:0] far_6_6269_1;    relay_conn far_6_6269_1_a(.in(far_6_6269_0[0]), .out(far_6_6269_1[0]));    relay_conn far_6_6269_1_b(.in(far_6_6269_0[1]), .out(far_6_6269_1[1]));
    assign layer_6[149] = ~(far_6_6269_1[0] & far_6_6269_1[1]); 
    assign layer_6[150] = ~layer_5[77]; 
    wire [1:0] far_6_6271_0;    relay_conn far_6_6271_0_a(.in(layer_5[509]), .out(far_6_6271_0[0]));    relay_conn far_6_6271_0_b(.in(layer_5[627]), .out(far_6_6271_0[1]));
    wire [1:0] far_6_6271_1;    relay_conn far_6_6271_1_a(.in(far_6_6271_0[0]), .out(far_6_6271_1[0]));    relay_conn far_6_6271_1_b(.in(far_6_6271_0[1]), .out(far_6_6271_1[1]));
    wire [1:0] far_6_6271_2;    relay_conn far_6_6271_2_a(.in(far_6_6271_1[0]), .out(far_6_6271_2[0]));    relay_conn far_6_6271_2_b(.in(far_6_6271_1[1]), .out(far_6_6271_2[1]));
    assign layer_6[151] = ~(far_6_6271_2[0] ^ far_6_6271_2[1]); 
    wire [1:0] far_6_6272_0;    relay_conn far_6_6272_0_a(.in(layer_5[818]), .out(far_6_6272_0[0]));    relay_conn far_6_6272_0_b(.in(layer_5[945]), .out(far_6_6272_0[1]));
    wire [1:0] far_6_6272_1;    relay_conn far_6_6272_1_a(.in(far_6_6272_0[0]), .out(far_6_6272_1[0]));    relay_conn far_6_6272_1_b(.in(far_6_6272_0[1]), .out(far_6_6272_1[1]));
    wire [1:0] far_6_6272_2;    relay_conn far_6_6272_2_a(.in(far_6_6272_1[0]), .out(far_6_6272_2[0]));    relay_conn far_6_6272_2_b(.in(far_6_6272_1[1]), .out(far_6_6272_2[1]));
    assign layer_6[152] = far_6_6272_2[1]; 
    wire [1:0] far_6_6273_0;    relay_conn far_6_6273_0_a(.in(layer_5[54]), .out(far_6_6273_0[0]));    relay_conn far_6_6273_0_b(.in(layer_5[115]), .out(far_6_6273_0[1]));
    assign layer_6[153] = ~far_6_6273_0[1]; 
    wire [1:0] far_6_6274_0;    relay_conn far_6_6274_0_a(.in(layer_5[348]), .out(far_6_6274_0[0]));    relay_conn far_6_6274_0_b(.in(layer_5[226]), .out(far_6_6274_0[1]));
    wire [1:0] far_6_6274_1;    relay_conn far_6_6274_1_a(.in(far_6_6274_0[0]), .out(far_6_6274_1[0]));    relay_conn far_6_6274_1_b(.in(far_6_6274_0[1]), .out(far_6_6274_1[1]));
    wire [1:0] far_6_6274_2;    relay_conn far_6_6274_2_a(.in(far_6_6274_1[0]), .out(far_6_6274_2[0]));    relay_conn far_6_6274_2_b(.in(far_6_6274_1[1]), .out(far_6_6274_2[1]));
    assign layer_6[154] = ~(far_6_6274_2[0] ^ far_6_6274_2[1]); 
    wire [1:0] far_6_6275_0;    relay_conn far_6_6275_0_a(.in(layer_5[336]), .out(far_6_6275_0[0]));    relay_conn far_6_6275_0_b(.in(layer_5[230]), .out(far_6_6275_0[1]));
    wire [1:0] far_6_6275_1;    relay_conn far_6_6275_1_a(.in(far_6_6275_0[0]), .out(far_6_6275_1[0]));    relay_conn far_6_6275_1_b(.in(far_6_6275_0[1]), .out(far_6_6275_1[1]));
    wire [1:0] far_6_6275_2;    relay_conn far_6_6275_2_a(.in(far_6_6275_1[0]), .out(far_6_6275_2[0]));    relay_conn far_6_6275_2_b(.in(far_6_6275_1[1]), .out(far_6_6275_2[1]));
    assign layer_6[155] = ~far_6_6275_2[1]; 
    wire [1:0] far_6_6276_0;    relay_conn far_6_6276_0_a(.in(layer_5[984]), .out(far_6_6276_0[0]));    relay_conn far_6_6276_0_b(.in(layer_5[933]), .out(far_6_6276_0[1]));
    assign layer_6[156] = far_6_6276_0[0] & ~far_6_6276_0[1]; 
    wire [1:0] far_6_6277_0;    relay_conn far_6_6277_0_a(.in(layer_5[687]), .out(far_6_6277_0[0]));    relay_conn far_6_6277_0_b(.in(layer_5[584]), .out(far_6_6277_0[1]));
    wire [1:0] far_6_6277_1;    relay_conn far_6_6277_1_a(.in(far_6_6277_0[0]), .out(far_6_6277_1[0]));    relay_conn far_6_6277_1_b(.in(far_6_6277_0[1]), .out(far_6_6277_1[1]));
    wire [1:0] far_6_6277_2;    relay_conn far_6_6277_2_a(.in(far_6_6277_1[0]), .out(far_6_6277_2[0]));    relay_conn far_6_6277_2_b(.in(far_6_6277_1[1]), .out(far_6_6277_2[1]));
    assign layer_6[157] = far_6_6277_2[1] & ~far_6_6277_2[0]; 
    wire [1:0] far_6_6278_0;    relay_conn far_6_6278_0_a(.in(layer_5[798]), .out(far_6_6278_0[0]));    relay_conn far_6_6278_0_b(.in(layer_5[865]), .out(far_6_6278_0[1]));
    wire [1:0] far_6_6278_1;    relay_conn far_6_6278_1_a(.in(far_6_6278_0[0]), .out(far_6_6278_1[0]));    relay_conn far_6_6278_1_b(.in(far_6_6278_0[1]), .out(far_6_6278_1[1]));
    assign layer_6[158] = ~far_6_6278_1[0] | (far_6_6278_1[0] & far_6_6278_1[1]); 
    wire [1:0] far_6_6279_0;    relay_conn far_6_6279_0_a(.in(layer_5[258]), .out(far_6_6279_0[0]));    relay_conn far_6_6279_0_b(.in(layer_5[216]), .out(far_6_6279_0[1]));
    assign layer_6[159] = far_6_6279_0[0] | far_6_6279_0[1]; 
    assign layer_6[160] = layer_5[234]; 
    assign layer_6[161] = layer_5[876] & ~layer_5[871]; 
    assign layer_6[162] = ~(layer_5[958] ^ layer_5[961]); 
    wire [1:0] far_6_6283_0;    relay_conn far_6_6283_0_a(.in(layer_5[657]), .out(far_6_6283_0[0]));    relay_conn far_6_6283_0_b(.in(layer_5[560]), .out(far_6_6283_0[1]));
    wire [1:0] far_6_6283_1;    relay_conn far_6_6283_1_a(.in(far_6_6283_0[0]), .out(far_6_6283_1[0]));    relay_conn far_6_6283_1_b(.in(far_6_6283_0[1]), .out(far_6_6283_1[1]));
    wire [1:0] far_6_6283_2;    relay_conn far_6_6283_2_a(.in(far_6_6283_1[0]), .out(far_6_6283_2[0]));    relay_conn far_6_6283_2_b(.in(far_6_6283_1[1]), .out(far_6_6283_2[1]));
    assign layer_6[163] = far_6_6283_2[0]; 
    wire [1:0] far_6_6284_0;    relay_conn far_6_6284_0_a(.in(layer_5[124]), .out(far_6_6284_0[0]));    relay_conn far_6_6284_0_b(.in(layer_5[222]), .out(far_6_6284_0[1]));
    wire [1:0] far_6_6284_1;    relay_conn far_6_6284_1_a(.in(far_6_6284_0[0]), .out(far_6_6284_1[0]));    relay_conn far_6_6284_1_b(.in(far_6_6284_0[1]), .out(far_6_6284_1[1]));
    wire [1:0] far_6_6284_2;    relay_conn far_6_6284_2_a(.in(far_6_6284_1[0]), .out(far_6_6284_2[0]));    relay_conn far_6_6284_2_b(.in(far_6_6284_1[1]), .out(far_6_6284_2[1]));
    assign layer_6[164] = far_6_6284_2[0] & far_6_6284_2[1]; 
    wire [1:0] far_6_6285_0;    relay_conn far_6_6285_0_a(.in(layer_5[94]), .out(far_6_6285_0[0]));    relay_conn far_6_6285_0_b(.in(layer_5[7]), .out(far_6_6285_0[1]));
    wire [1:0] far_6_6285_1;    relay_conn far_6_6285_1_a(.in(far_6_6285_0[0]), .out(far_6_6285_1[0]));    relay_conn far_6_6285_1_b(.in(far_6_6285_0[1]), .out(far_6_6285_1[1]));
    assign layer_6[165] = far_6_6285_1[1]; 
    wire [1:0] far_6_6286_0;    relay_conn far_6_6286_0_a(.in(layer_5[553]), .out(far_6_6286_0[0]));    relay_conn far_6_6286_0_b(.in(layer_5[667]), .out(far_6_6286_0[1]));
    wire [1:0] far_6_6286_1;    relay_conn far_6_6286_1_a(.in(far_6_6286_0[0]), .out(far_6_6286_1[0]));    relay_conn far_6_6286_1_b(.in(far_6_6286_0[1]), .out(far_6_6286_1[1]));
    wire [1:0] far_6_6286_2;    relay_conn far_6_6286_2_a(.in(far_6_6286_1[0]), .out(far_6_6286_2[0]));    relay_conn far_6_6286_2_b(.in(far_6_6286_1[1]), .out(far_6_6286_2[1]));
    assign layer_6[166] = ~(far_6_6286_2[0] & far_6_6286_2[1]); 
    wire [1:0] far_6_6287_0;    relay_conn far_6_6287_0_a(.in(layer_5[490]), .out(far_6_6287_0[0]));    relay_conn far_6_6287_0_b(.in(layer_5[533]), .out(far_6_6287_0[1]));
    assign layer_6[167] = ~far_6_6287_0[0] | (far_6_6287_0[0] & far_6_6287_0[1]); 
    assign layer_6[168] = layer_5[993]; 
    wire [1:0] far_6_6289_0;    relay_conn far_6_6289_0_a(.in(layer_5[57]), .out(far_6_6289_0[0]));    relay_conn far_6_6289_0_b(.in(layer_5[115]), .out(far_6_6289_0[1]));
    assign layer_6[169] = far_6_6289_0[0] | far_6_6289_0[1]; 
    wire [1:0] far_6_6290_0;    relay_conn far_6_6290_0_a(.in(layer_5[550]), .out(far_6_6290_0[0]));    relay_conn far_6_6290_0_b(.in(layer_5[477]), .out(far_6_6290_0[1]));
    wire [1:0] far_6_6290_1;    relay_conn far_6_6290_1_a(.in(far_6_6290_0[0]), .out(far_6_6290_1[0]));    relay_conn far_6_6290_1_b(.in(far_6_6290_0[1]), .out(far_6_6290_1[1]));
    assign layer_6[170] = ~(far_6_6290_1[0] ^ far_6_6290_1[1]); 
    wire [1:0] far_6_6291_0;    relay_conn far_6_6291_0_a(.in(layer_5[685]), .out(far_6_6291_0[0]));    relay_conn far_6_6291_0_b(.in(layer_5[722]), .out(far_6_6291_0[1]));
    assign layer_6[171] = far_6_6291_0[0] & far_6_6291_0[1]; 
    wire [1:0] far_6_6292_0;    relay_conn far_6_6292_0_a(.in(layer_5[860]), .out(far_6_6292_0[0]));    relay_conn far_6_6292_0_b(.in(layer_5[765]), .out(far_6_6292_0[1]));
    wire [1:0] far_6_6292_1;    relay_conn far_6_6292_1_a(.in(far_6_6292_0[0]), .out(far_6_6292_1[0]));    relay_conn far_6_6292_1_b(.in(far_6_6292_0[1]), .out(far_6_6292_1[1]));
    assign layer_6[172] = ~far_6_6292_1[1]; 
    wire [1:0] far_6_6293_0;    relay_conn far_6_6293_0_a(.in(layer_5[35]), .out(far_6_6293_0[0]));    relay_conn far_6_6293_0_b(.in(layer_5[157]), .out(far_6_6293_0[1]));
    wire [1:0] far_6_6293_1;    relay_conn far_6_6293_1_a(.in(far_6_6293_0[0]), .out(far_6_6293_1[0]));    relay_conn far_6_6293_1_b(.in(far_6_6293_0[1]), .out(far_6_6293_1[1]));
    wire [1:0] far_6_6293_2;    relay_conn far_6_6293_2_a(.in(far_6_6293_1[0]), .out(far_6_6293_2[0]));    relay_conn far_6_6293_2_b(.in(far_6_6293_1[1]), .out(far_6_6293_2[1]));
    assign layer_6[173] = ~far_6_6293_2[1]; 
    wire [1:0] far_6_6294_0;    relay_conn far_6_6294_0_a(.in(layer_5[454]), .out(far_6_6294_0[0]));    relay_conn far_6_6294_0_b(.in(layer_5[352]), .out(far_6_6294_0[1]));
    wire [1:0] far_6_6294_1;    relay_conn far_6_6294_1_a(.in(far_6_6294_0[0]), .out(far_6_6294_1[0]));    relay_conn far_6_6294_1_b(.in(far_6_6294_0[1]), .out(far_6_6294_1[1]));
    wire [1:0] far_6_6294_2;    relay_conn far_6_6294_2_a(.in(far_6_6294_1[0]), .out(far_6_6294_2[0]));    relay_conn far_6_6294_2_b(.in(far_6_6294_1[1]), .out(far_6_6294_2[1]));
    assign layer_6[174] = far_6_6294_2[0] & ~far_6_6294_2[1]; 
    wire [1:0] far_6_6295_0;    relay_conn far_6_6295_0_a(.in(layer_5[716]), .out(far_6_6295_0[0]));    relay_conn far_6_6295_0_b(.in(layer_5[645]), .out(far_6_6295_0[1]));
    wire [1:0] far_6_6295_1;    relay_conn far_6_6295_1_a(.in(far_6_6295_0[0]), .out(far_6_6295_1[0]));    relay_conn far_6_6295_1_b(.in(far_6_6295_0[1]), .out(far_6_6295_1[1]));
    assign layer_6[175] = ~far_6_6295_1[0]; 
    wire [1:0] far_6_6296_0;    relay_conn far_6_6296_0_a(.in(layer_5[521]), .out(far_6_6296_0[0]));    relay_conn far_6_6296_0_b(.in(layer_5[487]), .out(far_6_6296_0[1]));
    assign layer_6[176] = far_6_6296_0[0]; 
    wire [1:0] far_6_6297_0;    relay_conn far_6_6297_0_a(.in(layer_5[63]), .out(far_6_6297_0[0]));    relay_conn far_6_6297_0_b(.in(layer_5[98]), .out(far_6_6297_0[1]));
    assign layer_6[177] = far_6_6297_0[0] & far_6_6297_0[1]; 
    wire [1:0] far_6_6298_0;    relay_conn far_6_6298_0_a(.in(layer_5[233]), .out(far_6_6298_0[0]));    relay_conn far_6_6298_0_b(.in(layer_5[127]), .out(far_6_6298_0[1]));
    wire [1:0] far_6_6298_1;    relay_conn far_6_6298_1_a(.in(far_6_6298_0[0]), .out(far_6_6298_1[0]));    relay_conn far_6_6298_1_b(.in(far_6_6298_0[1]), .out(far_6_6298_1[1]));
    wire [1:0] far_6_6298_2;    relay_conn far_6_6298_2_a(.in(far_6_6298_1[0]), .out(far_6_6298_2[0]));    relay_conn far_6_6298_2_b(.in(far_6_6298_1[1]), .out(far_6_6298_2[1]));
    assign layer_6[178] = ~far_6_6298_2[0] | (far_6_6298_2[0] & far_6_6298_2[1]); 
    wire [1:0] far_6_6299_0;    relay_conn far_6_6299_0_a(.in(layer_5[730]), .out(far_6_6299_0[0]));    relay_conn far_6_6299_0_b(.in(layer_5[816]), .out(far_6_6299_0[1]));
    wire [1:0] far_6_6299_1;    relay_conn far_6_6299_1_a(.in(far_6_6299_0[0]), .out(far_6_6299_1[0]));    relay_conn far_6_6299_1_b(.in(far_6_6299_0[1]), .out(far_6_6299_1[1]));
    assign layer_6[179] = far_6_6299_1[1]; 
    wire [1:0] far_6_6300_0;    relay_conn far_6_6300_0_a(.in(layer_5[845]), .out(far_6_6300_0[0]));    relay_conn far_6_6300_0_b(.in(layer_5[746]), .out(far_6_6300_0[1]));
    wire [1:0] far_6_6300_1;    relay_conn far_6_6300_1_a(.in(far_6_6300_0[0]), .out(far_6_6300_1[0]));    relay_conn far_6_6300_1_b(.in(far_6_6300_0[1]), .out(far_6_6300_1[1]));
    wire [1:0] far_6_6300_2;    relay_conn far_6_6300_2_a(.in(far_6_6300_1[0]), .out(far_6_6300_2[0]));    relay_conn far_6_6300_2_b(.in(far_6_6300_1[1]), .out(far_6_6300_2[1]));
    assign layer_6[180] = far_6_6300_2[1] & ~far_6_6300_2[0]; 
    wire [1:0] far_6_6301_0;    relay_conn far_6_6301_0_a(.in(layer_5[498]), .out(far_6_6301_0[0]));    relay_conn far_6_6301_0_b(.in(layer_5[584]), .out(far_6_6301_0[1]));
    wire [1:0] far_6_6301_1;    relay_conn far_6_6301_1_a(.in(far_6_6301_0[0]), .out(far_6_6301_1[0]));    relay_conn far_6_6301_1_b(.in(far_6_6301_0[1]), .out(far_6_6301_1[1]));
    assign layer_6[181] = far_6_6301_1[1]; 
    assign layer_6[182] = ~layer_5[910]; 
    wire [1:0] far_6_6303_0;    relay_conn far_6_6303_0_a(.in(layer_5[875]), .out(far_6_6303_0[0]));    relay_conn far_6_6303_0_b(.in(layer_5[983]), .out(far_6_6303_0[1]));
    wire [1:0] far_6_6303_1;    relay_conn far_6_6303_1_a(.in(far_6_6303_0[0]), .out(far_6_6303_1[0]));    relay_conn far_6_6303_1_b(.in(far_6_6303_0[1]), .out(far_6_6303_1[1]));
    wire [1:0] far_6_6303_2;    relay_conn far_6_6303_2_a(.in(far_6_6303_1[0]), .out(far_6_6303_2[0]));    relay_conn far_6_6303_2_b(.in(far_6_6303_1[1]), .out(far_6_6303_2[1]));
    assign layer_6[183] = ~far_6_6303_2[1] | (far_6_6303_2[0] & far_6_6303_2[1]); 
    wire [1:0] far_6_6304_0;    relay_conn far_6_6304_0_a(.in(layer_5[773]), .out(far_6_6304_0[0]));    relay_conn far_6_6304_0_b(.in(layer_5[689]), .out(far_6_6304_0[1]));
    wire [1:0] far_6_6304_1;    relay_conn far_6_6304_1_a(.in(far_6_6304_0[0]), .out(far_6_6304_1[0]));    relay_conn far_6_6304_1_b(.in(far_6_6304_0[1]), .out(far_6_6304_1[1]));
    assign layer_6[184] = far_6_6304_1[1] & ~far_6_6304_1[0]; 
    assign layer_6[185] = layer_5[759] & layer_5[728]; 
    assign layer_6[186] = ~(layer_5[152] | layer_5[156]); 
    wire [1:0] far_6_6307_0;    relay_conn far_6_6307_0_a(.in(layer_5[1002]), .out(far_6_6307_0[0]));    relay_conn far_6_6307_0_b(.in(layer_5[922]), .out(far_6_6307_0[1]));
    wire [1:0] far_6_6307_1;    relay_conn far_6_6307_1_a(.in(far_6_6307_0[0]), .out(far_6_6307_1[0]));    relay_conn far_6_6307_1_b(.in(far_6_6307_0[1]), .out(far_6_6307_1[1]));
    assign layer_6[187] = far_6_6307_1[0] | far_6_6307_1[1]; 
    wire [1:0] far_6_6308_0;    relay_conn far_6_6308_0_a(.in(layer_5[51]), .out(far_6_6308_0[0]));    relay_conn far_6_6308_0_b(.in(layer_5[165]), .out(far_6_6308_0[1]));
    wire [1:0] far_6_6308_1;    relay_conn far_6_6308_1_a(.in(far_6_6308_0[0]), .out(far_6_6308_1[0]));    relay_conn far_6_6308_1_b(.in(far_6_6308_0[1]), .out(far_6_6308_1[1]));
    wire [1:0] far_6_6308_2;    relay_conn far_6_6308_2_a(.in(far_6_6308_1[0]), .out(far_6_6308_2[0]));    relay_conn far_6_6308_2_b(.in(far_6_6308_1[1]), .out(far_6_6308_2[1]));
    assign layer_6[188] = ~(far_6_6308_2[0] & far_6_6308_2[1]); 
    wire [1:0] far_6_6309_0;    relay_conn far_6_6309_0_a(.in(layer_5[439]), .out(far_6_6309_0[0]));    relay_conn far_6_6309_0_b(.in(layer_5[507]), .out(far_6_6309_0[1]));
    wire [1:0] far_6_6309_1;    relay_conn far_6_6309_1_a(.in(far_6_6309_0[0]), .out(far_6_6309_1[0]));    relay_conn far_6_6309_1_b(.in(far_6_6309_0[1]), .out(far_6_6309_1[1]));
    assign layer_6[189] = ~far_6_6309_1[1]; 
    wire [1:0] far_6_6310_0;    relay_conn far_6_6310_0_a(.in(layer_5[980]), .out(far_6_6310_0[0]));    relay_conn far_6_6310_0_b(.in(layer_5[887]), .out(far_6_6310_0[1]));
    wire [1:0] far_6_6310_1;    relay_conn far_6_6310_1_a(.in(far_6_6310_0[0]), .out(far_6_6310_1[0]));    relay_conn far_6_6310_1_b(.in(far_6_6310_0[1]), .out(far_6_6310_1[1]));
    assign layer_6[190] = ~far_6_6310_1[0]; 
    assign layer_6[191] = layer_5[1012]; 
    assign layer_6[192] = layer_5[620] & layer_5[636]; 
    assign layer_6[193] = ~(layer_5[942] | layer_5[917]); 
    wire [1:0] far_6_6314_0;    relay_conn far_6_6314_0_a(.in(layer_5[501]), .out(far_6_6314_0[0]));    relay_conn far_6_6314_0_b(.in(layer_5[424]), .out(far_6_6314_0[1]));
    wire [1:0] far_6_6314_1;    relay_conn far_6_6314_1_a(.in(far_6_6314_0[0]), .out(far_6_6314_1[0]));    relay_conn far_6_6314_1_b(.in(far_6_6314_0[1]), .out(far_6_6314_1[1]));
    assign layer_6[194] = far_6_6314_1[1]; 
    wire [1:0] far_6_6315_0;    relay_conn far_6_6315_0_a(.in(layer_5[339]), .out(far_6_6315_0[0]));    relay_conn far_6_6315_0_b(.in(layer_5[253]), .out(far_6_6315_0[1]));
    wire [1:0] far_6_6315_1;    relay_conn far_6_6315_1_a(.in(far_6_6315_0[0]), .out(far_6_6315_1[0]));    relay_conn far_6_6315_1_b(.in(far_6_6315_0[1]), .out(far_6_6315_1[1]));
    assign layer_6[195] = ~far_6_6315_1[0]; 
    wire [1:0] far_6_6316_0;    relay_conn far_6_6316_0_a(.in(layer_5[426]), .out(far_6_6316_0[0]));    relay_conn far_6_6316_0_b(.in(layer_5[473]), .out(far_6_6316_0[1]));
    assign layer_6[196] = far_6_6316_0[0]; 
    wire [1:0] far_6_6317_0;    relay_conn far_6_6317_0_a(.in(layer_5[817]), .out(far_6_6317_0[0]));    relay_conn far_6_6317_0_b(.in(layer_5[885]), .out(far_6_6317_0[1]));
    wire [1:0] far_6_6317_1;    relay_conn far_6_6317_1_a(.in(far_6_6317_0[0]), .out(far_6_6317_1[0]));    relay_conn far_6_6317_1_b(.in(far_6_6317_0[1]), .out(far_6_6317_1[1]));
    assign layer_6[197] = far_6_6317_1[0]; 
    wire [1:0] far_6_6318_0;    relay_conn far_6_6318_0_a(.in(layer_5[501]), .out(far_6_6318_0[0]));    relay_conn far_6_6318_0_b(.in(layer_5[549]), .out(far_6_6318_0[1]));
    assign layer_6[198] = ~(far_6_6318_0[0] & far_6_6318_0[1]); 
    wire [1:0] far_6_6319_0;    relay_conn far_6_6319_0_a(.in(layer_5[542]), .out(far_6_6319_0[0]));    relay_conn far_6_6319_0_b(.in(layer_5[461]), .out(far_6_6319_0[1]));
    wire [1:0] far_6_6319_1;    relay_conn far_6_6319_1_a(.in(far_6_6319_0[0]), .out(far_6_6319_1[0]));    relay_conn far_6_6319_1_b(.in(far_6_6319_0[1]), .out(far_6_6319_1[1]));
    assign layer_6[199] = far_6_6319_1[0]; 
    wire [1:0] far_6_6320_0;    relay_conn far_6_6320_0_a(.in(layer_5[180]), .out(far_6_6320_0[0]));    relay_conn far_6_6320_0_b(.in(layer_5[52]), .out(far_6_6320_0[1]));
    wire [1:0] far_6_6320_1;    relay_conn far_6_6320_1_a(.in(far_6_6320_0[0]), .out(far_6_6320_1[0]));    relay_conn far_6_6320_1_b(.in(far_6_6320_0[1]), .out(far_6_6320_1[1]));
    wire [1:0] far_6_6320_2;    relay_conn far_6_6320_2_a(.in(far_6_6320_1[0]), .out(far_6_6320_2[0]));    relay_conn far_6_6320_2_b(.in(far_6_6320_1[1]), .out(far_6_6320_2[1]));
    wire [1:0] far_6_6320_3;    relay_conn far_6_6320_3_a(.in(far_6_6320_2[0]), .out(far_6_6320_3[0]));    relay_conn far_6_6320_3_b(.in(far_6_6320_2[1]), .out(far_6_6320_3[1]));
    assign layer_6[200] = far_6_6320_3[0] ^ far_6_6320_3[1]; 
    assign layer_6[201] = ~(layer_5[800] ^ layer_5[804]); 
    assign layer_6[202] = ~(layer_5[643] | layer_5[674]); 
    wire [1:0] far_6_6323_0;    relay_conn far_6_6323_0_a(.in(layer_5[135]), .out(far_6_6323_0[0]));    relay_conn far_6_6323_0_b(.in(layer_5[231]), .out(far_6_6323_0[1]));
    wire [1:0] far_6_6323_1;    relay_conn far_6_6323_1_a(.in(far_6_6323_0[0]), .out(far_6_6323_1[0]));    relay_conn far_6_6323_1_b(.in(far_6_6323_0[1]), .out(far_6_6323_1[1]));
    wire [1:0] far_6_6323_2;    relay_conn far_6_6323_2_a(.in(far_6_6323_1[0]), .out(far_6_6323_2[0]));    relay_conn far_6_6323_2_b(.in(far_6_6323_1[1]), .out(far_6_6323_2[1]));
    assign layer_6[203] = far_6_6323_2[0] | far_6_6323_2[1]; 
    wire [1:0] far_6_6324_0;    relay_conn far_6_6324_0_a(.in(layer_5[424]), .out(far_6_6324_0[0]));    relay_conn far_6_6324_0_b(.in(layer_5[378]), .out(far_6_6324_0[1]));
    assign layer_6[204] = ~far_6_6324_0[1] | (far_6_6324_0[0] & far_6_6324_0[1]); 
    wire [1:0] far_6_6325_0;    relay_conn far_6_6325_0_a(.in(layer_5[201]), .out(far_6_6325_0[0]));    relay_conn far_6_6325_0_b(.in(layer_5[296]), .out(far_6_6325_0[1]));
    wire [1:0] far_6_6325_1;    relay_conn far_6_6325_1_a(.in(far_6_6325_0[0]), .out(far_6_6325_1[0]));    relay_conn far_6_6325_1_b(.in(far_6_6325_0[1]), .out(far_6_6325_1[1]));
    assign layer_6[205] = far_6_6325_1[0]; 
    assign layer_6[206] = layer_5[312]; 
    wire [1:0] far_6_6327_0;    relay_conn far_6_6327_0_a(.in(layer_5[953]), .out(far_6_6327_0[0]));    relay_conn far_6_6327_0_b(.in(layer_5[985]), .out(far_6_6327_0[1]));
    assign layer_6[207] = ~(far_6_6327_0[0] & far_6_6327_0[1]); 
    assign layer_6[208] = ~layer_5[159]; 
    assign layer_6[209] = layer_5[79] & ~layer_5[63]; 
    wire [1:0] far_6_6330_0;    relay_conn far_6_6330_0_a(.in(layer_5[424]), .out(far_6_6330_0[0]));    relay_conn far_6_6330_0_b(.in(layer_5[457]), .out(far_6_6330_0[1]));
    assign layer_6[210] = ~(far_6_6330_0[0] | far_6_6330_0[1]); 
    wire [1:0] far_6_6331_0;    relay_conn far_6_6331_0_a(.in(layer_5[92]), .out(far_6_6331_0[0]));    relay_conn far_6_6331_0_b(.in(layer_5[7]), .out(far_6_6331_0[1]));
    wire [1:0] far_6_6331_1;    relay_conn far_6_6331_1_a(.in(far_6_6331_0[0]), .out(far_6_6331_1[0]));    relay_conn far_6_6331_1_b(.in(far_6_6331_0[1]), .out(far_6_6331_1[1]));
    assign layer_6[211] = far_6_6331_1[0] ^ far_6_6331_1[1]; 
    wire [1:0] far_6_6332_0;    relay_conn far_6_6332_0_a(.in(layer_5[26]), .out(far_6_6332_0[0]));    relay_conn far_6_6332_0_b(.in(layer_5[126]), .out(far_6_6332_0[1]));
    wire [1:0] far_6_6332_1;    relay_conn far_6_6332_1_a(.in(far_6_6332_0[0]), .out(far_6_6332_1[0]));    relay_conn far_6_6332_1_b(.in(far_6_6332_0[1]), .out(far_6_6332_1[1]));
    wire [1:0] far_6_6332_2;    relay_conn far_6_6332_2_a(.in(far_6_6332_1[0]), .out(far_6_6332_2[0]));    relay_conn far_6_6332_2_b(.in(far_6_6332_1[1]), .out(far_6_6332_2[1]));
    assign layer_6[212] = far_6_6332_2[1]; 
    wire [1:0] far_6_6333_0;    relay_conn far_6_6333_0_a(.in(layer_5[560]), .out(far_6_6333_0[0]));    relay_conn far_6_6333_0_b(.in(layer_5[613]), .out(far_6_6333_0[1]));
    assign layer_6[213] = ~(far_6_6333_0[0] | far_6_6333_0[1]); 
    wire [1:0] far_6_6334_0;    relay_conn far_6_6334_0_a(.in(layer_5[16]), .out(far_6_6334_0[0]));    relay_conn far_6_6334_0_b(.in(layer_5[127]), .out(far_6_6334_0[1]));
    wire [1:0] far_6_6334_1;    relay_conn far_6_6334_1_a(.in(far_6_6334_0[0]), .out(far_6_6334_1[0]));    relay_conn far_6_6334_1_b(.in(far_6_6334_0[1]), .out(far_6_6334_1[1]));
    wire [1:0] far_6_6334_2;    relay_conn far_6_6334_2_a(.in(far_6_6334_1[0]), .out(far_6_6334_2[0]));    relay_conn far_6_6334_2_b(.in(far_6_6334_1[1]), .out(far_6_6334_2[1]));
    assign layer_6[214] = far_6_6334_2[0]; 
    wire [1:0] far_6_6335_0;    relay_conn far_6_6335_0_a(.in(layer_5[63]), .out(far_6_6335_0[0]));    relay_conn far_6_6335_0_b(.in(layer_5[190]), .out(far_6_6335_0[1]));
    wire [1:0] far_6_6335_1;    relay_conn far_6_6335_1_a(.in(far_6_6335_0[0]), .out(far_6_6335_1[0]));    relay_conn far_6_6335_1_b(.in(far_6_6335_0[1]), .out(far_6_6335_1[1]));
    wire [1:0] far_6_6335_2;    relay_conn far_6_6335_2_a(.in(far_6_6335_1[0]), .out(far_6_6335_2[0]));    relay_conn far_6_6335_2_b(.in(far_6_6335_1[1]), .out(far_6_6335_2[1]));
    assign layer_6[215] = ~far_6_6335_2[1] | (far_6_6335_2[0] & far_6_6335_2[1]); 
    wire [1:0] far_6_6336_0;    relay_conn far_6_6336_0_a(.in(layer_5[136]), .out(far_6_6336_0[0]));    relay_conn far_6_6336_0_b(.in(layer_5[64]), .out(far_6_6336_0[1]));
    wire [1:0] far_6_6336_1;    relay_conn far_6_6336_1_a(.in(far_6_6336_0[0]), .out(far_6_6336_1[0]));    relay_conn far_6_6336_1_b(.in(far_6_6336_0[1]), .out(far_6_6336_1[1]));
    assign layer_6[216] = ~(far_6_6336_1[0] & far_6_6336_1[1]); 
    assign layer_6[217] = ~(layer_5[928] & layer_5[911]); 
    wire [1:0] far_6_6338_0;    relay_conn far_6_6338_0_a(.in(layer_5[773]), .out(far_6_6338_0[0]));    relay_conn far_6_6338_0_b(.in(layer_5[720]), .out(far_6_6338_0[1]));
    assign layer_6[218] = far_6_6338_0[0] & ~far_6_6338_0[1]; 
    wire [1:0] far_6_6339_0;    relay_conn far_6_6339_0_a(.in(layer_5[178]), .out(far_6_6339_0[0]));    relay_conn far_6_6339_0_b(.in(layer_5[86]), .out(far_6_6339_0[1]));
    wire [1:0] far_6_6339_1;    relay_conn far_6_6339_1_a(.in(far_6_6339_0[0]), .out(far_6_6339_1[0]));    relay_conn far_6_6339_1_b(.in(far_6_6339_0[1]), .out(far_6_6339_1[1]));
    assign layer_6[219] = far_6_6339_1[0] & ~far_6_6339_1[1]; 
    assign layer_6[220] = ~(layer_5[179] | layer_5[201]); 
    wire [1:0] far_6_6341_0;    relay_conn far_6_6341_0_a(.in(layer_5[525]), .out(far_6_6341_0[0]));    relay_conn far_6_6341_0_b(.in(layer_5[469]), .out(far_6_6341_0[1]));
    assign layer_6[221] = far_6_6341_0[1] & ~far_6_6341_0[0]; 
    wire [1:0] far_6_6342_0;    relay_conn far_6_6342_0_a(.in(layer_5[663]), .out(far_6_6342_0[0]));    relay_conn far_6_6342_0_b(.in(layer_5[733]), .out(far_6_6342_0[1]));
    wire [1:0] far_6_6342_1;    relay_conn far_6_6342_1_a(.in(far_6_6342_0[0]), .out(far_6_6342_1[0]));    relay_conn far_6_6342_1_b(.in(far_6_6342_0[1]), .out(far_6_6342_1[1]));
    assign layer_6[222] = ~far_6_6342_1[1]; 
    assign layer_6[223] = layer_5[291]; 
    wire [1:0] far_6_6344_0;    relay_conn far_6_6344_0_a(.in(layer_5[222]), .out(far_6_6344_0[0]));    relay_conn far_6_6344_0_b(.in(layer_5[276]), .out(far_6_6344_0[1]));
    assign layer_6[224] = far_6_6344_0[0] & ~far_6_6344_0[1]; 
    assign layer_6[225] = layer_5[791] & ~layer_5[765]; 
    wire [1:0] far_6_6346_0;    relay_conn far_6_6346_0_a(.in(layer_5[20]), .out(far_6_6346_0[0]));    relay_conn far_6_6346_0_b(.in(layer_5[136]), .out(far_6_6346_0[1]));
    wire [1:0] far_6_6346_1;    relay_conn far_6_6346_1_a(.in(far_6_6346_0[0]), .out(far_6_6346_1[0]));    relay_conn far_6_6346_1_b(.in(far_6_6346_0[1]), .out(far_6_6346_1[1]));
    wire [1:0] far_6_6346_2;    relay_conn far_6_6346_2_a(.in(far_6_6346_1[0]), .out(far_6_6346_2[0]));    relay_conn far_6_6346_2_b(.in(far_6_6346_1[1]), .out(far_6_6346_2[1]));
    assign layer_6[226] = ~far_6_6346_2[1]; 
    assign layer_6[227] = ~layer_5[956] | (layer_5[956] & layer_5[958]); 
    wire [1:0] far_6_6348_0;    relay_conn far_6_6348_0_a(.in(layer_5[107]), .out(far_6_6348_0[0]));    relay_conn far_6_6348_0_b(.in(layer_5[161]), .out(far_6_6348_0[1]));
    assign layer_6[228] = far_6_6348_0[1]; 
    wire [1:0] far_6_6349_0;    relay_conn far_6_6349_0_a(.in(layer_5[827]), .out(far_6_6349_0[0]));    relay_conn far_6_6349_0_b(.in(layer_5[891]), .out(far_6_6349_0[1]));
    wire [1:0] far_6_6349_1;    relay_conn far_6_6349_1_a(.in(far_6_6349_0[0]), .out(far_6_6349_1[0]));    relay_conn far_6_6349_1_b(.in(far_6_6349_0[1]), .out(far_6_6349_1[1]));
    assign layer_6[229] = far_6_6349_1[0] & far_6_6349_1[1]; 
    assign layer_6[230] = layer_5[28]; 
    wire [1:0] far_6_6351_0;    relay_conn far_6_6351_0_a(.in(layer_5[939]), .out(far_6_6351_0[0]));    relay_conn far_6_6351_0_b(.in(layer_5[832]), .out(far_6_6351_0[1]));
    wire [1:0] far_6_6351_1;    relay_conn far_6_6351_1_a(.in(far_6_6351_0[0]), .out(far_6_6351_1[0]));    relay_conn far_6_6351_1_b(.in(far_6_6351_0[1]), .out(far_6_6351_1[1]));
    wire [1:0] far_6_6351_2;    relay_conn far_6_6351_2_a(.in(far_6_6351_1[0]), .out(far_6_6351_2[0]));    relay_conn far_6_6351_2_b(.in(far_6_6351_1[1]), .out(far_6_6351_2[1]));
    assign layer_6[231] = ~(far_6_6351_2[0] | far_6_6351_2[1]); 
    assign layer_6[232] = ~(layer_5[773] ^ layer_5[798]); 
    assign layer_6[233] = ~(layer_5[772] ^ layer_5[774]); 
    wire [1:0] far_6_6354_0;    relay_conn far_6_6354_0_a(.in(layer_5[352]), .out(far_6_6354_0[0]));    relay_conn far_6_6354_0_b(.in(layer_5[227]), .out(far_6_6354_0[1]));
    wire [1:0] far_6_6354_1;    relay_conn far_6_6354_1_a(.in(far_6_6354_0[0]), .out(far_6_6354_1[0]));    relay_conn far_6_6354_1_b(.in(far_6_6354_0[1]), .out(far_6_6354_1[1]));
    wire [1:0] far_6_6354_2;    relay_conn far_6_6354_2_a(.in(far_6_6354_1[0]), .out(far_6_6354_2[0]));    relay_conn far_6_6354_2_b(.in(far_6_6354_1[1]), .out(far_6_6354_2[1]));
    assign layer_6[234] = far_6_6354_2[0] & ~far_6_6354_2[1]; 
    assign layer_6[235] = layer_5[427] & layer_5[405]; 
    assign layer_6[236] = ~layer_5[759]; 
    wire [1:0] far_6_6357_0;    relay_conn far_6_6357_0_a(.in(layer_5[83]), .out(far_6_6357_0[0]));    relay_conn far_6_6357_0_b(.in(layer_5[204]), .out(far_6_6357_0[1]));
    wire [1:0] far_6_6357_1;    relay_conn far_6_6357_1_a(.in(far_6_6357_0[0]), .out(far_6_6357_1[0]));    relay_conn far_6_6357_1_b(.in(far_6_6357_0[1]), .out(far_6_6357_1[1]));
    wire [1:0] far_6_6357_2;    relay_conn far_6_6357_2_a(.in(far_6_6357_1[0]), .out(far_6_6357_2[0]));    relay_conn far_6_6357_2_b(.in(far_6_6357_1[1]), .out(far_6_6357_2[1]));
    assign layer_6[237] = ~far_6_6357_2[0]; 
    wire [1:0] far_6_6358_0;    relay_conn far_6_6358_0_a(.in(layer_5[977]), .out(far_6_6358_0[0]));    relay_conn far_6_6358_0_b(.in(layer_5[899]), .out(far_6_6358_0[1]));
    wire [1:0] far_6_6358_1;    relay_conn far_6_6358_1_a(.in(far_6_6358_0[0]), .out(far_6_6358_1[0]));    relay_conn far_6_6358_1_b(.in(far_6_6358_0[1]), .out(far_6_6358_1[1]));
    assign layer_6[238] = far_6_6358_1[0]; 
    wire [1:0] far_6_6359_0;    relay_conn far_6_6359_0_a(.in(layer_5[139]), .out(far_6_6359_0[0]));    relay_conn far_6_6359_0_b(.in(layer_5[54]), .out(far_6_6359_0[1]));
    wire [1:0] far_6_6359_1;    relay_conn far_6_6359_1_a(.in(far_6_6359_0[0]), .out(far_6_6359_1[0]));    relay_conn far_6_6359_1_b(.in(far_6_6359_0[1]), .out(far_6_6359_1[1]));
    assign layer_6[239] = far_6_6359_1[0] | far_6_6359_1[1]; 
    wire [1:0] far_6_6360_0;    relay_conn far_6_6360_0_a(.in(layer_5[870]), .out(far_6_6360_0[0]));    relay_conn far_6_6360_0_b(.in(layer_5[749]), .out(far_6_6360_0[1]));
    wire [1:0] far_6_6360_1;    relay_conn far_6_6360_1_a(.in(far_6_6360_0[0]), .out(far_6_6360_1[0]));    relay_conn far_6_6360_1_b(.in(far_6_6360_0[1]), .out(far_6_6360_1[1]));
    wire [1:0] far_6_6360_2;    relay_conn far_6_6360_2_a(.in(far_6_6360_1[0]), .out(far_6_6360_2[0]));    relay_conn far_6_6360_2_b(.in(far_6_6360_1[1]), .out(far_6_6360_2[1]));
    assign layer_6[240] = far_6_6360_2[1]; 
    wire [1:0] far_6_6361_0;    relay_conn far_6_6361_0_a(.in(layer_5[250]), .out(far_6_6361_0[0]));    relay_conn far_6_6361_0_b(.in(layer_5[374]), .out(far_6_6361_0[1]));
    wire [1:0] far_6_6361_1;    relay_conn far_6_6361_1_a(.in(far_6_6361_0[0]), .out(far_6_6361_1[0]));    relay_conn far_6_6361_1_b(.in(far_6_6361_0[1]), .out(far_6_6361_1[1]));
    wire [1:0] far_6_6361_2;    relay_conn far_6_6361_2_a(.in(far_6_6361_1[0]), .out(far_6_6361_2[0]));    relay_conn far_6_6361_2_b(.in(far_6_6361_1[1]), .out(far_6_6361_2[1]));
    assign layer_6[241] = ~far_6_6361_2[1] | (far_6_6361_2[0] & far_6_6361_2[1]); 
    wire [1:0] far_6_6362_0;    relay_conn far_6_6362_0_a(.in(layer_5[875]), .out(far_6_6362_0[0]));    relay_conn far_6_6362_0_b(.in(layer_5[773]), .out(far_6_6362_0[1]));
    wire [1:0] far_6_6362_1;    relay_conn far_6_6362_1_a(.in(far_6_6362_0[0]), .out(far_6_6362_1[0]));    relay_conn far_6_6362_1_b(.in(far_6_6362_0[1]), .out(far_6_6362_1[1]));
    wire [1:0] far_6_6362_2;    relay_conn far_6_6362_2_a(.in(far_6_6362_1[0]), .out(far_6_6362_2[0]));    relay_conn far_6_6362_2_b(.in(far_6_6362_1[1]), .out(far_6_6362_2[1]));
    assign layer_6[242] = ~far_6_6362_2[1] | (far_6_6362_2[0] & far_6_6362_2[1]); 
    wire [1:0] far_6_6363_0;    relay_conn far_6_6363_0_a(.in(layer_5[901]), .out(far_6_6363_0[0]));    relay_conn far_6_6363_0_b(.in(layer_5[956]), .out(far_6_6363_0[1]));
    assign layer_6[243] = ~far_6_6363_0[1] | (far_6_6363_0[0] & far_6_6363_0[1]); 
    wire [1:0] far_6_6364_0;    relay_conn far_6_6364_0_a(.in(layer_5[85]), .out(far_6_6364_0[0]));    relay_conn far_6_6364_0_b(.in(layer_5[25]), .out(far_6_6364_0[1]));
    assign layer_6[244] = ~far_6_6364_0[1] | (far_6_6364_0[0] & far_6_6364_0[1]); 
    wire [1:0] far_6_6365_0;    relay_conn far_6_6365_0_a(.in(layer_5[743]), .out(far_6_6365_0[0]));    relay_conn far_6_6365_0_b(.in(layer_5[779]), .out(far_6_6365_0[1]));
    assign layer_6[245] = far_6_6365_0[0] ^ far_6_6365_0[1]; 
    wire [1:0] far_6_6366_0;    relay_conn far_6_6366_0_a(.in(layer_5[63]), .out(far_6_6366_0[0]));    relay_conn far_6_6366_0_b(.in(layer_5[121]), .out(far_6_6366_0[1]));
    assign layer_6[246] = ~(far_6_6366_0[0] | far_6_6366_0[1]); 
    wire [1:0] far_6_6367_0;    relay_conn far_6_6367_0_a(.in(layer_5[440]), .out(far_6_6367_0[0]));    relay_conn far_6_6367_0_b(.in(layer_5[533]), .out(far_6_6367_0[1]));
    wire [1:0] far_6_6367_1;    relay_conn far_6_6367_1_a(.in(far_6_6367_0[0]), .out(far_6_6367_1[0]));    relay_conn far_6_6367_1_b(.in(far_6_6367_0[1]), .out(far_6_6367_1[1]));
    assign layer_6[247] = far_6_6367_1[0]; 
    assign layer_6[248] = layer_5[724] ^ layer_5[711]; 
    assign layer_6[249] = ~layer_5[20] | (layer_5[20] & layer_5[40]); 
    wire [1:0] far_6_6370_0;    relay_conn far_6_6370_0_a(.in(layer_5[437]), .out(far_6_6370_0[0]));    relay_conn far_6_6370_0_b(.in(layer_5[330]), .out(far_6_6370_0[1]));
    wire [1:0] far_6_6370_1;    relay_conn far_6_6370_1_a(.in(far_6_6370_0[0]), .out(far_6_6370_1[0]));    relay_conn far_6_6370_1_b(.in(far_6_6370_0[1]), .out(far_6_6370_1[1]));
    wire [1:0] far_6_6370_2;    relay_conn far_6_6370_2_a(.in(far_6_6370_1[0]), .out(far_6_6370_2[0]));    relay_conn far_6_6370_2_b(.in(far_6_6370_1[1]), .out(far_6_6370_2[1]));
    assign layer_6[250] = far_6_6370_2[0] & ~far_6_6370_2[1]; 
    assign layer_6[251] = layer_5[272]; 
    assign layer_6[252] = layer_5[16]; 
    wire [1:0] far_6_6373_0;    relay_conn far_6_6373_0_a(.in(layer_5[569]), .out(far_6_6373_0[0]));    relay_conn far_6_6373_0_b(.in(layer_5[663]), .out(far_6_6373_0[1]));
    wire [1:0] far_6_6373_1;    relay_conn far_6_6373_1_a(.in(far_6_6373_0[0]), .out(far_6_6373_1[0]));    relay_conn far_6_6373_1_b(.in(far_6_6373_0[1]), .out(far_6_6373_1[1]));
    assign layer_6[253] = ~far_6_6373_1[0] | (far_6_6373_1[0] & far_6_6373_1[1]); 
    wire [1:0] far_6_6374_0;    relay_conn far_6_6374_0_a(.in(layer_5[176]), .out(far_6_6374_0[0]));    relay_conn far_6_6374_0_b(.in(layer_5[117]), .out(far_6_6374_0[1]));
    assign layer_6[254] = ~far_6_6374_0[0]; 
    wire [1:0] far_6_6375_0;    relay_conn far_6_6375_0_a(.in(layer_5[963]), .out(far_6_6375_0[0]));    relay_conn far_6_6375_0_b(.in(layer_5[867]), .out(far_6_6375_0[1]));
    wire [1:0] far_6_6375_1;    relay_conn far_6_6375_1_a(.in(far_6_6375_0[0]), .out(far_6_6375_1[0]));    relay_conn far_6_6375_1_b(.in(far_6_6375_0[1]), .out(far_6_6375_1[1]));
    wire [1:0] far_6_6375_2;    relay_conn far_6_6375_2_a(.in(far_6_6375_1[0]), .out(far_6_6375_2[0]));    relay_conn far_6_6375_2_b(.in(far_6_6375_1[1]), .out(far_6_6375_2[1]));
    assign layer_6[255] = ~far_6_6375_2[1] | (far_6_6375_2[0] & far_6_6375_2[1]); 
    wire [1:0] far_6_6376_0;    relay_conn far_6_6376_0_a(.in(layer_5[547]), .out(far_6_6376_0[0]));    relay_conn far_6_6376_0_b(.in(layer_5[435]), .out(far_6_6376_0[1]));
    wire [1:0] far_6_6376_1;    relay_conn far_6_6376_1_a(.in(far_6_6376_0[0]), .out(far_6_6376_1[0]));    relay_conn far_6_6376_1_b(.in(far_6_6376_0[1]), .out(far_6_6376_1[1]));
    wire [1:0] far_6_6376_2;    relay_conn far_6_6376_2_a(.in(far_6_6376_1[0]), .out(far_6_6376_2[0]));    relay_conn far_6_6376_2_b(.in(far_6_6376_1[1]), .out(far_6_6376_2[1]));
    assign layer_6[256] = far_6_6376_2[0] & ~far_6_6376_2[1]; 
    wire [1:0] far_6_6377_0;    relay_conn far_6_6377_0_a(.in(layer_5[983]), .out(far_6_6377_0[0]));    relay_conn far_6_6377_0_b(.in(layer_5[890]), .out(far_6_6377_0[1]));
    wire [1:0] far_6_6377_1;    relay_conn far_6_6377_1_a(.in(far_6_6377_0[0]), .out(far_6_6377_1[0]));    relay_conn far_6_6377_1_b(.in(far_6_6377_0[1]), .out(far_6_6377_1[1]));
    assign layer_6[257] = ~far_6_6377_1[1]; 
    wire [1:0] far_6_6378_0;    relay_conn far_6_6378_0_a(.in(layer_5[862]), .out(far_6_6378_0[0]));    relay_conn far_6_6378_0_b(.in(layer_5[959]), .out(far_6_6378_0[1]));
    wire [1:0] far_6_6378_1;    relay_conn far_6_6378_1_a(.in(far_6_6378_0[0]), .out(far_6_6378_1[0]));    relay_conn far_6_6378_1_b(.in(far_6_6378_0[1]), .out(far_6_6378_1[1]));
    wire [1:0] far_6_6378_2;    relay_conn far_6_6378_2_a(.in(far_6_6378_1[0]), .out(far_6_6378_2[0]));    relay_conn far_6_6378_2_b(.in(far_6_6378_1[1]), .out(far_6_6378_2[1]));
    assign layer_6[258] = far_6_6378_2[0] ^ far_6_6378_2[1]; 
    wire [1:0] far_6_6379_0;    relay_conn far_6_6379_0_a(.in(layer_5[513]), .out(far_6_6379_0[0]));    relay_conn far_6_6379_0_b(.in(layer_5[412]), .out(far_6_6379_0[1]));
    wire [1:0] far_6_6379_1;    relay_conn far_6_6379_1_a(.in(far_6_6379_0[0]), .out(far_6_6379_1[0]));    relay_conn far_6_6379_1_b(.in(far_6_6379_0[1]), .out(far_6_6379_1[1]));
    wire [1:0] far_6_6379_2;    relay_conn far_6_6379_2_a(.in(far_6_6379_1[0]), .out(far_6_6379_2[0]));    relay_conn far_6_6379_2_b(.in(far_6_6379_1[1]), .out(far_6_6379_2[1]));
    assign layer_6[259] = far_6_6379_2[0] ^ far_6_6379_2[1]; 
    wire [1:0] far_6_6380_0;    relay_conn far_6_6380_0_a(.in(layer_5[333]), .out(far_6_6380_0[0]));    relay_conn far_6_6380_0_b(.in(layer_5[452]), .out(far_6_6380_0[1]));
    wire [1:0] far_6_6380_1;    relay_conn far_6_6380_1_a(.in(far_6_6380_0[0]), .out(far_6_6380_1[0]));    relay_conn far_6_6380_1_b(.in(far_6_6380_0[1]), .out(far_6_6380_1[1]));
    wire [1:0] far_6_6380_2;    relay_conn far_6_6380_2_a(.in(far_6_6380_1[0]), .out(far_6_6380_2[0]));    relay_conn far_6_6380_2_b(.in(far_6_6380_1[1]), .out(far_6_6380_2[1]));
    assign layer_6[260] = ~far_6_6380_2[1]; 
    assign layer_6[261] = ~layer_5[706]; 
    wire [1:0] far_6_6382_0;    relay_conn far_6_6382_0_a(.in(layer_5[104]), .out(far_6_6382_0[0]));    relay_conn far_6_6382_0_b(.in(layer_5[159]), .out(far_6_6382_0[1]));
    assign layer_6[262] = ~far_6_6382_0[0]; 
    wire [1:0] far_6_6383_0;    relay_conn far_6_6383_0_a(.in(layer_5[10]), .out(far_6_6383_0[0]));    relay_conn far_6_6383_0_b(.in(layer_5[45]), .out(far_6_6383_0[1]));
    assign layer_6[263] = far_6_6383_0[0] & far_6_6383_0[1]; 
    assign layer_6[264] = layer_5[469] & ~layer_5[480]; 
    wire [1:0] far_6_6385_0;    relay_conn far_6_6385_0_a(.in(layer_5[101]), .out(far_6_6385_0[0]));    relay_conn far_6_6385_0_b(.in(layer_5[69]), .out(far_6_6385_0[1]));
    assign layer_6[265] = far_6_6385_0[0] & far_6_6385_0[1]; 
    assign layer_6[266] = ~layer_5[77] | (layer_5[95] & layer_5[77]); 
    wire [1:0] far_6_6387_0;    relay_conn far_6_6387_0_a(.in(layer_5[169]), .out(far_6_6387_0[0]));    relay_conn far_6_6387_0_b(.in(layer_5[231]), .out(far_6_6387_0[1]));
    assign layer_6[267] = ~far_6_6387_0[0]; 
    assign layer_6[268] = ~layer_5[675] | (layer_5[675] & layer_5[673]); 
    assign layer_6[269] = ~layer_5[54] | (layer_5[83] & layer_5[54]); 
    wire [1:0] far_6_6390_0;    relay_conn far_6_6390_0_a(.in(layer_5[290]), .out(far_6_6390_0[0]));    relay_conn far_6_6390_0_b(.in(layer_5[220]), .out(far_6_6390_0[1]));
    wire [1:0] far_6_6390_1;    relay_conn far_6_6390_1_a(.in(far_6_6390_0[0]), .out(far_6_6390_1[0]));    relay_conn far_6_6390_1_b(.in(far_6_6390_0[1]), .out(far_6_6390_1[1]));
    assign layer_6[270] = far_6_6390_1[0]; 
    wire [1:0] far_6_6391_0;    relay_conn far_6_6391_0_a(.in(layer_5[363]), .out(far_6_6391_0[0]));    relay_conn far_6_6391_0_b(.in(layer_5[430]), .out(far_6_6391_0[1]));
    wire [1:0] far_6_6391_1;    relay_conn far_6_6391_1_a(.in(far_6_6391_0[0]), .out(far_6_6391_1[0]));    relay_conn far_6_6391_1_b(.in(far_6_6391_0[1]), .out(far_6_6391_1[1]));
    assign layer_6[271] = ~far_6_6391_1[0]; 
    wire [1:0] far_6_6392_0;    relay_conn far_6_6392_0_a(.in(layer_5[124]), .out(far_6_6392_0[0]));    relay_conn far_6_6392_0_b(.in(layer_5[90]), .out(far_6_6392_0[1]));
    assign layer_6[272] = far_6_6392_0[1] & ~far_6_6392_0[0]; 
    wire [1:0] far_6_6393_0;    relay_conn far_6_6393_0_a(.in(layer_5[520]), .out(far_6_6393_0[0]));    relay_conn far_6_6393_0_b(.in(layer_5[597]), .out(far_6_6393_0[1]));
    wire [1:0] far_6_6393_1;    relay_conn far_6_6393_1_a(.in(far_6_6393_0[0]), .out(far_6_6393_1[0]));    relay_conn far_6_6393_1_b(.in(far_6_6393_0[1]), .out(far_6_6393_1[1]));
    assign layer_6[273] = far_6_6393_1[0]; 
    wire [1:0] far_6_6394_0;    relay_conn far_6_6394_0_a(.in(layer_5[312]), .out(far_6_6394_0[0]));    relay_conn far_6_6394_0_b(.in(layer_5[351]), .out(far_6_6394_0[1]));
    assign layer_6[274] = ~far_6_6394_0[1] | (far_6_6394_0[0] & far_6_6394_0[1]); 
    wire [1:0] far_6_6395_0;    relay_conn far_6_6395_0_a(.in(layer_5[22]), .out(far_6_6395_0[0]));    relay_conn far_6_6395_0_b(.in(layer_5[83]), .out(far_6_6395_0[1]));
    assign layer_6[275] = ~(far_6_6395_0[0] ^ far_6_6395_0[1]); 
    wire [1:0] far_6_6396_0;    relay_conn far_6_6396_0_a(.in(layer_5[102]), .out(far_6_6396_0[0]));    relay_conn far_6_6396_0_b(.in(layer_5[190]), .out(far_6_6396_0[1]));
    wire [1:0] far_6_6396_1;    relay_conn far_6_6396_1_a(.in(far_6_6396_0[0]), .out(far_6_6396_1[0]));    relay_conn far_6_6396_1_b(.in(far_6_6396_0[1]), .out(far_6_6396_1[1]));
    assign layer_6[276] = ~far_6_6396_1[1] | (far_6_6396_1[0] & far_6_6396_1[1]); 
    wire [1:0] far_6_6397_0;    relay_conn far_6_6397_0_a(.in(layer_5[437]), .out(far_6_6397_0[0]));    relay_conn far_6_6397_0_b(.in(layer_5[473]), .out(far_6_6397_0[1]));
    assign layer_6[277] = far_6_6397_0[0]; 
    wire [1:0] far_6_6398_0;    relay_conn far_6_6398_0_a(.in(layer_5[525]), .out(far_6_6398_0[0]));    relay_conn far_6_6398_0_b(.in(layer_5[584]), .out(far_6_6398_0[1]));
    assign layer_6[278] = far_6_6398_0[0] | far_6_6398_0[1]; 
    wire [1:0] far_6_6399_0;    relay_conn far_6_6399_0_a(.in(layer_5[289]), .out(far_6_6399_0[0]));    relay_conn far_6_6399_0_b(.in(layer_5[363]), .out(far_6_6399_0[1]));
    wire [1:0] far_6_6399_1;    relay_conn far_6_6399_1_a(.in(far_6_6399_0[0]), .out(far_6_6399_1[0]));    relay_conn far_6_6399_1_b(.in(far_6_6399_0[1]), .out(far_6_6399_1[1]));
    assign layer_6[279] = far_6_6399_1[0]; 
    wire [1:0] far_6_6400_0;    relay_conn far_6_6400_0_a(.in(layer_5[714]), .out(far_6_6400_0[0]));    relay_conn far_6_6400_0_b(.in(layer_5[644]), .out(far_6_6400_0[1]));
    wire [1:0] far_6_6400_1;    relay_conn far_6_6400_1_a(.in(far_6_6400_0[0]), .out(far_6_6400_1[0]));    relay_conn far_6_6400_1_b(.in(far_6_6400_0[1]), .out(far_6_6400_1[1]));
    assign layer_6[280] = far_6_6400_1[0] & far_6_6400_1[1]; 
    wire [1:0] far_6_6401_0;    relay_conn far_6_6401_0_a(.in(layer_5[291]), .out(far_6_6401_0[0]));    relay_conn far_6_6401_0_b(.in(layer_5[418]), .out(far_6_6401_0[1]));
    wire [1:0] far_6_6401_1;    relay_conn far_6_6401_1_a(.in(far_6_6401_0[0]), .out(far_6_6401_1[0]));    relay_conn far_6_6401_1_b(.in(far_6_6401_0[1]), .out(far_6_6401_1[1]));
    wire [1:0] far_6_6401_2;    relay_conn far_6_6401_2_a(.in(far_6_6401_1[0]), .out(far_6_6401_2[0]));    relay_conn far_6_6401_2_b(.in(far_6_6401_1[1]), .out(far_6_6401_2[1]));
    assign layer_6[281] = ~far_6_6401_2[0] | (far_6_6401_2[0] & far_6_6401_2[1]); 
    wire [1:0] far_6_6402_0;    relay_conn far_6_6402_0_a(.in(layer_5[777]), .out(far_6_6402_0[0]));    relay_conn far_6_6402_0_b(.in(layer_5[653]), .out(far_6_6402_0[1]));
    wire [1:0] far_6_6402_1;    relay_conn far_6_6402_1_a(.in(far_6_6402_0[0]), .out(far_6_6402_1[0]));    relay_conn far_6_6402_1_b(.in(far_6_6402_0[1]), .out(far_6_6402_1[1]));
    wire [1:0] far_6_6402_2;    relay_conn far_6_6402_2_a(.in(far_6_6402_1[0]), .out(far_6_6402_2[0]));    relay_conn far_6_6402_2_b(.in(far_6_6402_1[1]), .out(far_6_6402_2[1]));
    assign layer_6[282] = ~far_6_6402_2[1] | (far_6_6402_2[0] & far_6_6402_2[1]); 
    wire [1:0] far_6_6403_0;    relay_conn far_6_6403_0_a(.in(layer_5[629]), .out(far_6_6403_0[0]));    relay_conn far_6_6403_0_b(.in(layer_5[741]), .out(far_6_6403_0[1]));
    wire [1:0] far_6_6403_1;    relay_conn far_6_6403_1_a(.in(far_6_6403_0[0]), .out(far_6_6403_1[0]));    relay_conn far_6_6403_1_b(.in(far_6_6403_0[1]), .out(far_6_6403_1[1]));
    wire [1:0] far_6_6403_2;    relay_conn far_6_6403_2_a(.in(far_6_6403_1[0]), .out(far_6_6403_2[0]));    relay_conn far_6_6403_2_b(.in(far_6_6403_1[1]), .out(far_6_6403_2[1]));
    assign layer_6[283] = far_6_6403_2[0] | far_6_6403_2[1]; 
    wire [1:0] far_6_6404_0;    relay_conn far_6_6404_0_a(.in(layer_5[149]), .out(far_6_6404_0[0]));    relay_conn far_6_6404_0_b(.in(layer_5[230]), .out(far_6_6404_0[1]));
    wire [1:0] far_6_6404_1;    relay_conn far_6_6404_1_a(.in(far_6_6404_0[0]), .out(far_6_6404_1[0]));    relay_conn far_6_6404_1_b(.in(far_6_6404_0[1]), .out(far_6_6404_1[1]));
    assign layer_6[284] = far_6_6404_1[1]; 
    wire [1:0] far_6_6405_0;    relay_conn far_6_6405_0_a(.in(layer_5[180]), .out(far_6_6405_0[0]));    relay_conn far_6_6405_0_b(.in(layer_5[219]), .out(far_6_6405_0[1]));
    assign layer_6[285] = ~far_6_6405_0[1]; 
    wire [1:0] far_6_6406_0;    relay_conn far_6_6406_0_a(.in(layer_5[402]), .out(far_6_6406_0[0]));    relay_conn far_6_6406_0_b(.in(layer_5[468]), .out(far_6_6406_0[1]));
    wire [1:0] far_6_6406_1;    relay_conn far_6_6406_1_a(.in(far_6_6406_0[0]), .out(far_6_6406_1[0]));    relay_conn far_6_6406_1_b(.in(far_6_6406_0[1]), .out(far_6_6406_1[1]));
    assign layer_6[286] = far_6_6406_1[1]; 
    assign layer_6[287] = ~(layer_5[95] ^ layer_5[104]); 
    assign layer_6[288] = layer_5[452] & layer_5[469]; 
    wire [1:0] far_6_6409_0;    relay_conn far_6_6409_0_a(.in(layer_5[432]), .out(far_6_6409_0[0]));    relay_conn far_6_6409_0_b(.in(layer_5[494]), .out(far_6_6409_0[1]));
    assign layer_6[289] = far_6_6409_0[0]; 
    wire [1:0] far_6_6410_0;    relay_conn far_6_6410_0_a(.in(layer_5[201]), .out(far_6_6410_0[0]));    relay_conn far_6_6410_0_b(.in(layer_5[236]), .out(far_6_6410_0[1]));
    assign layer_6[290] = far_6_6410_0[1] & ~far_6_6410_0[0]; 
    wire [1:0] far_6_6411_0;    relay_conn far_6_6411_0_a(.in(layer_5[194]), .out(far_6_6411_0[0]));    relay_conn far_6_6411_0_b(.in(layer_5[93]), .out(far_6_6411_0[1]));
    wire [1:0] far_6_6411_1;    relay_conn far_6_6411_1_a(.in(far_6_6411_0[0]), .out(far_6_6411_1[0]));    relay_conn far_6_6411_1_b(.in(far_6_6411_0[1]), .out(far_6_6411_1[1]));
    wire [1:0] far_6_6411_2;    relay_conn far_6_6411_2_a(.in(far_6_6411_1[0]), .out(far_6_6411_2[0]));    relay_conn far_6_6411_2_b(.in(far_6_6411_1[1]), .out(far_6_6411_2[1]));
    assign layer_6[291] = far_6_6411_2[0] ^ far_6_6411_2[1]; 
    wire [1:0] far_6_6412_0;    relay_conn far_6_6412_0_a(.in(layer_5[196]), .out(far_6_6412_0[0]));    relay_conn far_6_6412_0_b(.in(layer_5[92]), .out(far_6_6412_0[1]));
    wire [1:0] far_6_6412_1;    relay_conn far_6_6412_1_a(.in(far_6_6412_0[0]), .out(far_6_6412_1[0]));    relay_conn far_6_6412_1_b(.in(far_6_6412_0[1]), .out(far_6_6412_1[1]));
    wire [1:0] far_6_6412_2;    relay_conn far_6_6412_2_a(.in(far_6_6412_1[0]), .out(far_6_6412_2[0]));    relay_conn far_6_6412_2_b(.in(far_6_6412_1[1]), .out(far_6_6412_2[1]));
    assign layer_6[292] = ~far_6_6412_2[0]; 
    wire [1:0] far_6_6413_0;    relay_conn far_6_6413_0_a(.in(layer_5[341]), .out(far_6_6413_0[0]));    relay_conn far_6_6413_0_b(.in(layer_5[288]), .out(far_6_6413_0[1]));
    assign layer_6[293] = far_6_6413_0[0]; 
    wire [1:0] far_6_6414_0;    relay_conn far_6_6414_0_a(.in(layer_5[584]), .out(far_6_6414_0[0]));    relay_conn far_6_6414_0_b(.in(layer_5[692]), .out(far_6_6414_0[1]));
    wire [1:0] far_6_6414_1;    relay_conn far_6_6414_1_a(.in(far_6_6414_0[0]), .out(far_6_6414_1[0]));    relay_conn far_6_6414_1_b(.in(far_6_6414_0[1]), .out(far_6_6414_1[1]));
    wire [1:0] far_6_6414_2;    relay_conn far_6_6414_2_a(.in(far_6_6414_1[0]), .out(far_6_6414_2[0]));    relay_conn far_6_6414_2_b(.in(far_6_6414_1[1]), .out(far_6_6414_2[1]));
    assign layer_6[294] = far_6_6414_2[0] | far_6_6414_2[1]; 
    wire [1:0] far_6_6415_0;    relay_conn far_6_6415_0_a(.in(layer_5[763]), .out(far_6_6415_0[0]));    relay_conn far_6_6415_0_b(.in(layer_5[860]), .out(far_6_6415_0[1]));
    wire [1:0] far_6_6415_1;    relay_conn far_6_6415_1_a(.in(far_6_6415_0[0]), .out(far_6_6415_1[0]));    relay_conn far_6_6415_1_b(.in(far_6_6415_0[1]), .out(far_6_6415_1[1]));
    wire [1:0] far_6_6415_2;    relay_conn far_6_6415_2_a(.in(far_6_6415_1[0]), .out(far_6_6415_2[0]));    relay_conn far_6_6415_2_b(.in(far_6_6415_1[1]), .out(far_6_6415_2[1]));
    assign layer_6[295] = far_6_6415_2[1]; 
    wire [1:0] far_6_6416_0;    relay_conn far_6_6416_0_a(.in(layer_5[434]), .out(far_6_6416_0[0]));    relay_conn far_6_6416_0_b(.in(layer_5[369]), .out(far_6_6416_0[1]));
    wire [1:0] far_6_6416_1;    relay_conn far_6_6416_1_a(.in(far_6_6416_0[0]), .out(far_6_6416_1[0]));    relay_conn far_6_6416_1_b(.in(far_6_6416_0[1]), .out(far_6_6416_1[1]));
    assign layer_6[296] = far_6_6416_1[0] & ~far_6_6416_1[1]; 
    wire [1:0] far_6_6417_0;    relay_conn far_6_6417_0_a(.in(layer_5[347]), .out(far_6_6417_0[0]));    relay_conn far_6_6417_0_b(.in(layer_5[454]), .out(far_6_6417_0[1]));
    wire [1:0] far_6_6417_1;    relay_conn far_6_6417_1_a(.in(far_6_6417_0[0]), .out(far_6_6417_1[0]));    relay_conn far_6_6417_1_b(.in(far_6_6417_0[1]), .out(far_6_6417_1[1]));
    wire [1:0] far_6_6417_2;    relay_conn far_6_6417_2_a(.in(far_6_6417_1[0]), .out(far_6_6417_2[0]));    relay_conn far_6_6417_2_b(.in(far_6_6417_1[1]), .out(far_6_6417_2[1]));
    assign layer_6[297] = far_6_6417_2[0]; 
    wire [1:0] far_6_6418_0;    relay_conn far_6_6418_0_a(.in(layer_5[636]), .out(far_6_6418_0[0]));    relay_conn far_6_6418_0_b(.in(layer_5[528]), .out(far_6_6418_0[1]));
    wire [1:0] far_6_6418_1;    relay_conn far_6_6418_1_a(.in(far_6_6418_0[0]), .out(far_6_6418_1[0]));    relay_conn far_6_6418_1_b(.in(far_6_6418_0[1]), .out(far_6_6418_1[1]));
    wire [1:0] far_6_6418_2;    relay_conn far_6_6418_2_a(.in(far_6_6418_1[0]), .out(far_6_6418_2[0]));    relay_conn far_6_6418_2_b(.in(far_6_6418_1[1]), .out(far_6_6418_2[1]));
    assign layer_6[298] = ~far_6_6418_2[1]; 
    wire [1:0] far_6_6419_0;    relay_conn far_6_6419_0_a(.in(layer_5[784]), .out(far_6_6419_0[0]));    relay_conn far_6_6419_0_b(.in(layer_5[704]), .out(far_6_6419_0[1]));
    wire [1:0] far_6_6419_1;    relay_conn far_6_6419_1_a(.in(far_6_6419_0[0]), .out(far_6_6419_1[0]));    relay_conn far_6_6419_1_b(.in(far_6_6419_0[1]), .out(far_6_6419_1[1]));
    assign layer_6[299] = far_6_6419_1[1]; 
    wire [1:0] far_6_6420_0;    relay_conn far_6_6420_0_a(.in(layer_5[636]), .out(far_6_6420_0[0]));    relay_conn far_6_6420_0_b(.in(layer_5[706]), .out(far_6_6420_0[1]));
    wire [1:0] far_6_6420_1;    relay_conn far_6_6420_1_a(.in(far_6_6420_0[0]), .out(far_6_6420_1[0]));    relay_conn far_6_6420_1_b(.in(far_6_6420_0[1]), .out(far_6_6420_1[1]));
    assign layer_6[300] = far_6_6420_1[0] ^ far_6_6420_1[1]; 
    wire [1:0] far_6_6421_0;    relay_conn far_6_6421_0_a(.in(layer_5[323]), .out(far_6_6421_0[0]));    relay_conn far_6_6421_0_b(.in(layer_5[258]), .out(far_6_6421_0[1]));
    wire [1:0] far_6_6421_1;    relay_conn far_6_6421_1_a(.in(far_6_6421_0[0]), .out(far_6_6421_1[0]));    relay_conn far_6_6421_1_b(.in(far_6_6421_0[1]), .out(far_6_6421_1[1]));
    assign layer_6[301] = ~far_6_6421_1[0] | (far_6_6421_1[0] & far_6_6421_1[1]); 
    wire [1:0] far_6_6422_0;    relay_conn far_6_6422_0_a(.in(layer_5[952]), .out(far_6_6422_0[0]));    relay_conn far_6_6422_0_b(.in(layer_5[993]), .out(far_6_6422_0[1]));
    assign layer_6[302] = ~(far_6_6422_0[0] ^ far_6_6422_0[1]); 
    wire [1:0] far_6_6423_0;    relay_conn far_6_6423_0_a(.in(layer_5[612]), .out(far_6_6423_0[0]));    relay_conn far_6_6423_0_b(.in(layer_5[710]), .out(far_6_6423_0[1]));
    wire [1:0] far_6_6423_1;    relay_conn far_6_6423_1_a(.in(far_6_6423_0[0]), .out(far_6_6423_1[0]));    relay_conn far_6_6423_1_b(.in(far_6_6423_0[1]), .out(far_6_6423_1[1]));
    wire [1:0] far_6_6423_2;    relay_conn far_6_6423_2_a(.in(far_6_6423_1[0]), .out(far_6_6423_2[0]));    relay_conn far_6_6423_2_b(.in(far_6_6423_1[1]), .out(far_6_6423_2[1]));
    assign layer_6[303] = far_6_6423_2[0]; 
    wire [1:0] far_6_6424_0;    relay_conn far_6_6424_0_a(.in(layer_5[612]), .out(far_6_6424_0[0]));    relay_conn far_6_6424_0_b(.in(layer_5[651]), .out(far_6_6424_0[1]));
    assign layer_6[304] = far_6_6424_0[1]; 
    assign layer_6[305] = layer_5[424] & layer_5[394]; 
    wire [1:0] far_6_6426_0;    relay_conn far_6_6426_0_a(.in(layer_5[440]), .out(far_6_6426_0[0]));    relay_conn far_6_6426_0_b(.in(layer_5[536]), .out(far_6_6426_0[1]));
    wire [1:0] far_6_6426_1;    relay_conn far_6_6426_1_a(.in(far_6_6426_0[0]), .out(far_6_6426_1[0]));    relay_conn far_6_6426_1_b(.in(far_6_6426_0[1]), .out(far_6_6426_1[1]));
    wire [1:0] far_6_6426_2;    relay_conn far_6_6426_2_a(.in(far_6_6426_1[0]), .out(far_6_6426_2[0]));    relay_conn far_6_6426_2_b(.in(far_6_6426_1[1]), .out(far_6_6426_2[1]));
    assign layer_6[306] = ~far_6_6426_2[1]; 
    wire [1:0] far_6_6427_0;    relay_conn far_6_6427_0_a(.in(layer_5[140]), .out(far_6_6427_0[0]));    relay_conn far_6_6427_0_b(.in(layer_5[196]), .out(far_6_6427_0[1]));
    assign layer_6[307] = ~far_6_6427_0[0] | (far_6_6427_0[0] & far_6_6427_0[1]); 
    wire [1:0] far_6_6428_0;    relay_conn far_6_6428_0_a(.in(layer_5[1012]), .out(far_6_6428_0[0]));    relay_conn far_6_6428_0_b(.in(layer_5[967]), .out(far_6_6428_0[1]));
    assign layer_6[308] = ~far_6_6428_0[0]; 
    wire [1:0] far_6_6429_0;    relay_conn far_6_6429_0_a(.in(layer_5[87]), .out(far_6_6429_0[0]));    relay_conn far_6_6429_0_b(.in(layer_5[47]), .out(far_6_6429_0[1]));
    assign layer_6[309] = ~far_6_6429_0[0]; 
    assign layer_6[310] = layer_5[760]; 
    assign layer_6[311] = layer_5[974]; 
    assign layer_6[312] = ~layer_5[770]; 
    assign layer_6[313] = layer_5[1002]; 
    assign layer_6[314] = layer_5[89]; 
    wire [1:0] far_6_6435_0;    relay_conn far_6_6435_0_a(.in(layer_5[678]), .out(far_6_6435_0[0]));    relay_conn far_6_6435_0_b(.in(layer_5[646]), .out(far_6_6435_0[1]));
    assign layer_6[315] = ~far_6_6435_0[0]; 
    wire [1:0] far_6_6436_0;    relay_conn far_6_6436_0_a(.in(layer_5[341]), .out(far_6_6436_0[0]));    relay_conn far_6_6436_0_b(.in(layer_5[375]), .out(far_6_6436_0[1]));
    assign layer_6[316] = ~(far_6_6436_0[0] | far_6_6436_0[1]); 
    wire [1:0] far_6_6437_0;    relay_conn far_6_6437_0_a(.in(layer_5[325]), .out(far_6_6437_0[0]));    relay_conn far_6_6437_0_b(.in(layer_5[424]), .out(far_6_6437_0[1]));
    wire [1:0] far_6_6437_1;    relay_conn far_6_6437_1_a(.in(far_6_6437_0[0]), .out(far_6_6437_1[0]));    relay_conn far_6_6437_1_b(.in(far_6_6437_0[1]), .out(far_6_6437_1[1]));
    wire [1:0] far_6_6437_2;    relay_conn far_6_6437_2_a(.in(far_6_6437_1[0]), .out(far_6_6437_2[0]));    relay_conn far_6_6437_2_b(.in(far_6_6437_1[1]), .out(far_6_6437_2[1]));
    assign layer_6[317] = far_6_6437_2[1] & ~far_6_6437_2[0]; 
    wire [1:0] far_6_6438_0;    relay_conn far_6_6438_0_a(.in(layer_5[921]), .out(far_6_6438_0[0]));    relay_conn far_6_6438_0_b(.in(layer_5[827]), .out(far_6_6438_0[1]));
    wire [1:0] far_6_6438_1;    relay_conn far_6_6438_1_a(.in(far_6_6438_0[0]), .out(far_6_6438_1[0]));    relay_conn far_6_6438_1_b(.in(far_6_6438_0[1]), .out(far_6_6438_1[1]));
    assign layer_6[318] = far_6_6438_1[0] | far_6_6438_1[1]; 
    assign layer_6[319] = layer_5[942]; 
    wire [1:0] far_6_6440_0;    relay_conn far_6_6440_0_a(.in(layer_5[44]), .out(far_6_6440_0[0]));    relay_conn far_6_6440_0_b(.in(layer_5[3]), .out(far_6_6440_0[1]));
    assign layer_6[320] = ~far_6_6440_0[0]; 
    wire [1:0] far_6_6441_0;    relay_conn far_6_6441_0_a(.in(layer_5[3]), .out(far_6_6441_0[0]));    relay_conn far_6_6441_0_b(.in(layer_5[57]), .out(far_6_6441_0[1]));
    assign layer_6[321] = ~(far_6_6441_0[0] & far_6_6441_0[1]); 
    wire [1:0] far_6_6442_0;    relay_conn far_6_6442_0_a(.in(layer_5[571]), .out(far_6_6442_0[0]));    relay_conn far_6_6442_0_b(.in(layer_5[609]), .out(far_6_6442_0[1]));
    assign layer_6[322] = ~(far_6_6442_0[0] | far_6_6442_0[1]); 
    wire [1:0] far_6_6443_0;    relay_conn far_6_6443_0_a(.in(layer_5[319]), .out(far_6_6443_0[0]));    relay_conn far_6_6443_0_b(.in(layer_5[352]), .out(far_6_6443_0[1]));
    assign layer_6[323] = far_6_6443_0[1] & ~far_6_6443_0[0]; 
    assign layer_6[324] = ~layer_5[432] | (layer_5[423] & layer_5[432]); 
    wire [1:0] far_6_6445_0;    relay_conn far_6_6445_0_a(.in(layer_5[360]), .out(far_6_6445_0[0]));    relay_conn far_6_6445_0_b(.in(layer_5[324]), .out(far_6_6445_0[1]));
    assign layer_6[325] = far_6_6445_0[0] & far_6_6445_0[1]; 
    assign layer_6[326] = ~(layer_5[733] & layer_5[764]); 
    wire [1:0] far_6_6447_0;    relay_conn far_6_6447_0_a(.in(layer_5[533]), .out(far_6_6447_0[0]));    relay_conn far_6_6447_0_b(.in(layer_5[602]), .out(far_6_6447_0[1]));
    wire [1:0] far_6_6447_1;    relay_conn far_6_6447_1_a(.in(far_6_6447_0[0]), .out(far_6_6447_1[0]));    relay_conn far_6_6447_1_b(.in(far_6_6447_0[1]), .out(far_6_6447_1[1]));
    assign layer_6[327] = ~far_6_6447_1[1] | (far_6_6447_1[0] & far_6_6447_1[1]); 
    wire [1:0] far_6_6448_0;    relay_conn far_6_6448_0_a(.in(layer_5[733]), .out(far_6_6448_0[0]));    relay_conn far_6_6448_0_b(.in(layer_5[645]), .out(far_6_6448_0[1]));
    wire [1:0] far_6_6448_1;    relay_conn far_6_6448_1_a(.in(far_6_6448_0[0]), .out(far_6_6448_1[0]));    relay_conn far_6_6448_1_b(.in(far_6_6448_0[1]), .out(far_6_6448_1[1]));
    assign layer_6[328] = ~far_6_6448_1[1]; 
    wire [1:0] far_6_6449_0;    relay_conn far_6_6449_0_a(.in(layer_5[399]), .out(far_6_6449_0[0]));    relay_conn far_6_6449_0_b(.in(layer_5[450]), .out(far_6_6449_0[1]));
    assign layer_6[329] = far_6_6449_0[0]; 
    wire [1:0] far_6_6450_0;    relay_conn far_6_6450_0_a(.in(layer_5[282]), .out(far_6_6450_0[0]));    relay_conn far_6_6450_0_b(.in(layer_5[330]), .out(far_6_6450_0[1]));
    assign layer_6[330] = ~(far_6_6450_0[0] | far_6_6450_0[1]); 
    assign layer_6[331] = ~layer_5[129]; 
    wire [1:0] far_6_6452_0;    relay_conn far_6_6452_0_a(.in(layer_5[282]), .out(far_6_6452_0[0]));    relay_conn far_6_6452_0_b(.in(layer_5[409]), .out(far_6_6452_0[1]));
    wire [1:0] far_6_6452_1;    relay_conn far_6_6452_1_a(.in(far_6_6452_0[0]), .out(far_6_6452_1[0]));    relay_conn far_6_6452_1_b(.in(far_6_6452_0[1]), .out(far_6_6452_1[1]));
    wire [1:0] far_6_6452_2;    relay_conn far_6_6452_2_a(.in(far_6_6452_1[0]), .out(far_6_6452_2[0]));    relay_conn far_6_6452_2_b(.in(far_6_6452_1[1]), .out(far_6_6452_2[1]));
    assign layer_6[332] = far_6_6452_2[0] ^ far_6_6452_2[1]; 
    assign layer_6[333] = layer_5[430]; 
    wire [1:0] far_6_6454_0;    relay_conn far_6_6454_0_a(.in(layer_5[520]), .out(far_6_6454_0[0]));    relay_conn far_6_6454_0_b(.in(layer_5[423]), .out(far_6_6454_0[1]));
    wire [1:0] far_6_6454_1;    relay_conn far_6_6454_1_a(.in(far_6_6454_0[0]), .out(far_6_6454_1[0]));    relay_conn far_6_6454_1_b(.in(far_6_6454_0[1]), .out(far_6_6454_1[1]));
    wire [1:0] far_6_6454_2;    relay_conn far_6_6454_2_a(.in(far_6_6454_1[0]), .out(far_6_6454_2[0]));    relay_conn far_6_6454_2_b(.in(far_6_6454_1[1]), .out(far_6_6454_2[1]));
    assign layer_6[334] = far_6_6454_2[1]; 
    assign layer_6[335] = ~layer_5[691]; 
    wire [1:0] far_6_6456_0;    relay_conn far_6_6456_0_a(.in(layer_5[243]), .out(far_6_6456_0[0]));    relay_conn far_6_6456_0_b(.in(layer_5[168]), .out(far_6_6456_0[1]));
    wire [1:0] far_6_6456_1;    relay_conn far_6_6456_1_a(.in(far_6_6456_0[0]), .out(far_6_6456_1[0]));    relay_conn far_6_6456_1_b(.in(far_6_6456_0[1]), .out(far_6_6456_1[1]));
    assign layer_6[336] = far_6_6456_1[0] & far_6_6456_1[1]; 
    wire [1:0] far_6_6457_0;    relay_conn far_6_6457_0_a(.in(layer_5[111]), .out(far_6_6457_0[0]));    relay_conn far_6_6457_0_b(.in(layer_5[165]), .out(far_6_6457_0[1]));
    assign layer_6[337] = far_6_6457_0[0]; 
    wire [1:0] far_6_6458_0;    relay_conn far_6_6458_0_a(.in(layer_5[791]), .out(far_6_6458_0[0]));    relay_conn far_6_6458_0_b(.in(layer_5[886]), .out(far_6_6458_0[1]));
    wire [1:0] far_6_6458_1;    relay_conn far_6_6458_1_a(.in(far_6_6458_0[0]), .out(far_6_6458_1[0]));    relay_conn far_6_6458_1_b(.in(far_6_6458_0[1]), .out(far_6_6458_1[1]));
    assign layer_6[338] = ~far_6_6458_1[1]; 
    wire [1:0] far_6_6459_0;    relay_conn far_6_6459_0_a(.in(layer_5[718]), .out(far_6_6459_0[0]));    relay_conn far_6_6459_0_b(.in(layer_5[759]), .out(far_6_6459_0[1]));
    assign layer_6[339] = ~far_6_6459_0[0]; 
    assign layer_6[340] = layer_5[219] & ~layer_5[221]; 
    wire [1:0] far_6_6461_0;    relay_conn far_6_6461_0_a(.in(layer_5[627]), .out(far_6_6461_0[0]));    relay_conn far_6_6461_0_b(.in(layer_5[706]), .out(far_6_6461_0[1]));
    wire [1:0] far_6_6461_1;    relay_conn far_6_6461_1_a(.in(far_6_6461_0[0]), .out(far_6_6461_1[0]));    relay_conn far_6_6461_1_b(.in(far_6_6461_0[1]), .out(far_6_6461_1[1]));
    assign layer_6[341] = ~far_6_6461_1[0]; 
    wire [1:0] far_6_6462_0;    relay_conn far_6_6462_0_a(.in(layer_5[457]), .out(far_6_6462_0[0]));    relay_conn far_6_6462_0_b(.in(layer_5[366]), .out(far_6_6462_0[1]));
    wire [1:0] far_6_6462_1;    relay_conn far_6_6462_1_a(.in(far_6_6462_0[0]), .out(far_6_6462_1[0]));    relay_conn far_6_6462_1_b(.in(far_6_6462_0[1]), .out(far_6_6462_1[1]));
    assign layer_6[342] = far_6_6462_1[0]; 
    wire [1:0] far_6_6463_0;    relay_conn far_6_6463_0_a(.in(layer_5[53]), .out(far_6_6463_0[0]));    relay_conn far_6_6463_0_b(.in(layer_5[150]), .out(far_6_6463_0[1]));
    wire [1:0] far_6_6463_1;    relay_conn far_6_6463_1_a(.in(far_6_6463_0[0]), .out(far_6_6463_1[0]));    relay_conn far_6_6463_1_b(.in(far_6_6463_0[1]), .out(far_6_6463_1[1]));
    wire [1:0] far_6_6463_2;    relay_conn far_6_6463_2_a(.in(far_6_6463_1[0]), .out(far_6_6463_2[0]));    relay_conn far_6_6463_2_b(.in(far_6_6463_1[1]), .out(far_6_6463_2[1]));
    assign layer_6[343] = ~far_6_6463_2[1]; 
    wire [1:0] far_6_6464_0;    relay_conn far_6_6464_0_a(.in(layer_5[490]), .out(far_6_6464_0[0]));    relay_conn far_6_6464_0_b(.in(layer_5[369]), .out(far_6_6464_0[1]));
    wire [1:0] far_6_6464_1;    relay_conn far_6_6464_1_a(.in(far_6_6464_0[0]), .out(far_6_6464_1[0]));    relay_conn far_6_6464_1_b(.in(far_6_6464_0[1]), .out(far_6_6464_1[1]));
    wire [1:0] far_6_6464_2;    relay_conn far_6_6464_2_a(.in(far_6_6464_1[0]), .out(far_6_6464_2[0]));    relay_conn far_6_6464_2_b(.in(far_6_6464_1[1]), .out(far_6_6464_2[1]));
    assign layer_6[344] = ~far_6_6464_2[1] | (far_6_6464_2[0] & far_6_6464_2[1]); 
    wire [1:0] far_6_6465_0;    relay_conn far_6_6465_0_a(.in(layer_5[687]), .out(far_6_6465_0[0]));    relay_conn far_6_6465_0_b(.in(layer_5[578]), .out(far_6_6465_0[1]));
    wire [1:0] far_6_6465_1;    relay_conn far_6_6465_1_a(.in(far_6_6465_0[0]), .out(far_6_6465_1[0]));    relay_conn far_6_6465_1_b(.in(far_6_6465_0[1]), .out(far_6_6465_1[1]));
    wire [1:0] far_6_6465_2;    relay_conn far_6_6465_2_a(.in(far_6_6465_1[0]), .out(far_6_6465_2[0]));    relay_conn far_6_6465_2_b(.in(far_6_6465_1[1]), .out(far_6_6465_2[1]));
    assign layer_6[345] = ~far_6_6465_2[1] | (far_6_6465_2[0] & far_6_6465_2[1]); 
    wire [1:0] far_6_6466_0;    relay_conn far_6_6466_0_a(.in(layer_5[874]), .out(far_6_6466_0[0]));    relay_conn far_6_6466_0_b(.in(layer_5[959]), .out(far_6_6466_0[1]));
    wire [1:0] far_6_6466_1;    relay_conn far_6_6466_1_a(.in(far_6_6466_0[0]), .out(far_6_6466_1[0]));    relay_conn far_6_6466_1_b(.in(far_6_6466_0[1]), .out(far_6_6466_1[1]));
    assign layer_6[346] = far_6_6466_1[0] & ~far_6_6466_1[1]; 
    wire [1:0] far_6_6467_0;    relay_conn far_6_6467_0_a(.in(layer_5[562]), .out(far_6_6467_0[0]));    relay_conn far_6_6467_0_b(.in(layer_5[670]), .out(far_6_6467_0[1]));
    wire [1:0] far_6_6467_1;    relay_conn far_6_6467_1_a(.in(far_6_6467_0[0]), .out(far_6_6467_1[0]));    relay_conn far_6_6467_1_b(.in(far_6_6467_0[1]), .out(far_6_6467_1[1]));
    wire [1:0] far_6_6467_2;    relay_conn far_6_6467_2_a(.in(far_6_6467_1[0]), .out(far_6_6467_2[0]));    relay_conn far_6_6467_2_b(.in(far_6_6467_1[1]), .out(far_6_6467_2[1]));
    assign layer_6[347] = ~(far_6_6467_2[0] | far_6_6467_2[1]); 
    wire [1:0] far_6_6468_0;    relay_conn far_6_6468_0_a(.in(layer_5[36]), .out(far_6_6468_0[0]));    relay_conn far_6_6468_0_b(.in(layer_5[121]), .out(far_6_6468_0[1]));
    wire [1:0] far_6_6468_1;    relay_conn far_6_6468_1_a(.in(far_6_6468_0[0]), .out(far_6_6468_1[0]));    relay_conn far_6_6468_1_b(.in(far_6_6468_0[1]), .out(far_6_6468_1[1]));
    assign layer_6[348] = ~far_6_6468_1[1]; 
    wire [1:0] far_6_6469_0;    relay_conn far_6_6469_0_a(.in(layer_5[802]), .out(far_6_6469_0[0]));    relay_conn far_6_6469_0_b(.in(layer_5[845]), .out(far_6_6469_0[1]));
    assign layer_6[349] = far_6_6469_0[0] ^ far_6_6469_0[1]; 
    wire [1:0] far_6_6470_0;    relay_conn far_6_6470_0_a(.in(layer_5[70]), .out(far_6_6470_0[0]));    relay_conn far_6_6470_0_b(.in(layer_5[129]), .out(far_6_6470_0[1]));
    assign layer_6[350] = ~(far_6_6470_0[0] & far_6_6470_0[1]); 
    assign layer_6[351] = ~(layer_5[195] ^ layer_5[194]); 
    assign layer_6[352] = layer_5[657] & layer_5[651]; 
    wire [1:0] far_6_6473_0;    relay_conn far_6_6473_0_a(.in(layer_5[533]), .out(far_6_6473_0[0]));    relay_conn far_6_6473_0_b(.in(layer_5[644]), .out(far_6_6473_0[1]));
    wire [1:0] far_6_6473_1;    relay_conn far_6_6473_1_a(.in(far_6_6473_0[0]), .out(far_6_6473_1[0]));    relay_conn far_6_6473_1_b(.in(far_6_6473_0[1]), .out(far_6_6473_1[1]));
    wire [1:0] far_6_6473_2;    relay_conn far_6_6473_2_a(.in(far_6_6473_1[0]), .out(far_6_6473_2[0]));    relay_conn far_6_6473_2_b(.in(far_6_6473_1[1]), .out(far_6_6473_2[1]));
    assign layer_6[353] = far_6_6473_2[1] & ~far_6_6473_2[0]; 
    assign layer_6[354] = layer_5[547] | layer_5[571]; 
    wire [1:0] far_6_6475_0;    relay_conn far_6_6475_0_a(.in(layer_5[977]), .out(far_6_6475_0[0]));    relay_conn far_6_6475_0_b(.in(layer_5[915]), .out(far_6_6475_0[1]));
    assign layer_6[355] = ~far_6_6475_0[1] | (far_6_6475_0[0] & far_6_6475_0[1]); 
    wire [1:0] far_6_6476_0;    relay_conn far_6_6476_0_a(.in(layer_5[746]), .out(far_6_6476_0[0]));    relay_conn far_6_6476_0_b(.in(layer_5[648]), .out(far_6_6476_0[1]));
    wire [1:0] far_6_6476_1;    relay_conn far_6_6476_1_a(.in(far_6_6476_0[0]), .out(far_6_6476_1[0]));    relay_conn far_6_6476_1_b(.in(far_6_6476_0[1]), .out(far_6_6476_1[1]));
    wire [1:0] far_6_6476_2;    relay_conn far_6_6476_2_a(.in(far_6_6476_1[0]), .out(far_6_6476_2[0]));    relay_conn far_6_6476_2_b(.in(far_6_6476_1[1]), .out(far_6_6476_2[1]));
    assign layer_6[356] = far_6_6476_2[0] & far_6_6476_2[1]; 
    assign layer_6[357] = ~(layer_5[36] ^ layer_5[43]); 
    assign layer_6[358] = layer_5[334] & ~layer_5[330]; 
    assign layer_6[359] = layer_5[1] & layer_5[25]; 
    wire [1:0] far_6_6480_0;    relay_conn far_6_6480_0_a(.in(layer_5[689]), .out(far_6_6480_0[0]));    relay_conn far_6_6480_0_b(.in(layer_5[817]), .out(far_6_6480_0[1]));
    wire [1:0] far_6_6480_1;    relay_conn far_6_6480_1_a(.in(far_6_6480_0[0]), .out(far_6_6480_1[0]));    relay_conn far_6_6480_1_b(.in(far_6_6480_0[1]), .out(far_6_6480_1[1]));
    wire [1:0] far_6_6480_2;    relay_conn far_6_6480_2_a(.in(far_6_6480_1[0]), .out(far_6_6480_2[0]));    relay_conn far_6_6480_2_b(.in(far_6_6480_1[1]), .out(far_6_6480_2[1]));
    wire [1:0] far_6_6480_3;    relay_conn far_6_6480_3_a(.in(far_6_6480_2[0]), .out(far_6_6480_3[0]));    relay_conn far_6_6480_3_b(.in(far_6_6480_2[1]), .out(far_6_6480_3[1]));
    assign layer_6[360] = far_6_6480_3[0] & ~far_6_6480_3[1]; 
    wire [1:0] far_6_6481_0;    relay_conn far_6_6481_0_a(.in(layer_5[769]), .out(far_6_6481_0[0]));    relay_conn far_6_6481_0_b(.in(layer_5[837]), .out(far_6_6481_0[1]));
    wire [1:0] far_6_6481_1;    relay_conn far_6_6481_1_a(.in(far_6_6481_0[0]), .out(far_6_6481_1[0]));    relay_conn far_6_6481_1_b(.in(far_6_6481_0[1]), .out(far_6_6481_1[1]));
    assign layer_6[361] = far_6_6481_1[1] & ~far_6_6481_1[0]; 
    wire [1:0] far_6_6482_0;    relay_conn far_6_6482_0_a(.in(layer_5[743]), .out(far_6_6482_0[0]));    relay_conn far_6_6482_0_b(.in(layer_5[685]), .out(far_6_6482_0[1]));
    assign layer_6[362] = far_6_6482_0[1]; 
    wire [1:0] far_6_6483_0;    relay_conn far_6_6483_0_a(.in(layer_5[593]), .out(far_6_6483_0[0]));    relay_conn far_6_6483_0_b(.in(layer_5[543]), .out(far_6_6483_0[1]));
    assign layer_6[363] = ~far_6_6483_0[0]; 
    assign layer_6[364] = ~(layer_5[779] | layer_5[777]); 
    wire [1:0] far_6_6485_0;    relay_conn far_6_6485_0_a(.in(layer_5[685]), .out(far_6_6485_0[0]));    relay_conn far_6_6485_0_b(.in(layer_5[769]), .out(far_6_6485_0[1]));
    wire [1:0] far_6_6485_1;    relay_conn far_6_6485_1_a(.in(far_6_6485_0[0]), .out(far_6_6485_1[0]));    relay_conn far_6_6485_1_b(.in(far_6_6485_0[1]), .out(far_6_6485_1[1]));
    assign layer_6[365] = far_6_6485_1[0] & far_6_6485_1[1]; 
    wire [1:0] far_6_6486_0;    relay_conn far_6_6486_0_a(.in(layer_5[802]), .out(far_6_6486_0[0]));    relay_conn far_6_6486_0_b(.in(layer_5[891]), .out(far_6_6486_0[1]));
    wire [1:0] far_6_6486_1;    relay_conn far_6_6486_1_a(.in(far_6_6486_0[0]), .out(far_6_6486_1[0]));    relay_conn far_6_6486_1_b(.in(far_6_6486_0[1]), .out(far_6_6486_1[1]));
    assign layer_6[366] = far_6_6486_1[0]; 
    wire [1:0] far_6_6487_0;    relay_conn far_6_6487_0_a(.in(layer_5[95]), .out(far_6_6487_0[0]));    relay_conn far_6_6487_0_b(.in(layer_5[6]), .out(far_6_6487_0[1]));
    wire [1:0] far_6_6487_1;    relay_conn far_6_6487_1_a(.in(far_6_6487_0[0]), .out(far_6_6487_1[0]));    relay_conn far_6_6487_1_b(.in(far_6_6487_0[1]), .out(far_6_6487_1[1]));
    assign layer_6[367] = ~far_6_6487_1[0] | (far_6_6487_1[0] & far_6_6487_1[1]); 
    wire [1:0] far_6_6488_0;    relay_conn far_6_6488_0_a(.in(layer_5[666]), .out(far_6_6488_0[0]));    relay_conn far_6_6488_0_b(.in(layer_5[715]), .out(far_6_6488_0[1]));
    assign layer_6[368] = ~(far_6_6488_0[0] ^ far_6_6488_0[1]); 
    wire [1:0] far_6_6489_0;    relay_conn far_6_6489_0_a(.in(layer_5[63]), .out(far_6_6489_0[0]));    relay_conn far_6_6489_0_b(.in(layer_5[186]), .out(far_6_6489_0[1]));
    wire [1:0] far_6_6489_1;    relay_conn far_6_6489_1_a(.in(far_6_6489_0[0]), .out(far_6_6489_1[0]));    relay_conn far_6_6489_1_b(.in(far_6_6489_0[1]), .out(far_6_6489_1[1]));
    wire [1:0] far_6_6489_2;    relay_conn far_6_6489_2_a(.in(far_6_6489_1[0]), .out(far_6_6489_2[0]));    relay_conn far_6_6489_2_b(.in(far_6_6489_1[1]), .out(far_6_6489_2[1]));
    assign layer_6[369] = far_6_6489_2[0] & ~far_6_6489_2[1]; 
    assign layer_6[370] = layer_5[225]; 
    wire [1:0] far_6_6491_0;    relay_conn far_6_6491_0_a(.in(layer_5[224]), .out(far_6_6491_0[0]));    relay_conn far_6_6491_0_b(.in(layer_5[150]), .out(far_6_6491_0[1]));
    wire [1:0] far_6_6491_1;    relay_conn far_6_6491_1_a(.in(far_6_6491_0[0]), .out(far_6_6491_1[0]));    relay_conn far_6_6491_1_b(.in(far_6_6491_0[1]), .out(far_6_6491_1[1]));
    assign layer_6[371] = ~far_6_6491_1[0]; 
    wire [1:0] far_6_6492_0;    relay_conn far_6_6492_0_a(.in(layer_5[613]), .out(far_6_6492_0[0]));    relay_conn far_6_6492_0_b(.in(layer_5[487]), .out(far_6_6492_0[1]));
    wire [1:0] far_6_6492_1;    relay_conn far_6_6492_1_a(.in(far_6_6492_0[0]), .out(far_6_6492_1[0]));    relay_conn far_6_6492_1_b(.in(far_6_6492_0[1]), .out(far_6_6492_1[1]));
    wire [1:0] far_6_6492_2;    relay_conn far_6_6492_2_a(.in(far_6_6492_1[0]), .out(far_6_6492_2[0]));    relay_conn far_6_6492_2_b(.in(far_6_6492_1[1]), .out(far_6_6492_2[1]));
    assign layer_6[372] = ~(far_6_6492_2[0] & far_6_6492_2[1]); 
    wire [1:0] far_6_6493_0;    relay_conn far_6_6493_0_a(.in(layer_5[819]), .out(far_6_6493_0[0]));    relay_conn far_6_6493_0_b(.in(layer_5[865]), .out(far_6_6493_0[1]));
    assign layer_6[373] = ~(far_6_6493_0[0] | far_6_6493_0[1]); 
    wire [1:0] far_6_6494_0;    relay_conn far_6_6494_0_a(.in(layer_5[860]), .out(far_6_6494_0[0]));    relay_conn far_6_6494_0_b(.in(layer_5[779]), .out(far_6_6494_0[1]));
    wire [1:0] far_6_6494_1;    relay_conn far_6_6494_1_a(.in(far_6_6494_0[0]), .out(far_6_6494_1[0]));    relay_conn far_6_6494_1_b(.in(far_6_6494_0[1]), .out(far_6_6494_1[1]));
    assign layer_6[374] = ~(far_6_6494_1[0] | far_6_6494_1[1]); 
    assign layer_6[375] = ~layer_5[862] | (layer_5[862] & layer_5[850]); 
    wire [1:0] far_6_6496_0;    relay_conn far_6_6496_0_a(.in(layer_5[164]), .out(far_6_6496_0[0]));    relay_conn far_6_6496_0_b(.in(layer_5[83]), .out(far_6_6496_0[1]));
    wire [1:0] far_6_6496_1;    relay_conn far_6_6496_1_a(.in(far_6_6496_0[0]), .out(far_6_6496_1[0]));    relay_conn far_6_6496_1_b(.in(far_6_6496_0[1]), .out(far_6_6496_1[1]));
    assign layer_6[376] = far_6_6496_1[1]; 
    wire [1:0] far_6_6497_0;    relay_conn far_6_6497_0_a(.in(layer_5[87]), .out(far_6_6497_0[0]));    relay_conn far_6_6497_0_b(.in(layer_5[52]), .out(far_6_6497_0[1]));
    assign layer_6[377] = ~(far_6_6497_0[0] & far_6_6497_0[1]); 
    assign layer_6[378] = ~(layer_5[122] | layer_5[149]); 
    wire [1:0] far_6_6499_0;    relay_conn far_6_6499_0_a(.in(layer_5[520]), .out(far_6_6499_0[0]));    relay_conn far_6_6499_0_b(.in(layer_5[594]), .out(far_6_6499_0[1]));
    wire [1:0] far_6_6499_1;    relay_conn far_6_6499_1_a(.in(far_6_6499_0[0]), .out(far_6_6499_1[0]));    relay_conn far_6_6499_1_b(.in(far_6_6499_0[1]), .out(far_6_6499_1[1]));
    assign layer_6[379] = far_6_6499_1[1] & ~far_6_6499_1[0]; 
    wire [1:0] far_6_6500_0;    relay_conn far_6_6500_0_a(.in(layer_5[262]), .out(far_6_6500_0[0]));    relay_conn far_6_6500_0_b(.in(layer_5[209]), .out(far_6_6500_0[1]));
    assign layer_6[380] = ~(far_6_6500_0[0] & far_6_6500_0[1]); 
    wire [1:0] far_6_6501_0;    relay_conn far_6_6501_0_a(.in(layer_5[643]), .out(far_6_6501_0[0]));    relay_conn far_6_6501_0_b(.in(layer_5[600]), .out(far_6_6501_0[1]));
    assign layer_6[381] = ~far_6_6501_0[1]; 
    wire [1:0] far_6_6502_0;    relay_conn far_6_6502_0_a(.in(layer_5[60]), .out(far_6_6502_0[0]));    relay_conn far_6_6502_0_b(.in(layer_5[19]), .out(far_6_6502_0[1]));
    assign layer_6[382] = far_6_6502_0[0] & far_6_6502_0[1]; 
    wire [1:0] far_6_6503_0;    relay_conn far_6_6503_0_a(.in(layer_5[348]), .out(far_6_6503_0[0]));    relay_conn far_6_6503_0_b(.in(layer_5[281]), .out(far_6_6503_0[1]));
    wire [1:0] far_6_6503_1;    relay_conn far_6_6503_1_a(.in(far_6_6503_0[0]), .out(far_6_6503_1[0]));    relay_conn far_6_6503_1_b(.in(far_6_6503_0[1]), .out(far_6_6503_1[1]));
    assign layer_6[383] = far_6_6503_1[0]; 
    wire [1:0] far_6_6504_0;    relay_conn far_6_6504_0_a(.in(layer_5[218]), .out(far_6_6504_0[0]));    relay_conn far_6_6504_0_b(.in(layer_5[258]), .out(far_6_6504_0[1]));
    assign layer_6[384] = ~far_6_6504_0[0]; 
    wire [1:0] far_6_6505_0;    relay_conn far_6_6505_0_a(.in(layer_5[258]), .out(far_6_6505_0[0]));    relay_conn far_6_6505_0_b(.in(layer_5[305]), .out(far_6_6505_0[1]));
    assign layer_6[385] = far_6_6505_0[1]; 
    wire [1:0] far_6_6506_0;    relay_conn far_6_6506_0_a(.in(layer_5[1010]), .out(far_6_6506_0[0]));    relay_conn far_6_6506_0_b(.in(layer_5[953]), .out(far_6_6506_0[1]));
    assign layer_6[386] = far_6_6506_0[0]; 
    wire [1:0] far_6_6507_0;    relay_conn far_6_6507_0_a(.in(layer_5[58]), .out(far_6_6507_0[0]));    relay_conn far_6_6507_0_b(.in(layer_5[153]), .out(far_6_6507_0[1]));
    wire [1:0] far_6_6507_1;    relay_conn far_6_6507_1_a(.in(far_6_6507_0[0]), .out(far_6_6507_1[0]));    relay_conn far_6_6507_1_b(.in(far_6_6507_0[1]), .out(far_6_6507_1[1]));
    assign layer_6[387] = ~far_6_6507_1[0]; 
    wire [1:0] far_6_6508_0;    relay_conn far_6_6508_0_a(.in(layer_5[804]), .out(far_6_6508_0[0]));    relay_conn far_6_6508_0_b(.in(layer_5[883]), .out(far_6_6508_0[1]));
    wire [1:0] far_6_6508_1;    relay_conn far_6_6508_1_a(.in(far_6_6508_0[0]), .out(far_6_6508_1[0]));    relay_conn far_6_6508_1_b(.in(far_6_6508_0[1]), .out(far_6_6508_1[1]));
    assign layer_6[388] = far_6_6508_1[1]; 
    assign layer_6[389] = ~layer_5[518] | (layer_5[518] & layer_5[521]); 
    wire [1:0] far_6_6510_0;    relay_conn far_6_6510_0_a(.in(layer_5[215]), .out(far_6_6510_0[0]));    relay_conn far_6_6510_0_b(.in(layer_5[335]), .out(far_6_6510_0[1]));
    wire [1:0] far_6_6510_1;    relay_conn far_6_6510_1_a(.in(far_6_6510_0[0]), .out(far_6_6510_1[0]));    relay_conn far_6_6510_1_b(.in(far_6_6510_0[1]), .out(far_6_6510_1[1]));
    wire [1:0] far_6_6510_2;    relay_conn far_6_6510_2_a(.in(far_6_6510_1[0]), .out(far_6_6510_2[0]));    relay_conn far_6_6510_2_b(.in(far_6_6510_1[1]), .out(far_6_6510_2[1]));
    assign layer_6[390] = ~(far_6_6510_2[0] | far_6_6510_2[1]); 
    wire [1:0] far_6_6511_0;    relay_conn far_6_6511_0_a(.in(layer_5[19]), .out(far_6_6511_0[0]));    relay_conn far_6_6511_0_b(.in(layer_5[52]), .out(far_6_6511_0[1]));
    assign layer_6[391] = far_6_6511_0[0] & far_6_6511_0[1]; 
    wire [1:0] far_6_6512_0;    relay_conn far_6_6512_0_a(.in(layer_5[901]), .out(far_6_6512_0[0]));    relay_conn far_6_6512_0_b(.in(layer_5[847]), .out(far_6_6512_0[1]));
    assign layer_6[392] = ~far_6_6512_0[1]; 
    assign layer_6[393] = layer_5[430]; 
    wire [1:0] far_6_6514_0;    relay_conn far_6_6514_0_a(.in(layer_5[411]), .out(far_6_6514_0[0]));    relay_conn far_6_6514_0_b(.in(layer_5[346]), .out(far_6_6514_0[1]));
    wire [1:0] far_6_6514_1;    relay_conn far_6_6514_1_a(.in(far_6_6514_0[0]), .out(far_6_6514_1[0]));    relay_conn far_6_6514_1_b(.in(far_6_6514_0[1]), .out(far_6_6514_1[1]));
    assign layer_6[394] = far_6_6514_1[1]; 
    wire [1:0] far_6_6515_0;    relay_conn far_6_6515_0_a(.in(layer_5[730]), .out(far_6_6515_0[0]));    relay_conn far_6_6515_0_b(.in(layer_5[651]), .out(far_6_6515_0[1]));
    wire [1:0] far_6_6515_1;    relay_conn far_6_6515_1_a(.in(far_6_6515_0[0]), .out(far_6_6515_1[0]));    relay_conn far_6_6515_1_b(.in(far_6_6515_0[1]), .out(far_6_6515_1[1]));
    assign layer_6[395] = ~far_6_6515_1[1] | (far_6_6515_1[0] & far_6_6515_1[1]); 
    wire [1:0] far_6_6516_0;    relay_conn far_6_6516_0_a(.in(layer_5[736]), .out(far_6_6516_0[0]));    relay_conn far_6_6516_0_b(.in(layer_5[667]), .out(far_6_6516_0[1]));
    wire [1:0] far_6_6516_1;    relay_conn far_6_6516_1_a(.in(far_6_6516_0[0]), .out(far_6_6516_1[0]));    relay_conn far_6_6516_1_b(.in(far_6_6516_0[1]), .out(far_6_6516_1[1]));
    assign layer_6[396] = ~(far_6_6516_1[0] | far_6_6516_1[1]); 
    assign layer_6[397] = layer_5[54] & ~layer_5[58]; 
    wire [1:0] far_6_6518_0;    relay_conn far_6_6518_0_a(.in(layer_5[110]), .out(far_6_6518_0[0]));    relay_conn far_6_6518_0_b(.in(layer_5[205]), .out(far_6_6518_0[1]));
    wire [1:0] far_6_6518_1;    relay_conn far_6_6518_1_a(.in(far_6_6518_0[0]), .out(far_6_6518_1[0]));    relay_conn far_6_6518_1_b(.in(far_6_6518_0[1]), .out(far_6_6518_1[1]));
    assign layer_6[398] = far_6_6518_1[1] & ~far_6_6518_1[0]; 
    wire [1:0] far_6_6519_0;    relay_conn far_6_6519_0_a(.in(layer_5[305]), .out(far_6_6519_0[0]));    relay_conn far_6_6519_0_b(.in(layer_5[394]), .out(far_6_6519_0[1]));
    wire [1:0] far_6_6519_1;    relay_conn far_6_6519_1_a(.in(far_6_6519_0[0]), .out(far_6_6519_1[0]));    relay_conn far_6_6519_1_b(.in(far_6_6519_0[1]), .out(far_6_6519_1[1]));
    assign layer_6[399] = ~(far_6_6519_1[0] & far_6_6519_1[1]); 
    wire [1:0] far_6_6520_0;    relay_conn far_6_6520_0_a(.in(layer_5[471]), .out(far_6_6520_0[0]));    relay_conn far_6_6520_0_b(.in(layer_5[512]), .out(far_6_6520_0[1]));
    assign layer_6[400] = far_6_6520_0[1] & ~far_6_6520_0[0]; 
    wire [1:0] far_6_6521_0;    relay_conn far_6_6521_0_a(.in(layer_5[860]), .out(far_6_6521_0[0]));    relay_conn far_6_6521_0_b(.in(layer_5[761]), .out(far_6_6521_0[1]));
    wire [1:0] far_6_6521_1;    relay_conn far_6_6521_1_a(.in(far_6_6521_0[0]), .out(far_6_6521_1[0]));    relay_conn far_6_6521_1_b(.in(far_6_6521_0[1]), .out(far_6_6521_1[1]));
    wire [1:0] far_6_6521_2;    relay_conn far_6_6521_2_a(.in(far_6_6521_1[0]), .out(far_6_6521_2[0]));    relay_conn far_6_6521_2_b(.in(far_6_6521_1[1]), .out(far_6_6521_2[1]));
    assign layer_6[401] = far_6_6521_2[1] & ~far_6_6521_2[0]; 
    wire [1:0] far_6_6522_0;    relay_conn far_6_6522_0_a(.in(layer_5[596]), .out(far_6_6522_0[0]));    relay_conn far_6_6522_0_b(.in(layer_5[640]), .out(far_6_6522_0[1]));
    assign layer_6[402] = far_6_6522_0[0] & ~far_6_6522_0[1]; 
    wire [1:0] far_6_6523_0;    relay_conn far_6_6523_0_a(.in(layer_5[231]), .out(far_6_6523_0[0]));    relay_conn far_6_6523_0_b(.in(layer_5[120]), .out(far_6_6523_0[1]));
    wire [1:0] far_6_6523_1;    relay_conn far_6_6523_1_a(.in(far_6_6523_0[0]), .out(far_6_6523_1[0]));    relay_conn far_6_6523_1_b(.in(far_6_6523_0[1]), .out(far_6_6523_1[1]));
    wire [1:0] far_6_6523_2;    relay_conn far_6_6523_2_a(.in(far_6_6523_1[0]), .out(far_6_6523_2[0]));    relay_conn far_6_6523_2_b(.in(far_6_6523_1[1]), .out(far_6_6523_2[1]));
    assign layer_6[403] = ~(far_6_6523_2[0] ^ far_6_6523_2[1]); 
    wire [1:0] far_6_6524_0;    relay_conn far_6_6524_0_a(.in(layer_5[432]), .out(far_6_6524_0[0]));    relay_conn far_6_6524_0_b(.in(layer_5[502]), .out(far_6_6524_0[1]));
    wire [1:0] far_6_6524_1;    relay_conn far_6_6524_1_a(.in(far_6_6524_0[0]), .out(far_6_6524_1[0]));    relay_conn far_6_6524_1_b(.in(far_6_6524_0[1]), .out(far_6_6524_1[1]));
    assign layer_6[404] = far_6_6524_1[1]; 
    assign layer_6[405] = layer_5[975]; 
    wire [1:0] far_6_6526_0;    relay_conn far_6_6526_0_a(.in(layer_5[788]), .out(far_6_6526_0[0]));    relay_conn far_6_6526_0_b(.in(layer_5[860]), .out(far_6_6526_0[1]));
    wire [1:0] far_6_6526_1;    relay_conn far_6_6526_1_a(.in(far_6_6526_0[0]), .out(far_6_6526_1[0]));    relay_conn far_6_6526_1_b(.in(far_6_6526_0[1]), .out(far_6_6526_1[1]));
    assign layer_6[406] = ~far_6_6526_1[0]; 
    assign layer_6[407] = ~layer_5[426]; 
    wire [1:0] far_6_6528_0;    relay_conn far_6_6528_0_a(.in(layer_5[176]), .out(far_6_6528_0[0]));    relay_conn far_6_6528_0_b(.in(layer_5[288]), .out(far_6_6528_0[1]));
    wire [1:0] far_6_6528_1;    relay_conn far_6_6528_1_a(.in(far_6_6528_0[0]), .out(far_6_6528_1[0]));    relay_conn far_6_6528_1_b(.in(far_6_6528_0[1]), .out(far_6_6528_1[1]));
    wire [1:0] far_6_6528_2;    relay_conn far_6_6528_2_a(.in(far_6_6528_1[0]), .out(far_6_6528_2[0]));    relay_conn far_6_6528_2_b(.in(far_6_6528_1[1]), .out(far_6_6528_2[1]));
    assign layer_6[408] = ~(far_6_6528_2[0] | far_6_6528_2[1]); 
    wire [1:0] far_6_6529_0;    relay_conn far_6_6529_0_a(.in(layer_5[525]), .out(far_6_6529_0[0]));    relay_conn far_6_6529_0_b(.in(layer_5[617]), .out(far_6_6529_0[1]));
    wire [1:0] far_6_6529_1;    relay_conn far_6_6529_1_a(.in(far_6_6529_0[0]), .out(far_6_6529_1[0]));    relay_conn far_6_6529_1_b(.in(far_6_6529_0[1]), .out(far_6_6529_1[1]));
    assign layer_6[409] = far_6_6529_1[1]; 
    wire [1:0] far_6_6530_0;    relay_conn far_6_6530_0_a(.in(layer_5[384]), .out(far_6_6530_0[0]));    relay_conn far_6_6530_0_b(.in(layer_5[512]), .out(far_6_6530_0[1]));
    wire [1:0] far_6_6530_1;    relay_conn far_6_6530_1_a(.in(far_6_6530_0[0]), .out(far_6_6530_1[0]));    relay_conn far_6_6530_1_b(.in(far_6_6530_0[1]), .out(far_6_6530_1[1]));
    wire [1:0] far_6_6530_2;    relay_conn far_6_6530_2_a(.in(far_6_6530_1[0]), .out(far_6_6530_2[0]));    relay_conn far_6_6530_2_b(.in(far_6_6530_1[1]), .out(far_6_6530_2[1]));
    wire [1:0] far_6_6530_3;    relay_conn far_6_6530_3_a(.in(far_6_6530_2[0]), .out(far_6_6530_3[0]));    relay_conn far_6_6530_3_b(.in(far_6_6530_2[1]), .out(far_6_6530_3[1]));
    assign layer_6[410] = ~far_6_6530_3[1]; 
    wire [1:0] far_6_6531_0;    relay_conn far_6_6531_0_a(.in(layer_5[662]), .out(far_6_6531_0[0]));    relay_conn far_6_6531_0_b(.in(layer_5[629]), .out(far_6_6531_0[1]));
    assign layer_6[411] = far_6_6531_0[0]; 
    wire [1:0] far_6_6532_0;    relay_conn far_6_6532_0_a(.in(layer_5[668]), .out(far_6_6532_0[0]));    relay_conn far_6_6532_0_b(.in(layer_5[599]), .out(far_6_6532_0[1]));
    wire [1:0] far_6_6532_1;    relay_conn far_6_6532_1_a(.in(far_6_6532_0[0]), .out(far_6_6532_1[0]));    relay_conn far_6_6532_1_b(.in(far_6_6532_0[1]), .out(far_6_6532_1[1]));
    assign layer_6[412] = ~(far_6_6532_1[0] & far_6_6532_1[1]); 
    wire [1:0] far_6_6533_0;    relay_conn far_6_6533_0_a(.in(layer_5[695]), .out(far_6_6533_0[0]));    relay_conn far_6_6533_0_b(.in(layer_5[818]), .out(far_6_6533_0[1]));
    wire [1:0] far_6_6533_1;    relay_conn far_6_6533_1_a(.in(far_6_6533_0[0]), .out(far_6_6533_1[0]));    relay_conn far_6_6533_1_b(.in(far_6_6533_0[1]), .out(far_6_6533_1[1]));
    wire [1:0] far_6_6533_2;    relay_conn far_6_6533_2_a(.in(far_6_6533_1[0]), .out(far_6_6533_2[0]));    relay_conn far_6_6533_2_b(.in(far_6_6533_1[1]), .out(far_6_6533_2[1]));
    assign layer_6[413] = ~far_6_6533_2[0]; 
    wire [1:0] far_6_6534_0;    relay_conn far_6_6534_0_a(.in(layer_5[840]), .out(far_6_6534_0[0]));    relay_conn far_6_6534_0_b(.in(layer_5[725]), .out(far_6_6534_0[1]));
    wire [1:0] far_6_6534_1;    relay_conn far_6_6534_1_a(.in(far_6_6534_0[0]), .out(far_6_6534_1[0]));    relay_conn far_6_6534_1_b(.in(far_6_6534_0[1]), .out(far_6_6534_1[1]));
    wire [1:0] far_6_6534_2;    relay_conn far_6_6534_2_a(.in(far_6_6534_1[0]), .out(far_6_6534_2[0]));    relay_conn far_6_6534_2_b(.in(far_6_6534_1[1]), .out(far_6_6534_2[1]));
    assign layer_6[414] = ~far_6_6534_2[1]; 
    wire [1:0] far_6_6535_0;    relay_conn far_6_6535_0_a(.in(layer_5[458]), .out(far_6_6535_0[0]));    relay_conn far_6_6535_0_b(.in(layer_5[539]), .out(far_6_6535_0[1]));
    wire [1:0] far_6_6535_1;    relay_conn far_6_6535_1_a(.in(far_6_6535_0[0]), .out(far_6_6535_1[0]));    relay_conn far_6_6535_1_b(.in(far_6_6535_0[1]), .out(far_6_6535_1[1]));
    assign layer_6[415] = ~far_6_6535_1[0] | (far_6_6535_1[0] & far_6_6535_1[1]); 
    assign layer_6[416] = ~layer_5[763] | (layer_5[763] & layer_5[777]); 
    wire [1:0] far_6_6537_0;    relay_conn far_6_6537_0_a(.in(layer_5[878]), .out(far_6_6537_0[0]));    relay_conn far_6_6537_0_b(.in(layer_5[916]), .out(far_6_6537_0[1]));
    assign layer_6[417] = far_6_6537_0[0] | far_6_6537_0[1]; 
    wire [1:0] far_6_6538_0;    relay_conn far_6_6538_0_a(.in(layer_5[479]), .out(far_6_6538_0[0]));    relay_conn far_6_6538_0_b(.in(layer_5[540]), .out(far_6_6538_0[1]));
    assign layer_6[418] = ~far_6_6538_0[1]; 
    wire [1:0] far_6_6539_0;    relay_conn far_6_6539_0_a(.in(layer_5[684]), .out(far_6_6539_0[0]));    relay_conn far_6_6539_0_b(.in(layer_5[805]), .out(far_6_6539_0[1]));
    wire [1:0] far_6_6539_1;    relay_conn far_6_6539_1_a(.in(far_6_6539_0[0]), .out(far_6_6539_1[0]));    relay_conn far_6_6539_1_b(.in(far_6_6539_0[1]), .out(far_6_6539_1[1]));
    wire [1:0] far_6_6539_2;    relay_conn far_6_6539_2_a(.in(far_6_6539_1[0]), .out(far_6_6539_2[0]));    relay_conn far_6_6539_2_b(.in(far_6_6539_1[1]), .out(far_6_6539_2[1]));
    assign layer_6[419] = ~far_6_6539_2[0]; 
    wire [1:0] far_6_6540_0;    relay_conn far_6_6540_0_a(.in(layer_5[773]), .out(far_6_6540_0[0]));    relay_conn far_6_6540_0_b(.in(layer_5[653]), .out(far_6_6540_0[1]));
    wire [1:0] far_6_6540_1;    relay_conn far_6_6540_1_a(.in(far_6_6540_0[0]), .out(far_6_6540_1[0]));    relay_conn far_6_6540_1_b(.in(far_6_6540_0[1]), .out(far_6_6540_1[1]));
    wire [1:0] far_6_6540_2;    relay_conn far_6_6540_2_a(.in(far_6_6540_1[0]), .out(far_6_6540_2[0]));    relay_conn far_6_6540_2_b(.in(far_6_6540_1[1]), .out(far_6_6540_2[1]));
    assign layer_6[420] = ~far_6_6540_2[0] | (far_6_6540_2[0] & far_6_6540_2[1]); 
    assign layer_6[421] = ~layer_5[849] | (layer_5[849] & layer_5[840]); 
    assign layer_6[422] = layer_5[77]; 
    wire [1:0] far_6_6543_0;    relay_conn far_6_6543_0_a(.in(layer_5[694]), .out(far_6_6543_0[0]));    relay_conn far_6_6543_0_b(.in(layer_5[786]), .out(far_6_6543_0[1]));
    wire [1:0] far_6_6543_1;    relay_conn far_6_6543_1_a(.in(far_6_6543_0[0]), .out(far_6_6543_1[0]));    relay_conn far_6_6543_1_b(.in(far_6_6543_0[1]), .out(far_6_6543_1[1]));
    assign layer_6[423] = ~far_6_6543_1[1] | (far_6_6543_1[0] & far_6_6543_1[1]); 
    wire [1:0] far_6_6544_0;    relay_conn far_6_6544_0_a(.in(layer_5[482]), .out(far_6_6544_0[0]));    relay_conn far_6_6544_0_b(.in(layer_5[598]), .out(far_6_6544_0[1]));
    wire [1:0] far_6_6544_1;    relay_conn far_6_6544_1_a(.in(far_6_6544_0[0]), .out(far_6_6544_1[0]));    relay_conn far_6_6544_1_b(.in(far_6_6544_0[1]), .out(far_6_6544_1[1]));
    wire [1:0] far_6_6544_2;    relay_conn far_6_6544_2_a(.in(far_6_6544_1[0]), .out(far_6_6544_2[0]));    relay_conn far_6_6544_2_b(.in(far_6_6544_1[1]), .out(far_6_6544_2[1]));
    assign layer_6[424] = far_6_6544_2[1]; 
    wire [1:0] far_6_6545_0;    relay_conn far_6_6545_0_a(.in(layer_5[968]), .out(far_6_6545_0[0]));    relay_conn far_6_6545_0_b(.in(layer_5[1017]), .out(far_6_6545_0[1]));
    assign layer_6[425] = ~far_6_6545_0[0]; 
    wire [1:0] far_6_6546_0;    relay_conn far_6_6546_0_a(.in(layer_5[873]), .out(far_6_6546_0[0]));    relay_conn far_6_6546_0_b(.in(layer_5[824]), .out(far_6_6546_0[1]));
    assign layer_6[426] = ~far_6_6546_0[0] | (far_6_6546_0[0] & far_6_6546_0[1]); 
    wire [1:0] far_6_6547_0;    relay_conn far_6_6547_0_a(.in(layer_5[770]), .out(far_6_6547_0[0]));    relay_conn far_6_6547_0_b(.in(layer_5[875]), .out(far_6_6547_0[1]));
    wire [1:0] far_6_6547_1;    relay_conn far_6_6547_1_a(.in(far_6_6547_0[0]), .out(far_6_6547_1[0]));    relay_conn far_6_6547_1_b(.in(far_6_6547_0[1]), .out(far_6_6547_1[1]));
    wire [1:0] far_6_6547_2;    relay_conn far_6_6547_2_a(.in(far_6_6547_1[0]), .out(far_6_6547_2[0]));    relay_conn far_6_6547_2_b(.in(far_6_6547_1[1]), .out(far_6_6547_2[1]));
    assign layer_6[427] = far_6_6547_2[0] & ~far_6_6547_2[1]; 
    wire [1:0] far_6_6548_0;    relay_conn far_6_6548_0_a(.in(layer_5[667]), .out(far_6_6548_0[0]));    relay_conn far_6_6548_0_b(.in(layer_5[613]), .out(far_6_6548_0[1]));
    assign layer_6[428] = far_6_6548_0[0] & ~far_6_6548_0[1]; 
    wire [1:0] far_6_6549_0;    relay_conn far_6_6549_0_a(.in(layer_5[107]), .out(far_6_6549_0[0]));    relay_conn far_6_6549_0_b(.in(layer_5[203]), .out(far_6_6549_0[1]));
    wire [1:0] far_6_6549_1;    relay_conn far_6_6549_1_a(.in(far_6_6549_0[0]), .out(far_6_6549_1[0]));    relay_conn far_6_6549_1_b(.in(far_6_6549_0[1]), .out(far_6_6549_1[1]));
    wire [1:0] far_6_6549_2;    relay_conn far_6_6549_2_a(.in(far_6_6549_1[0]), .out(far_6_6549_2[0]));    relay_conn far_6_6549_2_b(.in(far_6_6549_1[1]), .out(far_6_6549_2[1]));
    assign layer_6[429] = far_6_6549_2[0] | far_6_6549_2[1]; 
    wire [1:0] far_6_6550_0;    relay_conn far_6_6550_0_a(.in(layer_5[480]), .out(far_6_6550_0[0]));    relay_conn far_6_6550_0_b(.in(layer_5[543]), .out(far_6_6550_0[1]));
    assign layer_6[430] = ~far_6_6550_0[1]; 
    wire [1:0] far_6_6551_0;    relay_conn far_6_6551_0_a(.in(layer_5[654]), .out(far_6_6551_0[0]));    relay_conn far_6_6551_0_b(.in(layer_5[561]), .out(far_6_6551_0[1]));
    wire [1:0] far_6_6551_1;    relay_conn far_6_6551_1_a(.in(far_6_6551_0[0]), .out(far_6_6551_1[0]));    relay_conn far_6_6551_1_b(.in(far_6_6551_0[1]), .out(far_6_6551_1[1]));
    assign layer_6[431] = ~(far_6_6551_1[0] | far_6_6551_1[1]); 
    wire [1:0] far_6_6552_0;    relay_conn far_6_6552_0_a(.in(layer_5[219]), .out(far_6_6552_0[0]));    relay_conn far_6_6552_0_b(.in(layer_5[128]), .out(far_6_6552_0[1]));
    wire [1:0] far_6_6552_1;    relay_conn far_6_6552_1_a(.in(far_6_6552_0[0]), .out(far_6_6552_1[0]));    relay_conn far_6_6552_1_b(.in(far_6_6552_0[1]), .out(far_6_6552_1[1]));
    assign layer_6[432] = ~far_6_6552_1[0]; 
    wire [1:0] far_6_6553_0;    relay_conn far_6_6553_0_a(.in(layer_5[457]), .out(far_6_6553_0[0]));    relay_conn far_6_6553_0_b(.in(layer_5[552]), .out(far_6_6553_0[1]));
    wire [1:0] far_6_6553_1;    relay_conn far_6_6553_1_a(.in(far_6_6553_0[0]), .out(far_6_6553_1[0]));    relay_conn far_6_6553_1_b(.in(far_6_6553_0[1]), .out(far_6_6553_1[1]));
    assign layer_6[433] = ~far_6_6553_1[1]; 
    wire [1:0] far_6_6554_0;    relay_conn far_6_6554_0_a(.in(layer_5[474]), .out(far_6_6554_0[0]));    relay_conn far_6_6554_0_b(.in(layer_5[423]), .out(far_6_6554_0[1]));
    assign layer_6[434] = far_6_6554_0[0] & ~far_6_6554_0[1]; 
    wire [1:0] far_6_6555_0;    relay_conn far_6_6555_0_a(.in(layer_5[823]), .out(far_6_6555_0[0]));    relay_conn far_6_6555_0_b(.in(layer_5[741]), .out(far_6_6555_0[1]));
    wire [1:0] far_6_6555_1;    relay_conn far_6_6555_1_a(.in(far_6_6555_0[0]), .out(far_6_6555_1[0]));    relay_conn far_6_6555_1_b(.in(far_6_6555_0[1]), .out(far_6_6555_1[1]));
    assign layer_6[435] = far_6_6555_1[0] & ~far_6_6555_1[1]; 
    wire [1:0] far_6_6556_0;    relay_conn far_6_6556_0_a(.in(layer_5[715]), .out(far_6_6556_0[0]));    relay_conn far_6_6556_0_b(.in(layer_5[637]), .out(far_6_6556_0[1]));
    wire [1:0] far_6_6556_1;    relay_conn far_6_6556_1_a(.in(far_6_6556_0[0]), .out(far_6_6556_1[0]));    relay_conn far_6_6556_1_b(.in(far_6_6556_0[1]), .out(far_6_6556_1[1]));
    assign layer_6[436] = far_6_6556_1[0] | far_6_6556_1[1]; 
    wire [1:0] far_6_6557_0;    relay_conn far_6_6557_0_a(.in(layer_5[615]), .out(far_6_6557_0[0]));    relay_conn far_6_6557_0_b(.in(layer_5[549]), .out(far_6_6557_0[1]));
    wire [1:0] far_6_6557_1;    relay_conn far_6_6557_1_a(.in(far_6_6557_0[0]), .out(far_6_6557_1[0]));    relay_conn far_6_6557_1_b(.in(far_6_6557_0[1]), .out(far_6_6557_1[1]));
    assign layer_6[437] = far_6_6557_1[0] | far_6_6557_1[1]; 
    wire [1:0] far_6_6558_0;    relay_conn far_6_6558_0_a(.in(layer_5[0]), .out(far_6_6558_0[0]));    relay_conn far_6_6558_0_b(.in(layer_5[58]), .out(far_6_6558_0[1]));
    assign layer_6[438] = ~far_6_6558_0[0] | (far_6_6558_0[0] & far_6_6558_0[1]); 
    assign layer_6[439] = layer_5[83]; 
    wire [1:0] far_6_6560_0;    relay_conn far_6_6560_0_a(.in(layer_5[653]), .out(far_6_6560_0[0]));    relay_conn far_6_6560_0_b(.in(layer_5[602]), .out(far_6_6560_0[1]));
    assign layer_6[440] = ~far_6_6560_0[1]; 
    wire [1:0] far_6_6561_0;    relay_conn far_6_6561_0_a(.in(layer_5[263]), .out(far_6_6561_0[0]));    relay_conn far_6_6561_0_b(.in(layer_5[374]), .out(far_6_6561_0[1]));
    wire [1:0] far_6_6561_1;    relay_conn far_6_6561_1_a(.in(far_6_6561_0[0]), .out(far_6_6561_1[0]));    relay_conn far_6_6561_1_b(.in(far_6_6561_0[1]), .out(far_6_6561_1[1]));
    wire [1:0] far_6_6561_2;    relay_conn far_6_6561_2_a(.in(far_6_6561_1[0]), .out(far_6_6561_2[0]));    relay_conn far_6_6561_2_b(.in(far_6_6561_1[1]), .out(far_6_6561_2[1]));
    assign layer_6[441] = ~(far_6_6561_2[0] ^ far_6_6561_2[1]); 
    wire [1:0] far_6_6562_0;    relay_conn far_6_6562_0_a(.in(layer_5[716]), .out(far_6_6562_0[0]));    relay_conn far_6_6562_0_b(.in(layer_5[613]), .out(far_6_6562_0[1]));
    wire [1:0] far_6_6562_1;    relay_conn far_6_6562_1_a(.in(far_6_6562_0[0]), .out(far_6_6562_1[0]));    relay_conn far_6_6562_1_b(.in(far_6_6562_0[1]), .out(far_6_6562_1[1]));
    wire [1:0] far_6_6562_2;    relay_conn far_6_6562_2_a(.in(far_6_6562_1[0]), .out(far_6_6562_2[0]));    relay_conn far_6_6562_2_b(.in(far_6_6562_1[1]), .out(far_6_6562_2[1]));
    assign layer_6[442] = ~far_6_6562_2[1] | (far_6_6562_2[0] & far_6_6562_2[1]); 
    wire [1:0] far_6_6563_0;    relay_conn far_6_6563_0_a(.in(layer_5[892]), .out(far_6_6563_0[0]));    relay_conn far_6_6563_0_b(.in(layer_5[769]), .out(far_6_6563_0[1]));
    wire [1:0] far_6_6563_1;    relay_conn far_6_6563_1_a(.in(far_6_6563_0[0]), .out(far_6_6563_1[0]));    relay_conn far_6_6563_1_b(.in(far_6_6563_0[1]), .out(far_6_6563_1[1]));
    wire [1:0] far_6_6563_2;    relay_conn far_6_6563_2_a(.in(far_6_6563_1[0]), .out(far_6_6563_2[0]));    relay_conn far_6_6563_2_b(.in(far_6_6563_1[1]), .out(far_6_6563_2[1]));
    assign layer_6[443] = ~far_6_6563_2[0]; 
    wire [1:0] far_6_6564_0;    relay_conn far_6_6564_0_a(.in(layer_5[738]), .out(far_6_6564_0[0]));    relay_conn far_6_6564_0_b(.in(layer_5[791]), .out(far_6_6564_0[1]));
    assign layer_6[444] = ~(far_6_6564_0[0] & far_6_6564_0[1]); 
    wire [1:0] far_6_6565_0;    relay_conn far_6_6565_0_a(.in(layer_5[720]), .out(far_6_6565_0[0]));    relay_conn far_6_6565_0_b(.in(layer_5[813]), .out(far_6_6565_0[1]));
    wire [1:0] far_6_6565_1;    relay_conn far_6_6565_1_a(.in(far_6_6565_0[0]), .out(far_6_6565_1[0]));    relay_conn far_6_6565_1_b(.in(far_6_6565_0[1]), .out(far_6_6565_1[1]));
    assign layer_6[445] = far_6_6565_1[0] | far_6_6565_1[1]; 
    wire [1:0] far_6_6566_0;    relay_conn far_6_6566_0_a(.in(layer_5[688]), .out(far_6_6566_0[0]));    relay_conn far_6_6566_0_b(.in(layer_5[760]), .out(far_6_6566_0[1]));
    wire [1:0] far_6_6566_1;    relay_conn far_6_6566_1_a(.in(far_6_6566_0[0]), .out(far_6_6566_1[0]));    relay_conn far_6_6566_1_b(.in(far_6_6566_0[1]), .out(far_6_6566_1[1]));
    assign layer_6[446] = ~far_6_6566_1[1]; 
    wire [1:0] far_6_6567_0;    relay_conn far_6_6567_0_a(.in(layer_5[619]), .out(far_6_6567_0[0]));    relay_conn far_6_6567_0_b(.in(layer_5[746]), .out(far_6_6567_0[1]));
    wire [1:0] far_6_6567_1;    relay_conn far_6_6567_1_a(.in(far_6_6567_0[0]), .out(far_6_6567_1[0]));    relay_conn far_6_6567_1_b(.in(far_6_6567_0[1]), .out(far_6_6567_1[1]));
    wire [1:0] far_6_6567_2;    relay_conn far_6_6567_2_a(.in(far_6_6567_1[0]), .out(far_6_6567_2[0]));    relay_conn far_6_6567_2_b(.in(far_6_6567_1[1]), .out(far_6_6567_2[1]));
    assign layer_6[447] = ~far_6_6567_2[0]; 
    wire [1:0] far_6_6568_0;    relay_conn far_6_6568_0_a(.in(layer_5[793]), .out(far_6_6568_0[0]));    relay_conn far_6_6568_0_b(.in(layer_5[894]), .out(far_6_6568_0[1]));
    wire [1:0] far_6_6568_1;    relay_conn far_6_6568_1_a(.in(far_6_6568_0[0]), .out(far_6_6568_1[0]));    relay_conn far_6_6568_1_b(.in(far_6_6568_0[1]), .out(far_6_6568_1[1]));
    wire [1:0] far_6_6568_2;    relay_conn far_6_6568_2_a(.in(far_6_6568_1[0]), .out(far_6_6568_2[0]));    relay_conn far_6_6568_2_b(.in(far_6_6568_1[1]), .out(far_6_6568_2[1]));
    assign layer_6[448] = far_6_6568_2[0] & far_6_6568_2[1]; 
    wire [1:0] far_6_6569_0;    relay_conn far_6_6569_0_a(.in(layer_5[865]), .out(far_6_6569_0[0]));    relay_conn far_6_6569_0_b(.in(layer_5[738]), .out(far_6_6569_0[1]));
    wire [1:0] far_6_6569_1;    relay_conn far_6_6569_1_a(.in(far_6_6569_0[0]), .out(far_6_6569_1[0]));    relay_conn far_6_6569_1_b(.in(far_6_6569_0[1]), .out(far_6_6569_1[1]));
    wire [1:0] far_6_6569_2;    relay_conn far_6_6569_2_a(.in(far_6_6569_1[0]), .out(far_6_6569_2[0]));    relay_conn far_6_6569_2_b(.in(far_6_6569_1[1]), .out(far_6_6569_2[1]));
    assign layer_6[449] = ~far_6_6569_2[0]; 
    wire [1:0] far_6_6570_0;    relay_conn far_6_6570_0_a(.in(layer_5[401]), .out(far_6_6570_0[0]));    relay_conn far_6_6570_0_b(.in(layer_5[505]), .out(far_6_6570_0[1]));
    wire [1:0] far_6_6570_1;    relay_conn far_6_6570_1_a(.in(far_6_6570_0[0]), .out(far_6_6570_1[0]));    relay_conn far_6_6570_1_b(.in(far_6_6570_0[1]), .out(far_6_6570_1[1]));
    wire [1:0] far_6_6570_2;    relay_conn far_6_6570_2_a(.in(far_6_6570_1[0]), .out(far_6_6570_2[0]));    relay_conn far_6_6570_2_b(.in(far_6_6570_1[1]), .out(far_6_6570_2[1]));
    assign layer_6[450] = far_6_6570_2[0] & ~far_6_6570_2[1]; 
    wire [1:0] far_6_6571_0;    relay_conn far_6_6571_0_a(.in(layer_5[793]), .out(far_6_6571_0[0]));    relay_conn far_6_6571_0_b(.in(layer_5[741]), .out(far_6_6571_0[1]));
    assign layer_6[451] = ~far_6_6571_0[1] | (far_6_6571_0[0] & far_6_6571_0[1]); 
    wire [1:0] far_6_6572_0;    relay_conn far_6_6572_0_a(.in(layer_5[689]), .out(far_6_6572_0[0]));    relay_conn far_6_6572_0_b(.in(layer_5[758]), .out(far_6_6572_0[1]));
    wire [1:0] far_6_6572_1;    relay_conn far_6_6572_1_a(.in(far_6_6572_0[0]), .out(far_6_6572_1[0]));    relay_conn far_6_6572_1_b(.in(far_6_6572_0[1]), .out(far_6_6572_1[1]));
    assign layer_6[452] = ~far_6_6572_1[1] | (far_6_6572_1[0] & far_6_6572_1[1]); 
    wire [1:0] far_6_6573_0;    relay_conn far_6_6573_0_a(.in(layer_5[401]), .out(far_6_6573_0[0]));    relay_conn far_6_6573_0_b(.in(layer_5[436]), .out(far_6_6573_0[1]));
    assign layer_6[453] = ~far_6_6573_0[0]; 
    wire [1:0] far_6_6574_0;    relay_conn far_6_6574_0_a(.in(layer_5[724]), .out(far_6_6574_0[0]));    relay_conn far_6_6574_0_b(.in(layer_5[758]), .out(far_6_6574_0[1]));
    assign layer_6[454] = ~(far_6_6574_0[0] & far_6_6574_0[1]); 
    wire [1:0] far_6_6575_0;    relay_conn far_6_6575_0_a(.in(layer_5[404]), .out(far_6_6575_0[0]));    relay_conn far_6_6575_0_b(.in(layer_5[504]), .out(far_6_6575_0[1]));
    wire [1:0] far_6_6575_1;    relay_conn far_6_6575_1_a(.in(far_6_6575_0[0]), .out(far_6_6575_1[0]));    relay_conn far_6_6575_1_b(.in(far_6_6575_0[1]), .out(far_6_6575_1[1]));
    wire [1:0] far_6_6575_2;    relay_conn far_6_6575_2_a(.in(far_6_6575_1[0]), .out(far_6_6575_2[0]));    relay_conn far_6_6575_2_b(.in(far_6_6575_1[1]), .out(far_6_6575_2[1]));
    assign layer_6[455] = far_6_6575_2[0]; 
    wire [1:0] far_6_6576_0;    relay_conn far_6_6576_0_a(.in(layer_5[125]), .out(far_6_6576_0[0]));    relay_conn far_6_6576_0_b(.in(layer_5[60]), .out(far_6_6576_0[1]));
    wire [1:0] far_6_6576_1;    relay_conn far_6_6576_1_a(.in(far_6_6576_0[0]), .out(far_6_6576_1[0]));    relay_conn far_6_6576_1_b(.in(far_6_6576_0[1]), .out(far_6_6576_1[1]));
    assign layer_6[456] = ~(far_6_6576_1[0] & far_6_6576_1[1]); 
    assign layer_6[457] = layer_5[1019] ^ layer_5[996]; 
    wire [1:0] far_6_6578_0;    relay_conn far_6_6578_0_a(.in(layer_5[552]), .out(far_6_6578_0[0]));    relay_conn far_6_6578_0_b(.in(layer_5[430]), .out(far_6_6578_0[1]));
    wire [1:0] far_6_6578_1;    relay_conn far_6_6578_1_a(.in(far_6_6578_0[0]), .out(far_6_6578_1[0]));    relay_conn far_6_6578_1_b(.in(far_6_6578_0[1]), .out(far_6_6578_1[1]));
    wire [1:0] far_6_6578_2;    relay_conn far_6_6578_2_a(.in(far_6_6578_1[0]), .out(far_6_6578_2[0]));    relay_conn far_6_6578_2_b(.in(far_6_6578_1[1]), .out(far_6_6578_2[1]));
    assign layer_6[458] = far_6_6578_2[1]; 
    assign layer_6[459] = ~layer_5[592] | (layer_5[567] & layer_5[592]); 
    wire [1:0] far_6_6580_0;    relay_conn far_6_6580_0_a(.in(layer_5[951]), .out(far_6_6580_0[0]));    relay_conn far_6_6580_0_b(.in(layer_5[888]), .out(far_6_6580_0[1]));
    assign layer_6[460] = far_6_6580_0[0]; 
    assign layer_6[461] = layer_5[187] & ~layer_5[203]; 
    assign layer_6[462] = ~(layer_5[888] | layer_5[858]); 
    assign layer_6[463] = ~(layer_5[396] | layer_5[424]); 
    wire [1:0] far_6_6584_0;    relay_conn far_6_6584_0_a(.in(layer_5[558]), .out(far_6_6584_0[0]));    relay_conn far_6_6584_0_b(.in(layer_5[454]), .out(far_6_6584_0[1]));
    wire [1:0] far_6_6584_1;    relay_conn far_6_6584_1_a(.in(far_6_6584_0[0]), .out(far_6_6584_1[0]));    relay_conn far_6_6584_1_b(.in(far_6_6584_0[1]), .out(far_6_6584_1[1]));
    wire [1:0] far_6_6584_2;    relay_conn far_6_6584_2_a(.in(far_6_6584_1[0]), .out(far_6_6584_2[0]));    relay_conn far_6_6584_2_b(.in(far_6_6584_1[1]), .out(far_6_6584_2[1]));
    assign layer_6[464] = ~far_6_6584_2[1] | (far_6_6584_2[0] & far_6_6584_2[1]); 
    wire [1:0] far_6_6585_0;    relay_conn far_6_6585_0_a(.in(layer_5[480]), .out(far_6_6585_0[0]));    relay_conn far_6_6585_0_b(.in(layer_5[599]), .out(far_6_6585_0[1]));
    wire [1:0] far_6_6585_1;    relay_conn far_6_6585_1_a(.in(far_6_6585_0[0]), .out(far_6_6585_1[0]));    relay_conn far_6_6585_1_b(.in(far_6_6585_0[1]), .out(far_6_6585_1[1]));
    wire [1:0] far_6_6585_2;    relay_conn far_6_6585_2_a(.in(far_6_6585_1[0]), .out(far_6_6585_2[0]));    relay_conn far_6_6585_2_b(.in(far_6_6585_1[1]), .out(far_6_6585_2[1]));
    assign layer_6[465] = ~far_6_6585_2[1]; 
    wire [1:0] far_6_6586_0;    relay_conn far_6_6586_0_a(.in(layer_5[185]), .out(far_6_6586_0[0]));    relay_conn far_6_6586_0_b(.in(layer_5[153]), .out(far_6_6586_0[1]));
    assign layer_6[466] = ~(far_6_6586_0[0] ^ far_6_6586_0[1]); 
    wire [1:0] far_6_6587_0;    relay_conn far_6_6587_0_a(.in(layer_5[149]), .out(far_6_6587_0[0]));    relay_conn far_6_6587_0_b(.in(layer_5[107]), .out(far_6_6587_0[1]));
    assign layer_6[467] = ~(far_6_6587_0[0] & far_6_6587_0[1]); 
    wire [1:0] far_6_6588_0;    relay_conn far_6_6588_0_a(.in(layer_5[190]), .out(far_6_6588_0[0]));    relay_conn far_6_6588_0_b(.in(layer_5[315]), .out(far_6_6588_0[1]));
    wire [1:0] far_6_6588_1;    relay_conn far_6_6588_1_a(.in(far_6_6588_0[0]), .out(far_6_6588_1[0]));    relay_conn far_6_6588_1_b(.in(far_6_6588_0[1]), .out(far_6_6588_1[1]));
    wire [1:0] far_6_6588_2;    relay_conn far_6_6588_2_a(.in(far_6_6588_1[0]), .out(far_6_6588_2[0]));    relay_conn far_6_6588_2_b(.in(far_6_6588_1[1]), .out(far_6_6588_2[1]));
    assign layer_6[468] = ~(far_6_6588_2[0] & far_6_6588_2[1]); 
    wire [1:0] far_6_6589_0;    relay_conn far_6_6589_0_a(.in(layer_5[772]), .out(far_6_6589_0[0]));    relay_conn far_6_6589_0_b(.in(layer_5[886]), .out(far_6_6589_0[1]));
    wire [1:0] far_6_6589_1;    relay_conn far_6_6589_1_a(.in(far_6_6589_0[0]), .out(far_6_6589_1[0]));    relay_conn far_6_6589_1_b(.in(far_6_6589_0[1]), .out(far_6_6589_1[1]));
    wire [1:0] far_6_6589_2;    relay_conn far_6_6589_2_a(.in(far_6_6589_1[0]), .out(far_6_6589_2[0]));    relay_conn far_6_6589_2_b(.in(far_6_6589_1[1]), .out(far_6_6589_2[1]));
    assign layer_6[469] = ~far_6_6589_2[1] | (far_6_6589_2[0] & far_6_6589_2[1]); 
    assign layer_6[470] = ~layer_5[640]; 
    assign layer_6[471] = ~layer_5[790]; 
    assign layer_6[472] = layer_5[246]; 
    assign layer_6[473] = ~layer_5[79] | (layer_5[98] & layer_5[79]); 
    assign layer_6[474] = ~(layer_5[748] ^ layer_5[717]); 
    assign layer_6[475] = ~layer_5[178]; 
    assign layer_6[476] = layer_5[956]; 
    wire [1:0] far_6_6597_0;    relay_conn far_6_6597_0_a(.in(layer_5[777]), .out(far_6_6597_0[0]));    relay_conn far_6_6597_0_b(.in(layer_5[734]), .out(far_6_6597_0[1]));
    assign layer_6[477] = ~far_6_6597_0[1] | (far_6_6597_0[0] & far_6_6597_0[1]); 
    wire [1:0] far_6_6598_0;    relay_conn far_6_6598_0_a(.in(layer_5[631]), .out(far_6_6598_0[0]));    relay_conn far_6_6598_0_b(.in(layer_5[598]), .out(far_6_6598_0[1]));
    assign layer_6[478] = ~far_6_6598_0[0]; 
    assign layer_6[479] = layer_5[746] & layer_5[755]; 
    wire [1:0] far_6_6600_0;    relay_conn far_6_6600_0_a(.in(layer_5[197]), .out(far_6_6600_0[0]));    relay_conn far_6_6600_0_b(.in(layer_5[254]), .out(far_6_6600_0[1]));
    assign layer_6[480] = ~far_6_6600_0[1]; 
    assign layer_6[481] = ~layer_5[161]; 
    wire [1:0] far_6_6602_0;    relay_conn far_6_6602_0_a(.in(layer_5[961]), .out(far_6_6602_0[0]));    relay_conn far_6_6602_0_b(.in(layer_5[862]), .out(far_6_6602_0[1]));
    wire [1:0] far_6_6602_1;    relay_conn far_6_6602_1_a(.in(far_6_6602_0[0]), .out(far_6_6602_1[0]));    relay_conn far_6_6602_1_b(.in(far_6_6602_0[1]), .out(far_6_6602_1[1]));
    wire [1:0] far_6_6602_2;    relay_conn far_6_6602_2_a(.in(far_6_6602_1[0]), .out(far_6_6602_2[0]));    relay_conn far_6_6602_2_b(.in(far_6_6602_1[1]), .out(far_6_6602_2[1]));
    assign layer_6[482] = ~(far_6_6602_2[0] | far_6_6602_2[1]); 
    wire [1:0] far_6_6603_0;    relay_conn far_6_6603_0_a(.in(layer_5[83]), .out(far_6_6603_0[0]));    relay_conn far_6_6603_0_b(.in(layer_5[45]), .out(far_6_6603_0[1]));
    assign layer_6[483] = ~(far_6_6603_0[0] & far_6_6603_0[1]); 
    wire [1:0] far_6_6604_0;    relay_conn far_6_6604_0_a(.in(layer_5[106]), .out(far_6_6604_0[0]));    relay_conn far_6_6604_0_b(.in(layer_5[218]), .out(far_6_6604_0[1]));
    wire [1:0] far_6_6604_1;    relay_conn far_6_6604_1_a(.in(far_6_6604_0[0]), .out(far_6_6604_1[0]));    relay_conn far_6_6604_1_b(.in(far_6_6604_0[1]), .out(far_6_6604_1[1]));
    wire [1:0] far_6_6604_2;    relay_conn far_6_6604_2_a(.in(far_6_6604_1[0]), .out(far_6_6604_2[0]));    relay_conn far_6_6604_2_b(.in(far_6_6604_1[1]), .out(far_6_6604_2[1]));
    assign layer_6[484] = ~far_6_6604_2[1]; 
    wire [1:0] far_6_6605_0;    relay_conn far_6_6605_0_a(.in(layer_5[922]), .out(far_6_6605_0[0]));    relay_conn far_6_6605_0_b(.in(layer_5[1002]), .out(far_6_6605_0[1]));
    wire [1:0] far_6_6605_1;    relay_conn far_6_6605_1_a(.in(far_6_6605_0[0]), .out(far_6_6605_1[0]));    relay_conn far_6_6605_1_b(.in(far_6_6605_0[1]), .out(far_6_6605_1[1]));
    assign layer_6[485] = far_6_6605_1[0]; 
    wire [1:0] far_6_6606_0;    relay_conn far_6_6606_0_a(.in(layer_5[98]), .out(far_6_6606_0[0]));    relay_conn far_6_6606_0_b(.in(layer_5[196]), .out(far_6_6606_0[1]));
    wire [1:0] far_6_6606_1;    relay_conn far_6_6606_1_a(.in(far_6_6606_0[0]), .out(far_6_6606_1[0]));    relay_conn far_6_6606_1_b(.in(far_6_6606_0[1]), .out(far_6_6606_1[1]));
    wire [1:0] far_6_6606_2;    relay_conn far_6_6606_2_a(.in(far_6_6606_1[0]), .out(far_6_6606_2[0]));    relay_conn far_6_6606_2_b(.in(far_6_6606_1[1]), .out(far_6_6606_2[1]));
    assign layer_6[486] = far_6_6606_2[1]; 
    wire [1:0] far_6_6607_0;    relay_conn far_6_6607_0_a(.in(layer_5[469]), .out(far_6_6607_0[0]));    relay_conn far_6_6607_0_b(.in(layer_5[370]), .out(far_6_6607_0[1]));
    wire [1:0] far_6_6607_1;    relay_conn far_6_6607_1_a(.in(far_6_6607_0[0]), .out(far_6_6607_1[0]));    relay_conn far_6_6607_1_b(.in(far_6_6607_0[1]), .out(far_6_6607_1[1]));
    wire [1:0] far_6_6607_2;    relay_conn far_6_6607_2_a(.in(far_6_6607_1[0]), .out(far_6_6607_2[0]));    relay_conn far_6_6607_2_b(.in(far_6_6607_1[1]), .out(far_6_6607_2[1]));
    assign layer_6[487] = ~(far_6_6607_2[0] | far_6_6607_2[1]); 
    wire [1:0] far_6_6608_0;    relay_conn far_6_6608_0_a(.in(layer_5[804]), .out(far_6_6608_0[0]));    relay_conn far_6_6608_0_b(.in(layer_5[761]), .out(far_6_6608_0[1]));
    assign layer_6[488] = far_6_6608_0[0] | far_6_6608_0[1]; 
    wire [1:0] far_6_6609_0;    relay_conn far_6_6609_0_a(.in(layer_5[550]), .out(far_6_6609_0[0]));    relay_conn far_6_6609_0_b(.in(layer_5[471]), .out(far_6_6609_0[1]));
    wire [1:0] far_6_6609_1;    relay_conn far_6_6609_1_a(.in(far_6_6609_0[0]), .out(far_6_6609_1[0]));    relay_conn far_6_6609_1_b(.in(far_6_6609_0[1]), .out(far_6_6609_1[1]));
    assign layer_6[489] = ~far_6_6609_1[1]; 
    wire [1:0] far_6_6610_0;    relay_conn far_6_6610_0_a(.in(layer_5[147]), .out(far_6_6610_0[0]));    relay_conn far_6_6610_0_b(.in(layer_5[25]), .out(far_6_6610_0[1]));
    wire [1:0] far_6_6610_1;    relay_conn far_6_6610_1_a(.in(far_6_6610_0[0]), .out(far_6_6610_1[0]));    relay_conn far_6_6610_1_b(.in(far_6_6610_0[1]), .out(far_6_6610_1[1]));
    wire [1:0] far_6_6610_2;    relay_conn far_6_6610_2_a(.in(far_6_6610_1[0]), .out(far_6_6610_2[0]));    relay_conn far_6_6610_2_b(.in(far_6_6610_1[1]), .out(far_6_6610_2[1]));
    assign layer_6[490] = ~(far_6_6610_2[0] | far_6_6610_2[1]); 
    assign layer_6[491] = layer_5[621]; 
    assign layer_6[492] = ~layer_5[424]; 
    wire [1:0] far_6_6613_0;    relay_conn far_6_6613_0_a(.in(layer_5[394]), .out(far_6_6613_0[0]));    relay_conn far_6_6613_0_b(.in(layer_5[351]), .out(far_6_6613_0[1]));
    assign layer_6[493] = far_6_6613_0[1]; 
    assign layer_6[494] = ~layer_5[369] | (layer_5[394] & layer_5[369]); 
    wire [1:0] far_6_6615_0;    relay_conn far_6_6615_0_a(.in(layer_5[687]), .out(far_6_6615_0[0]));    relay_conn far_6_6615_0_b(.in(layer_5[759]), .out(far_6_6615_0[1]));
    wire [1:0] far_6_6615_1;    relay_conn far_6_6615_1_a(.in(far_6_6615_0[0]), .out(far_6_6615_1[0]));    relay_conn far_6_6615_1_b(.in(far_6_6615_0[1]), .out(far_6_6615_1[1]));
    assign layer_6[495] = ~far_6_6615_1[1] | (far_6_6615_1[0] & far_6_6615_1[1]); 
    wire [1:0] far_6_6616_0;    relay_conn far_6_6616_0_a(.in(layer_5[602]), .out(far_6_6616_0[0]));    relay_conn far_6_6616_0_b(.in(layer_5[505]), .out(far_6_6616_0[1]));
    wire [1:0] far_6_6616_1;    relay_conn far_6_6616_1_a(.in(far_6_6616_0[0]), .out(far_6_6616_1[0]));    relay_conn far_6_6616_1_b(.in(far_6_6616_0[1]), .out(far_6_6616_1[1]));
    wire [1:0] far_6_6616_2;    relay_conn far_6_6616_2_a(.in(far_6_6616_1[0]), .out(far_6_6616_2[0]));    relay_conn far_6_6616_2_b(.in(far_6_6616_1[1]), .out(far_6_6616_2[1]));
    assign layer_6[496] = ~far_6_6616_2[0] | (far_6_6616_2[0] & far_6_6616_2[1]); 
    wire [1:0] far_6_6617_0;    relay_conn far_6_6617_0_a(.in(layer_5[640]), .out(far_6_6617_0[0]));    relay_conn far_6_6617_0_b(.in(layer_5[746]), .out(far_6_6617_0[1]));
    wire [1:0] far_6_6617_1;    relay_conn far_6_6617_1_a(.in(far_6_6617_0[0]), .out(far_6_6617_1[0]));    relay_conn far_6_6617_1_b(.in(far_6_6617_0[1]), .out(far_6_6617_1[1]));
    wire [1:0] far_6_6617_2;    relay_conn far_6_6617_2_a(.in(far_6_6617_1[0]), .out(far_6_6617_2[0]));    relay_conn far_6_6617_2_b(.in(far_6_6617_1[1]), .out(far_6_6617_2[1]));
    assign layer_6[497] = ~far_6_6617_2[0]; 
    wire [1:0] far_6_6618_0;    relay_conn far_6_6618_0_a(.in(layer_5[60]), .out(far_6_6618_0[0]));    relay_conn far_6_6618_0_b(.in(layer_5[7]), .out(far_6_6618_0[1]));
    assign layer_6[498] = far_6_6618_0[0] | far_6_6618_0[1]; 
    wire [1:0] far_6_6619_0;    relay_conn far_6_6619_0_a(.in(layer_5[643]), .out(far_6_6619_0[0]));    relay_conn far_6_6619_0_b(.in(layer_5[588]), .out(far_6_6619_0[1]));
    assign layer_6[499] = ~(far_6_6619_0[0] ^ far_6_6619_0[1]); 
    wire [1:0] far_6_6620_0;    relay_conn far_6_6620_0_a(.in(layer_5[629]), .out(far_6_6620_0[0]));    relay_conn far_6_6620_0_b(.in(layer_5[748]), .out(far_6_6620_0[1]));
    wire [1:0] far_6_6620_1;    relay_conn far_6_6620_1_a(.in(far_6_6620_0[0]), .out(far_6_6620_1[0]));    relay_conn far_6_6620_1_b(.in(far_6_6620_0[1]), .out(far_6_6620_1[1]));
    wire [1:0] far_6_6620_2;    relay_conn far_6_6620_2_a(.in(far_6_6620_1[0]), .out(far_6_6620_2[0]));    relay_conn far_6_6620_2_b(.in(far_6_6620_1[1]), .out(far_6_6620_2[1]));
    assign layer_6[500] = ~far_6_6620_2[0]; 
    wire [1:0] far_6_6621_0;    relay_conn far_6_6621_0_a(.in(layer_5[258]), .out(far_6_6621_0[0]));    relay_conn far_6_6621_0_b(.in(layer_5[150]), .out(far_6_6621_0[1]));
    wire [1:0] far_6_6621_1;    relay_conn far_6_6621_1_a(.in(far_6_6621_0[0]), .out(far_6_6621_1[0]));    relay_conn far_6_6621_1_b(.in(far_6_6621_0[1]), .out(far_6_6621_1[1]));
    wire [1:0] far_6_6621_2;    relay_conn far_6_6621_2_a(.in(far_6_6621_1[0]), .out(far_6_6621_2[0]));    relay_conn far_6_6621_2_b(.in(far_6_6621_1[1]), .out(far_6_6621_2[1]));
    assign layer_6[501] = far_6_6621_2[0] ^ far_6_6621_2[1]; 
    assign layer_6[502] = ~(layer_5[758] & layer_5[730]); 
    wire [1:0] far_6_6623_0;    relay_conn far_6_6623_0_a(.in(layer_5[222]), .out(far_6_6623_0[0]));    relay_conn far_6_6623_0_b(.in(layer_5[168]), .out(far_6_6623_0[1]));
    assign layer_6[503] = far_6_6623_0[1]; 
    wire [1:0] far_6_6624_0;    relay_conn far_6_6624_0_a(.in(layer_5[585]), .out(far_6_6624_0[0]));    relay_conn far_6_6624_0_b(.in(layer_5[668]), .out(far_6_6624_0[1]));
    wire [1:0] far_6_6624_1;    relay_conn far_6_6624_1_a(.in(far_6_6624_0[0]), .out(far_6_6624_1[0]));    relay_conn far_6_6624_1_b(.in(far_6_6624_0[1]), .out(far_6_6624_1[1]));
    assign layer_6[504] = ~(far_6_6624_1[0] | far_6_6624_1[1]); 
    wire [1:0] far_6_6625_0;    relay_conn far_6_6625_0_a(.in(layer_5[913]), .out(far_6_6625_0[0]));    relay_conn far_6_6625_0_b(.in(layer_5[793]), .out(far_6_6625_0[1]));
    wire [1:0] far_6_6625_1;    relay_conn far_6_6625_1_a(.in(far_6_6625_0[0]), .out(far_6_6625_1[0]));    relay_conn far_6_6625_1_b(.in(far_6_6625_0[1]), .out(far_6_6625_1[1]));
    wire [1:0] far_6_6625_2;    relay_conn far_6_6625_2_a(.in(far_6_6625_1[0]), .out(far_6_6625_2[0]));    relay_conn far_6_6625_2_b(.in(far_6_6625_1[1]), .out(far_6_6625_2[1]));
    assign layer_6[505] = far_6_6625_2[1] & ~far_6_6625_2[0]; 
    wire [1:0] far_6_6626_0;    relay_conn far_6_6626_0_a(.in(layer_5[489]), .out(far_6_6626_0[0]));    relay_conn far_6_6626_0_b(.in(layer_5[590]), .out(far_6_6626_0[1]));
    wire [1:0] far_6_6626_1;    relay_conn far_6_6626_1_a(.in(far_6_6626_0[0]), .out(far_6_6626_1[0]));    relay_conn far_6_6626_1_b(.in(far_6_6626_0[1]), .out(far_6_6626_1[1]));
    wire [1:0] far_6_6626_2;    relay_conn far_6_6626_2_a(.in(far_6_6626_1[0]), .out(far_6_6626_2[0]));    relay_conn far_6_6626_2_b(.in(far_6_6626_1[1]), .out(far_6_6626_2[1]));
    assign layer_6[506] = far_6_6626_2[0] ^ far_6_6626_2[1]; 
    wire [1:0] far_6_6627_0;    relay_conn far_6_6627_0_a(.in(layer_5[717]), .out(far_6_6627_0[0]));    relay_conn far_6_6627_0_b(.in(layer_5[629]), .out(far_6_6627_0[1]));
    wire [1:0] far_6_6627_1;    relay_conn far_6_6627_1_a(.in(far_6_6627_0[0]), .out(far_6_6627_1[0]));    relay_conn far_6_6627_1_b(.in(far_6_6627_0[1]), .out(far_6_6627_1[1]));
    assign layer_6[507] = ~(far_6_6627_1[0] & far_6_6627_1[1]); 
    wire [1:0] far_6_6628_0;    relay_conn far_6_6628_0_a(.in(layer_5[535]), .out(far_6_6628_0[0]));    relay_conn far_6_6628_0_b(.in(layer_5[599]), .out(far_6_6628_0[1]));
    wire [1:0] far_6_6628_1;    relay_conn far_6_6628_1_a(.in(far_6_6628_0[0]), .out(far_6_6628_1[0]));    relay_conn far_6_6628_1_b(.in(far_6_6628_0[1]), .out(far_6_6628_1[1]));
    assign layer_6[508] = ~far_6_6628_1[0]; 
    wire [1:0] far_6_6629_0;    relay_conn far_6_6629_0_a(.in(layer_5[585]), .out(far_6_6629_0[0]));    relay_conn far_6_6629_0_b(.in(layer_5[537]), .out(far_6_6629_0[1]));
    assign layer_6[509] = far_6_6629_0[0] & far_6_6629_0[1]; 
    wire [1:0] far_6_6630_0;    relay_conn far_6_6630_0_a(.in(layer_5[424]), .out(far_6_6630_0[0]));    relay_conn far_6_6630_0_b(.in(layer_5[509]), .out(far_6_6630_0[1]));
    wire [1:0] far_6_6630_1;    relay_conn far_6_6630_1_a(.in(far_6_6630_0[0]), .out(far_6_6630_1[0]));    relay_conn far_6_6630_1_b(.in(far_6_6630_0[1]), .out(far_6_6630_1[1]));
    assign layer_6[510] = ~far_6_6630_1[0]; 
    wire [1:0] far_6_6631_0;    relay_conn far_6_6631_0_a(.in(layer_5[63]), .out(far_6_6631_0[0]));    relay_conn far_6_6631_0_b(.in(layer_5[122]), .out(far_6_6631_0[1]));
    assign layer_6[511] = far_6_6631_0[0] & far_6_6631_0[1]; 
    wire [1:0] far_6_6632_0;    relay_conn far_6_6632_0_a(.in(layer_5[547]), .out(far_6_6632_0[0]));    relay_conn far_6_6632_0_b(.in(layer_5[593]), .out(far_6_6632_0[1]));
    assign layer_6[512] = ~far_6_6632_0[0]; 
    wire [1:0] far_6_6633_0;    relay_conn far_6_6633_0_a(.in(layer_5[605]), .out(far_6_6633_0[0]));    relay_conn far_6_6633_0_b(.in(layer_5[550]), .out(far_6_6633_0[1]));
    assign layer_6[513] = far_6_6633_0[0]; 
    wire [1:0] far_6_6634_0;    relay_conn far_6_6634_0_a(.in(layer_5[101]), .out(far_6_6634_0[0]));    relay_conn far_6_6634_0_b(.in(layer_5[149]), .out(far_6_6634_0[1]));
    assign layer_6[514] = far_6_6634_0[0] & far_6_6634_0[1]; 
    wire [1:0] far_6_6635_0;    relay_conn far_6_6635_0_a(.in(layer_5[78]), .out(far_6_6635_0[0]));    relay_conn far_6_6635_0_b(.in(layer_5[111]), .out(far_6_6635_0[1]));
    assign layer_6[515] = ~(far_6_6635_0[0] | far_6_6635_0[1]); 
    wire [1:0] far_6_6636_0;    relay_conn far_6_6636_0_a(.in(layer_5[963]), .out(far_6_6636_0[0]));    relay_conn far_6_6636_0_b(.in(layer_5[871]), .out(far_6_6636_0[1]));
    wire [1:0] far_6_6636_1;    relay_conn far_6_6636_1_a(.in(far_6_6636_0[0]), .out(far_6_6636_1[0]));    relay_conn far_6_6636_1_b(.in(far_6_6636_0[1]), .out(far_6_6636_1[1]));
    assign layer_6[516] = ~far_6_6636_1[1]; 
    assign layer_6[517] = ~layer_5[362]; 
    wire [1:0] far_6_6638_0;    relay_conn far_6_6638_0_a(.in(layer_5[679]), .out(far_6_6638_0[0]));    relay_conn far_6_6638_0_b(.in(layer_5[765]), .out(far_6_6638_0[1]));
    wire [1:0] far_6_6638_1;    relay_conn far_6_6638_1_a(.in(far_6_6638_0[0]), .out(far_6_6638_1[0]));    relay_conn far_6_6638_1_b(.in(far_6_6638_0[1]), .out(far_6_6638_1[1]));
    assign layer_6[518] = ~(far_6_6638_1[0] ^ far_6_6638_1[1]); 
    wire [1:0] far_6_6639_0;    relay_conn far_6_6639_0_a(.in(layer_5[346]), .out(far_6_6639_0[0]));    relay_conn far_6_6639_0_b(.in(layer_5[430]), .out(far_6_6639_0[1]));
    wire [1:0] far_6_6639_1;    relay_conn far_6_6639_1_a(.in(far_6_6639_0[0]), .out(far_6_6639_1[0]));    relay_conn far_6_6639_1_b(.in(far_6_6639_0[1]), .out(far_6_6639_1[1]));
    assign layer_6[519] = far_6_6639_1[0] ^ far_6_6639_1[1]; 
    wire [1:0] far_6_6640_0;    relay_conn far_6_6640_0_a(.in(layer_5[660]), .out(far_6_6640_0[0]));    relay_conn far_6_6640_0_b(.in(layer_5[550]), .out(far_6_6640_0[1]));
    wire [1:0] far_6_6640_1;    relay_conn far_6_6640_1_a(.in(far_6_6640_0[0]), .out(far_6_6640_1[0]));    relay_conn far_6_6640_1_b(.in(far_6_6640_0[1]), .out(far_6_6640_1[1]));
    wire [1:0] far_6_6640_2;    relay_conn far_6_6640_2_a(.in(far_6_6640_1[0]), .out(far_6_6640_2[0]));    relay_conn far_6_6640_2_b(.in(far_6_6640_1[1]), .out(far_6_6640_2[1]));
    assign layer_6[520] = far_6_6640_2[0] ^ far_6_6640_2[1]; 
    wire [1:0] far_6_6641_0;    relay_conn far_6_6641_0_a(.in(layer_5[921]), .out(far_6_6641_0[0]));    relay_conn far_6_6641_0_b(.in(layer_5[845]), .out(far_6_6641_0[1]));
    wire [1:0] far_6_6641_1;    relay_conn far_6_6641_1_a(.in(far_6_6641_0[0]), .out(far_6_6641_1[0]));    relay_conn far_6_6641_1_b(.in(far_6_6641_0[1]), .out(far_6_6641_1[1]));
    assign layer_6[521] = far_6_6641_1[1]; 
    wire [1:0] far_6_6642_0;    relay_conn far_6_6642_0_a(.in(layer_5[875]), .out(far_6_6642_0[0]));    relay_conn far_6_6642_0_b(.in(layer_5[958]), .out(far_6_6642_0[1]));
    wire [1:0] far_6_6642_1;    relay_conn far_6_6642_1_a(.in(far_6_6642_0[0]), .out(far_6_6642_1[0]));    relay_conn far_6_6642_1_b(.in(far_6_6642_0[1]), .out(far_6_6642_1[1]));
    assign layer_6[522] = far_6_6642_1[1]; 
    wire [1:0] far_6_6643_0;    relay_conn far_6_6643_0_a(.in(layer_5[312]), .out(far_6_6643_0[0]));    relay_conn far_6_6643_0_b(.in(layer_5[396]), .out(far_6_6643_0[1]));
    wire [1:0] far_6_6643_1;    relay_conn far_6_6643_1_a(.in(far_6_6643_0[0]), .out(far_6_6643_1[0]));    relay_conn far_6_6643_1_b(.in(far_6_6643_0[1]), .out(far_6_6643_1[1]));
    assign layer_6[523] = ~far_6_6643_1[0]; 
    wire [1:0] far_6_6644_0;    relay_conn far_6_6644_0_a(.in(layer_5[25]), .out(far_6_6644_0[0]));    relay_conn far_6_6644_0_b(.in(layer_5[128]), .out(far_6_6644_0[1]));
    wire [1:0] far_6_6644_1;    relay_conn far_6_6644_1_a(.in(far_6_6644_0[0]), .out(far_6_6644_1[0]));    relay_conn far_6_6644_1_b(.in(far_6_6644_0[1]), .out(far_6_6644_1[1]));
    wire [1:0] far_6_6644_2;    relay_conn far_6_6644_2_a(.in(far_6_6644_1[0]), .out(far_6_6644_2[0]));    relay_conn far_6_6644_2_b(.in(far_6_6644_1[1]), .out(far_6_6644_2[1]));
    assign layer_6[524] = ~far_6_6644_2[0]; 
    assign layer_6[525] = layer_5[612]; 
    wire [1:0] far_6_6646_0;    relay_conn far_6_6646_0_a(.in(layer_5[985]), .out(far_6_6646_0[0]));    relay_conn far_6_6646_0_b(.in(layer_5[860]), .out(far_6_6646_0[1]));
    wire [1:0] far_6_6646_1;    relay_conn far_6_6646_1_a(.in(far_6_6646_0[0]), .out(far_6_6646_1[0]));    relay_conn far_6_6646_1_b(.in(far_6_6646_0[1]), .out(far_6_6646_1[1]));
    wire [1:0] far_6_6646_2;    relay_conn far_6_6646_2_a(.in(far_6_6646_1[0]), .out(far_6_6646_2[0]));    relay_conn far_6_6646_2_b(.in(far_6_6646_1[1]), .out(far_6_6646_2[1]));
    assign layer_6[526] = ~far_6_6646_2[0] | (far_6_6646_2[0] & far_6_6646_2[1]); 
    wire [1:0] far_6_6647_0;    relay_conn far_6_6647_0_a(.in(layer_5[689]), .out(far_6_6647_0[0]));    relay_conn far_6_6647_0_b(.in(layer_5[597]), .out(far_6_6647_0[1]));
    wire [1:0] far_6_6647_1;    relay_conn far_6_6647_1_a(.in(far_6_6647_0[0]), .out(far_6_6647_1[0]));    relay_conn far_6_6647_1_b(.in(far_6_6647_0[1]), .out(far_6_6647_1[1]));
    assign layer_6[527] = far_6_6647_1[0] & far_6_6647_1[1]; 
    wire [1:0] far_6_6648_0;    relay_conn far_6_6648_0_a(.in(layer_5[301]), .out(far_6_6648_0[0]));    relay_conn far_6_6648_0_b(.in(layer_5[222]), .out(far_6_6648_0[1]));
    wire [1:0] far_6_6648_1;    relay_conn far_6_6648_1_a(.in(far_6_6648_0[0]), .out(far_6_6648_1[0]));    relay_conn far_6_6648_1_b(.in(far_6_6648_0[1]), .out(far_6_6648_1[1]));
    assign layer_6[528] = far_6_6648_1[0] ^ far_6_6648_1[1]; 
    assign layer_6[529] = ~layer_5[460] | (layer_5[460] & layer_5[457]); 
    assign layer_6[530] = ~layer_5[39]; 
    wire [1:0] far_6_6651_0;    relay_conn far_6_6651_0_a(.in(layer_5[487]), .out(far_6_6651_0[0]));    relay_conn far_6_6651_0_b(.in(layer_5[538]), .out(far_6_6651_0[1]));
    assign layer_6[531] = ~(far_6_6651_0[0] | far_6_6651_0[1]); 
    wire [1:0] far_6_6652_0;    relay_conn far_6_6652_0_a(.in(layer_5[487]), .out(far_6_6652_0[0]));    relay_conn far_6_6652_0_b(.in(layer_5[527]), .out(far_6_6652_0[1]));
    assign layer_6[532] = ~far_6_6652_0[1] | (far_6_6652_0[0] & far_6_6652_0[1]); 
    assign layer_6[533] = layer_5[129]; 
    wire [1:0] far_6_6654_0;    relay_conn far_6_6654_0_a(.in(layer_5[574]), .out(far_6_6654_0[0]));    relay_conn far_6_6654_0_b(.in(layer_5[612]), .out(far_6_6654_0[1]));
    assign layer_6[534] = ~far_6_6654_0[0]; 
    wire [1:0] far_6_6655_0;    relay_conn far_6_6655_0_a(.in(layer_5[399]), .out(far_6_6655_0[0]));    relay_conn far_6_6655_0_b(.in(layer_5[274]), .out(far_6_6655_0[1]));
    wire [1:0] far_6_6655_1;    relay_conn far_6_6655_1_a(.in(far_6_6655_0[0]), .out(far_6_6655_1[0]));    relay_conn far_6_6655_1_b(.in(far_6_6655_0[1]), .out(far_6_6655_1[1]));
    wire [1:0] far_6_6655_2;    relay_conn far_6_6655_2_a(.in(far_6_6655_1[0]), .out(far_6_6655_2[0]));    relay_conn far_6_6655_2_b(.in(far_6_6655_1[1]), .out(far_6_6655_2[1]));
    assign layer_6[535] = ~far_6_6655_2[1] | (far_6_6655_2[0] & far_6_6655_2[1]); 
    assign layer_6[536] = ~(layer_5[57] & layer_5[26]); 
    wire [1:0] far_6_6657_0;    relay_conn far_6_6657_0_a(.in(layer_5[690]), .out(far_6_6657_0[0]));    relay_conn far_6_6657_0_b(.in(layer_5[593]), .out(far_6_6657_0[1]));
    wire [1:0] far_6_6657_1;    relay_conn far_6_6657_1_a(.in(far_6_6657_0[0]), .out(far_6_6657_1[0]));    relay_conn far_6_6657_1_b(.in(far_6_6657_0[1]), .out(far_6_6657_1[1]));
    wire [1:0] far_6_6657_2;    relay_conn far_6_6657_2_a(.in(far_6_6657_1[0]), .out(far_6_6657_2[0]));    relay_conn far_6_6657_2_b(.in(far_6_6657_1[1]), .out(far_6_6657_2[1]));
    assign layer_6[537] = ~far_6_6657_2[1] | (far_6_6657_2[0] & far_6_6657_2[1]); 
    wire [1:0] far_6_6658_0;    relay_conn far_6_6658_0_a(.in(layer_5[514]), .out(far_6_6658_0[0]));    relay_conn far_6_6658_0_b(.in(layer_5[550]), .out(far_6_6658_0[1]));
    assign layer_6[538] = far_6_6658_0[0]; 
    wire [1:0] far_6_6659_0;    relay_conn far_6_6659_0_a(.in(layer_5[300]), .out(far_6_6659_0[0]));    relay_conn far_6_6659_0_b(.in(layer_5[215]), .out(far_6_6659_0[1]));
    wire [1:0] far_6_6659_1;    relay_conn far_6_6659_1_a(.in(far_6_6659_0[0]), .out(far_6_6659_1[0]));    relay_conn far_6_6659_1_b(.in(far_6_6659_0[1]), .out(far_6_6659_1[1]));
    assign layer_6[539] = ~(far_6_6659_1[0] | far_6_6659_1[1]); 
    wire [1:0] far_6_6660_0;    relay_conn far_6_6660_0_a(.in(layer_5[571]), .out(far_6_6660_0[0]));    relay_conn far_6_6660_0_b(.in(layer_5[522]), .out(far_6_6660_0[1]));
    assign layer_6[540] = ~far_6_6660_0[1]; 
    wire [1:0] far_6_6661_0;    relay_conn far_6_6661_0_a(.in(layer_5[913]), .out(far_6_6661_0[0]));    relay_conn far_6_6661_0_b(.in(layer_5[977]), .out(far_6_6661_0[1]));
    wire [1:0] far_6_6661_1;    relay_conn far_6_6661_1_a(.in(far_6_6661_0[0]), .out(far_6_6661_1[0]));    relay_conn far_6_6661_1_b(.in(far_6_6661_0[1]), .out(far_6_6661_1[1]));
    assign layer_6[541] = far_6_6661_1[0] & far_6_6661_1[1]; 
    wire [1:0] far_6_6662_0;    relay_conn far_6_6662_0_a(.in(layer_5[668]), .out(far_6_6662_0[0]));    relay_conn far_6_6662_0_b(.in(layer_5[542]), .out(far_6_6662_0[1]));
    wire [1:0] far_6_6662_1;    relay_conn far_6_6662_1_a(.in(far_6_6662_0[0]), .out(far_6_6662_1[0]));    relay_conn far_6_6662_1_b(.in(far_6_6662_0[1]), .out(far_6_6662_1[1]));
    wire [1:0] far_6_6662_2;    relay_conn far_6_6662_2_a(.in(far_6_6662_1[0]), .out(far_6_6662_2[0]));    relay_conn far_6_6662_2_b(.in(far_6_6662_1[1]), .out(far_6_6662_2[1]));
    assign layer_6[542] = far_6_6662_2[1] & ~far_6_6662_2[0]; 
    wire [1:0] far_6_6663_0;    relay_conn far_6_6663_0_a(.in(layer_5[612]), .out(far_6_6663_0[0]));    relay_conn far_6_6663_0_b(.in(layer_5[722]), .out(far_6_6663_0[1]));
    wire [1:0] far_6_6663_1;    relay_conn far_6_6663_1_a(.in(far_6_6663_0[0]), .out(far_6_6663_1[0]));    relay_conn far_6_6663_1_b(.in(far_6_6663_0[1]), .out(far_6_6663_1[1]));
    wire [1:0] far_6_6663_2;    relay_conn far_6_6663_2_a(.in(far_6_6663_1[0]), .out(far_6_6663_2[0]));    relay_conn far_6_6663_2_b(.in(far_6_6663_1[1]), .out(far_6_6663_2[1]));
    assign layer_6[543] = far_6_6663_2[0] & ~far_6_6663_2[1]; 
    assign layer_6[544] = ~layer_5[172] | (layer_5[172] & layer_5[150]); 
    wire [1:0] far_6_6665_0;    relay_conn far_6_6665_0_a(.in(layer_5[619]), .out(far_6_6665_0[0]));    relay_conn far_6_6665_0_b(.in(layer_5[564]), .out(far_6_6665_0[1]));
    assign layer_6[545] = ~far_6_6665_0[1]; 
    wire [1:0] far_6_6666_0;    relay_conn far_6_6666_0_a(.in(layer_5[723]), .out(far_6_6666_0[0]));    relay_conn far_6_6666_0_b(.in(layer_5[781]), .out(far_6_6666_0[1]));
    assign layer_6[546] = ~(far_6_6666_0[0] | far_6_6666_0[1]); 
    wire [1:0] far_6_6667_0;    relay_conn far_6_6667_0_a(.in(layer_5[319]), .out(far_6_6667_0[0]));    relay_conn far_6_6667_0_b(.in(layer_5[253]), .out(far_6_6667_0[1]));
    wire [1:0] far_6_6667_1;    relay_conn far_6_6667_1_a(.in(far_6_6667_0[0]), .out(far_6_6667_1[0]));    relay_conn far_6_6667_1_b(.in(far_6_6667_0[1]), .out(far_6_6667_1[1]));
    assign layer_6[547] = far_6_6667_1[1]; 
    wire [1:0] far_6_6668_0;    relay_conn far_6_6668_0_a(.in(layer_5[147]), .out(far_6_6668_0[0]));    relay_conn far_6_6668_0_b(.in(layer_5[19]), .out(far_6_6668_0[1]));
    wire [1:0] far_6_6668_1;    relay_conn far_6_6668_1_a(.in(far_6_6668_0[0]), .out(far_6_6668_1[0]));    relay_conn far_6_6668_1_b(.in(far_6_6668_0[1]), .out(far_6_6668_1[1]));
    wire [1:0] far_6_6668_2;    relay_conn far_6_6668_2_a(.in(far_6_6668_1[0]), .out(far_6_6668_2[0]));    relay_conn far_6_6668_2_b(.in(far_6_6668_1[1]), .out(far_6_6668_2[1]));
    wire [1:0] far_6_6668_3;    relay_conn far_6_6668_3_a(.in(far_6_6668_2[0]), .out(far_6_6668_3[0]));    relay_conn far_6_6668_3_b(.in(far_6_6668_2[1]), .out(far_6_6668_3[1]));
    assign layer_6[548] = ~far_6_6668_3[0] | (far_6_6668_3[0] & far_6_6668_3[1]); 
    wire [1:0] far_6_6669_0;    relay_conn far_6_6669_0_a(.in(layer_5[437]), .out(far_6_6669_0[0]));    relay_conn far_6_6669_0_b(.in(layer_5[384]), .out(far_6_6669_0[1]));
    assign layer_6[549] = far_6_6669_0[1]; 
    wire [1:0] far_6_6670_0;    relay_conn far_6_6670_0_a(.in(layer_5[296]), .out(far_6_6670_0[0]));    relay_conn far_6_6670_0_b(.in(layer_5[422]), .out(far_6_6670_0[1]));
    wire [1:0] far_6_6670_1;    relay_conn far_6_6670_1_a(.in(far_6_6670_0[0]), .out(far_6_6670_1[0]));    relay_conn far_6_6670_1_b(.in(far_6_6670_0[1]), .out(far_6_6670_1[1]));
    wire [1:0] far_6_6670_2;    relay_conn far_6_6670_2_a(.in(far_6_6670_1[0]), .out(far_6_6670_2[0]));    relay_conn far_6_6670_2_b(.in(far_6_6670_1[1]), .out(far_6_6670_2[1]));
    assign layer_6[550] = ~far_6_6670_2[1] | (far_6_6670_2[0] & far_6_6670_2[1]); 
    wire [1:0] far_6_6671_0;    relay_conn far_6_6671_0_a(.in(layer_5[981]), .out(far_6_6671_0[0]));    relay_conn far_6_6671_0_b(.in(layer_5[857]), .out(far_6_6671_0[1]));
    wire [1:0] far_6_6671_1;    relay_conn far_6_6671_1_a(.in(far_6_6671_0[0]), .out(far_6_6671_1[0]));    relay_conn far_6_6671_1_b(.in(far_6_6671_0[1]), .out(far_6_6671_1[1]));
    wire [1:0] far_6_6671_2;    relay_conn far_6_6671_2_a(.in(far_6_6671_1[0]), .out(far_6_6671_2[0]));    relay_conn far_6_6671_2_b(.in(far_6_6671_1[1]), .out(far_6_6671_2[1]));
    assign layer_6[551] = far_6_6671_2[0] & ~far_6_6671_2[1]; 
    assign layer_6[552] = layer_5[886]; 
    wire [1:0] far_6_6673_0;    relay_conn far_6_6673_0_a(.in(layer_5[224]), .out(far_6_6673_0[0]));    relay_conn far_6_6673_0_b(.in(layer_5[148]), .out(far_6_6673_0[1]));
    wire [1:0] far_6_6673_1;    relay_conn far_6_6673_1_a(.in(far_6_6673_0[0]), .out(far_6_6673_1[0]));    relay_conn far_6_6673_1_b(.in(far_6_6673_0[1]), .out(far_6_6673_1[1]));
    assign layer_6[553] = ~far_6_6673_1[0]; 
    assign layer_6[554] = ~layer_5[786]; 
    assign layer_6[555] = layer_5[983] & ~layer_5[988]; 
    wire [1:0] far_6_6676_0;    relay_conn far_6_6676_0_a(.in(layer_5[512]), .out(far_6_6676_0[0]));    relay_conn far_6_6676_0_b(.in(layer_5[435]), .out(far_6_6676_0[1]));
    wire [1:0] far_6_6676_1;    relay_conn far_6_6676_1_a(.in(far_6_6676_0[0]), .out(far_6_6676_1[0]));    relay_conn far_6_6676_1_b(.in(far_6_6676_0[1]), .out(far_6_6676_1[1]));
    assign layer_6[556] = far_6_6676_1[1] & ~far_6_6676_1[0]; 
    wire [1:0] far_6_6677_0;    relay_conn far_6_6677_0_a(.in(layer_5[977]), .out(far_6_6677_0[0]));    relay_conn far_6_6677_0_b(.in(layer_5[876]), .out(far_6_6677_0[1]));
    wire [1:0] far_6_6677_1;    relay_conn far_6_6677_1_a(.in(far_6_6677_0[0]), .out(far_6_6677_1[0]));    relay_conn far_6_6677_1_b(.in(far_6_6677_0[1]), .out(far_6_6677_1[1]));
    wire [1:0] far_6_6677_2;    relay_conn far_6_6677_2_a(.in(far_6_6677_1[0]), .out(far_6_6677_2[0]));    relay_conn far_6_6677_2_b(.in(far_6_6677_1[1]), .out(far_6_6677_2[1]));
    assign layer_6[557] = far_6_6677_2[0]; 
    wire [1:0] far_6_6678_0;    relay_conn far_6_6678_0_a(.in(layer_5[664]), .out(far_6_6678_0[0]));    relay_conn far_6_6678_0_b(.in(layer_5[766]), .out(far_6_6678_0[1]));
    wire [1:0] far_6_6678_1;    relay_conn far_6_6678_1_a(.in(far_6_6678_0[0]), .out(far_6_6678_1[0]));    relay_conn far_6_6678_1_b(.in(far_6_6678_0[1]), .out(far_6_6678_1[1]));
    wire [1:0] far_6_6678_2;    relay_conn far_6_6678_2_a(.in(far_6_6678_1[0]), .out(far_6_6678_2[0]));    relay_conn far_6_6678_2_b(.in(far_6_6678_1[1]), .out(far_6_6678_2[1]));
    assign layer_6[558] = far_6_6678_2[0] | far_6_6678_2[1]; 
    wire [1:0] far_6_6679_0;    relay_conn far_6_6679_0_a(.in(layer_5[440]), .out(far_6_6679_0[0]));    relay_conn far_6_6679_0_b(.in(layer_5[363]), .out(far_6_6679_0[1]));
    wire [1:0] far_6_6679_1;    relay_conn far_6_6679_1_a(.in(far_6_6679_0[0]), .out(far_6_6679_1[0]));    relay_conn far_6_6679_1_b(.in(far_6_6679_0[1]), .out(far_6_6679_1[1]));
    assign layer_6[559] = far_6_6679_1[1] & ~far_6_6679_1[0]; 
    wire [1:0] far_6_6680_0;    relay_conn far_6_6680_0_a(.in(layer_5[938]), .out(far_6_6680_0[0]));    relay_conn far_6_6680_0_b(.in(layer_5[995]), .out(far_6_6680_0[1]));
    assign layer_6[560] = ~far_6_6680_0[1] | (far_6_6680_0[0] & far_6_6680_0[1]); 
    wire [1:0] far_6_6681_0;    relay_conn far_6_6681_0_a(.in(layer_5[751]), .out(far_6_6681_0[0]));    relay_conn far_6_6681_0_b(.in(layer_5[856]), .out(far_6_6681_0[1]));
    wire [1:0] far_6_6681_1;    relay_conn far_6_6681_1_a(.in(far_6_6681_0[0]), .out(far_6_6681_1[0]));    relay_conn far_6_6681_1_b(.in(far_6_6681_0[1]), .out(far_6_6681_1[1]));
    wire [1:0] far_6_6681_2;    relay_conn far_6_6681_2_a(.in(far_6_6681_1[0]), .out(far_6_6681_2[0]));    relay_conn far_6_6681_2_b(.in(far_6_6681_1[1]), .out(far_6_6681_2[1]));
    assign layer_6[561] = ~far_6_6681_2[1]; 
    wire [1:0] far_6_6682_0;    relay_conn far_6_6682_0_a(.in(layer_5[291]), .out(far_6_6682_0[0]));    relay_conn far_6_6682_0_b(.in(layer_5[368]), .out(far_6_6682_0[1]));
    wire [1:0] far_6_6682_1;    relay_conn far_6_6682_1_a(.in(far_6_6682_0[0]), .out(far_6_6682_1[0]));    relay_conn far_6_6682_1_b(.in(far_6_6682_0[1]), .out(far_6_6682_1[1]));
    assign layer_6[562] = ~(far_6_6682_1[0] ^ far_6_6682_1[1]); 
    assign layer_6[563] = layer_5[23] | layer_5[22]; 
    assign layer_6[564] = layer_5[522] & layer_5[516]; 
    assign layer_6[565] = ~layer_5[454] | (layer_5[423] & layer_5[454]); 
    assign layer_6[566] = ~(layer_5[26] | layer_5[57]); 
    wire [1:0] far_6_6687_0;    relay_conn far_6_6687_0_a(.in(layer_5[515]), .out(far_6_6687_0[0]));    relay_conn far_6_6687_0_b(.in(layer_5[465]), .out(far_6_6687_0[1]));
    assign layer_6[567] = ~far_6_6687_0[0] | (far_6_6687_0[0] & far_6_6687_0[1]); 
    wire [1:0] far_6_6688_0;    relay_conn far_6_6688_0_a(.in(layer_5[928]), .out(far_6_6688_0[0]));    relay_conn far_6_6688_0_b(.in(layer_5[834]), .out(far_6_6688_0[1]));
    wire [1:0] far_6_6688_1;    relay_conn far_6_6688_1_a(.in(far_6_6688_0[0]), .out(far_6_6688_1[0]));    relay_conn far_6_6688_1_b(.in(far_6_6688_0[1]), .out(far_6_6688_1[1]));
    assign layer_6[568] = far_6_6688_1[1] & ~far_6_6688_1[0]; 
    assign layer_6[569] = ~layer_5[1016]; 
    wire [1:0] far_6_6690_0;    relay_conn far_6_6690_0_a(.in(layer_5[296]), .out(far_6_6690_0[0]));    relay_conn far_6_6690_0_b(.in(layer_5[233]), .out(far_6_6690_0[1]));
    assign layer_6[570] = ~far_6_6690_0[1] | (far_6_6690_0[0] & far_6_6690_0[1]); 
    wire [1:0] far_6_6691_0;    relay_conn far_6_6691_0_a(.in(layer_5[289]), .out(far_6_6691_0[0]));    relay_conn far_6_6691_0_b(.in(layer_5[373]), .out(far_6_6691_0[1]));
    wire [1:0] far_6_6691_1;    relay_conn far_6_6691_1_a(.in(far_6_6691_0[0]), .out(far_6_6691_1[0]));    relay_conn far_6_6691_1_b(.in(far_6_6691_0[1]), .out(far_6_6691_1[1]));
    assign layer_6[571] = far_6_6691_1[0]; 
    wire [1:0] far_6_6692_0;    relay_conn far_6_6692_0_a(.in(layer_5[557]), .out(far_6_6692_0[0]));    relay_conn far_6_6692_0_b(.in(layer_5[509]), .out(far_6_6692_0[1]));
    assign layer_6[572] = ~far_6_6692_0[1]; 
    wire [1:0] far_6_6693_0;    relay_conn far_6_6693_0_a(.in(layer_5[684]), .out(far_6_6693_0[0]));    relay_conn far_6_6693_0_b(.in(layer_5[731]), .out(far_6_6693_0[1]));
    assign layer_6[573] = ~(far_6_6693_0[0] | far_6_6693_0[1]); 
    wire [1:0] far_6_6694_0;    relay_conn far_6_6694_0_a(.in(layer_5[425]), .out(far_6_6694_0[0]));    relay_conn far_6_6694_0_b(.in(layer_5[384]), .out(far_6_6694_0[1]));
    assign layer_6[574] = far_6_6694_0[1]; 
    wire [1:0] far_6_6695_0;    relay_conn far_6_6695_0_a(.in(layer_5[276]), .out(far_6_6695_0[0]));    relay_conn far_6_6695_0_b(.in(layer_5[400]), .out(far_6_6695_0[1]));
    wire [1:0] far_6_6695_1;    relay_conn far_6_6695_1_a(.in(far_6_6695_0[0]), .out(far_6_6695_1[0]));    relay_conn far_6_6695_1_b(.in(far_6_6695_0[1]), .out(far_6_6695_1[1]));
    wire [1:0] far_6_6695_2;    relay_conn far_6_6695_2_a(.in(far_6_6695_1[0]), .out(far_6_6695_2[0]));    relay_conn far_6_6695_2_b(.in(far_6_6695_1[1]), .out(far_6_6695_2[1]));
    assign layer_6[575] = ~(far_6_6695_2[0] | far_6_6695_2[1]); 
    wire [1:0] far_6_6696_0;    relay_conn far_6_6696_0_a(.in(layer_5[505]), .out(far_6_6696_0[0]));    relay_conn far_6_6696_0_b(.in(layer_5[424]), .out(far_6_6696_0[1]));
    wire [1:0] far_6_6696_1;    relay_conn far_6_6696_1_a(.in(far_6_6696_0[0]), .out(far_6_6696_1[0]));    relay_conn far_6_6696_1_b(.in(far_6_6696_0[1]), .out(far_6_6696_1[1]));
    assign layer_6[576] = far_6_6696_1[0] | far_6_6696_1[1]; 
    wire [1:0] far_6_6697_0;    relay_conn far_6_6697_0_a(.in(layer_5[28]), .out(far_6_6697_0[0]));    relay_conn far_6_6697_0_b(.in(layer_5[149]), .out(far_6_6697_0[1]));
    wire [1:0] far_6_6697_1;    relay_conn far_6_6697_1_a(.in(far_6_6697_0[0]), .out(far_6_6697_1[0]));    relay_conn far_6_6697_1_b(.in(far_6_6697_0[1]), .out(far_6_6697_1[1]));
    wire [1:0] far_6_6697_2;    relay_conn far_6_6697_2_a(.in(far_6_6697_1[0]), .out(far_6_6697_2[0]));    relay_conn far_6_6697_2_b(.in(far_6_6697_1[1]), .out(far_6_6697_2[1]));
    assign layer_6[577] = ~far_6_6697_2[0]; 
    wire [1:0] far_6_6698_0;    relay_conn far_6_6698_0_a(.in(layer_5[706]), .out(far_6_6698_0[0]));    relay_conn far_6_6698_0_b(.in(layer_5[827]), .out(far_6_6698_0[1]));
    wire [1:0] far_6_6698_1;    relay_conn far_6_6698_1_a(.in(far_6_6698_0[0]), .out(far_6_6698_1[0]));    relay_conn far_6_6698_1_b(.in(far_6_6698_0[1]), .out(far_6_6698_1[1]));
    wire [1:0] far_6_6698_2;    relay_conn far_6_6698_2_a(.in(far_6_6698_1[0]), .out(far_6_6698_2[0]));    relay_conn far_6_6698_2_b(.in(far_6_6698_1[1]), .out(far_6_6698_2[1]));
    assign layer_6[578] = ~far_6_6698_2[0]; 
    wire [1:0] far_6_6699_0;    relay_conn far_6_6699_0_a(.in(layer_5[180]), .out(far_6_6699_0[0]));    relay_conn far_6_6699_0_b(.in(layer_5[227]), .out(far_6_6699_0[1]));
    assign layer_6[579] = far_6_6699_0[0]; 
    wire [1:0] far_6_6700_0;    relay_conn far_6_6700_0_a(.in(layer_5[1019]), .out(far_6_6700_0[0]));    relay_conn far_6_6700_0_b(.in(layer_5[921]), .out(far_6_6700_0[1]));
    wire [1:0] far_6_6700_1;    relay_conn far_6_6700_1_a(.in(far_6_6700_0[0]), .out(far_6_6700_1[0]));    relay_conn far_6_6700_1_b(.in(far_6_6700_0[1]), .out(far_6_6700_1[1]));
    wire [1:0] far_6_6700_2;    relay_conn far_6_6700_2_a(.in(far_6_6700_1[0]), .out(far_6_6700_2[0]));    relay_conn far_6_6700_2_b(.in(far_6_6700_1[1]), .out(far_6_6700_2[1]));
    assign layer_6[580] = ~far_6_6700_2[0]; 
    assign layer_6[581] = layer_5[668]; 
    wire [1:0] far_6_6702_0;    relay_conn far_6_6702_0_a(.in(layer_5[225]), .out(far_6_6702_0[0]));    relay_conn far_6_6702_0_b(.in(layer_5[182]), .out(far_6_6702_0[1]));
    assign layer_6[582] = ~far_6_6702_0[1]; 
    assign layer_6[583] = layer_5[505]; 
    wire [1:0] far_6_6704_0;    relay_conn far_6_6704_0_a(.in(layer_5[164]), .out(far_6_6704_0[0]));    relay_conn far_6_6704_0_b(.in(layer_5[76]), .out(far_6_6704_0[1]));
    wire [1:0] far_6_6704_1;    relay_conn far_6_6704_1_a(.in(far_6_6704_0[0]), .out(far_6_6704_1[0]));    relay_conn far_6_6704_1_b(.in(far_6_6704_0[1]), .out(far_6_6704_1[1]));
    assign layer_6[584] = far_6_6704_1[0] & ~far_6_6704_1[1]; 
    wire [1:0] far_6_6705_0;    relay_conn far_6_6705_0_a(.in(layer_5[78]), .out(far_6_6705_0[0]));    relay_conn far_6_6705_0_b(.in(layer_5[127]), .out(far_6_6705_0[1]));
    assign layer_6[585] = ~far_6_6705_0[0]; 
    wire [1:0] far_6_6706_0;    relay_conn far_6_6706_0_a(.in(layer_5[762]), .out(far_6_6706_0[0]));    relay_conn far_6_6706_0_b(.in(layer_5[656]), .out(far_6_6706_0[1]));
    wire [1:0] far_6_6706_1;    relay_conn far_6_6706_1_a(.in(far_6_6706_0[0]), .out(far_6_6706_1[0]));    relay_conn far_6_6706_1_b(.in(far_6_6706_0[1]), .out(far_6_6706_1[1]));
    wire [1:0] far_6_6706_2;    relay_conn far_6_6706_2_a(.in(far_6_6706_1[0]), .out(far_6_6706_2[0]));    relay_conn far_6_6706_2_b(.in(far_6_6706_1[1]), .out(far_6_6706_2[1]));
    assign layer_6[586] = ~(far_6_6706_2[0] | far_6_6706_2[1]); 
    wire [1:0] far_6_6707_0;    relay_conn far_6_6707_0_a(.in(layer_5[360]), .out(far_6_6707_0[0]));    relay_conn far_6_6707_0_b(.in(layer_5[418]), .out(far_6_6707_0[1]));
    assign layer_6[587] = far_6_6707_0[0]; 
    assign layer_6[588] = ~layer_5[225] | (layer_5[225] & layer_5[222]); 
    wire [1:0] far_6_6709_0;    relay_conn far_6_6709_0_a(.in(layer_5[754]), .out(far_6_6709_0[0]));    relay_conn far_6_6709_0_b(.in(layer_5[643]), .out(far_6_6709_0[1]));
    wire [1:0] far_6_6709_1;    relay_conn far_6_6709_1_a(.in(far_6_6709_0[0]), .out(far_6_6709_1[0]));    relay_conn far_6_6709_1_b(.in(far_6_6709_0[1]), .out(far_6_6709_1[1]));
    wire [1:0] far_6_6709_2;    relay_conn far_6_6709_2_a(.in(far_6_6709_1[0]), .out(far_6_6709_2[0]));    relay_conn far_6_6709_2_b(.in(far_6_6709_1[1]), .out(far_6_6709_2[1]));
    assign layer_6[589] = ~(far_6_6709_2[0] & far_6_6709_2[1]); 
    wire [1:0] far_6_6710_0;    relay_conn far_6_6710_0_a(.in(layer_5[490]), .out(far_6_6710_0[0]));    relay_conn far_6_6710_0_b(.in(layer_5[369]), .out(far_6_6710_0[1]));
    wire [1:0] far_6_6710_1;    relay_conn far_6_6710_1_a(.in(far_6_6710_0[0]), .out(far_6_6710_1[0]));    relay_conn far_6_6710_1_b(.in(far_6_6710_0[1]), .out(far_6_6710_1[1]));
    wire [1:0] far_6_6710_2;    relay_conn far_6_6710_2_a(.in(far_6_6710_1[0]), .out(far_6_6710_2[0]));    relay_conn far_6_6710_2_b(.in(far_6_6710_1[1]), .out(far_6_6710_2[1]));
    assign layer_6[590] = far_6_6710_2[1]; 
    wire [1:0] far_6_6711_0;    relay_conn far_6_6711_0_a(.in(layer_5[436]), .out(far_6_6711_0[0]));    relay_conn far_6_6711_0_b(.in(layer_5[516]), .out(far_6_6711_0[1]));
    wire [1:0] far_6_6711_1;    relay_conn far_6_6711_1_a(.in(far_6_6711_0[0]), .out(far_6_6711_1[0]));    relay_conn far_6_6711_1_b(.in(far_6_6711_0[1]), .out(far_6_6711_1[1]));
    assign layer_6[591] = far_6_6711_1[0]; 
    assign layer_6[592] = layer_5[840] & ~layer_5[810]; 
    wire [1:0] far_6_6713_0;    relay_conn far_6_6713_0_a(.in(layer_5[256]), .out(far_6_6713_0[0]));    relay_conn far_6_6713_0_b(.in(layer_5[222]), .out(far_6_6713_0[1]));
    assign layer_6[593] = ~far_6_6713_0[1] | (far_6_6713_0[0] & far_6_6713_0[1]); 
    assign layer_6[594] = ~(layer_5[659] | layer_5[688]); 
    assign layer_6[595] = ~layer_5[865] | (layer_5[865] & layer_5[881]); 
    wire [1:0] far_6_6716_0;    relay_conn far_6_6716_0_a(.in(layer_5[424]), .out(far_6_6716_0[0]));    relay_conn far_6_6716_0_b(.in(layer_5[341]), .out(far_6_6716_0[1]));
    wire [1:0] far_6_6716_1;    relay_conn far_6_6716_1_a(.in(far_6_6716_0[0]), .out(far_6_6716_1[0]));    relay_conn far_6_6716_1_b(.in(far_6_6716_0[1]), .out(far_6_6716_1[1]));
    assign layer_6[596] = far_6_6716_1[0]; 
    wire [1:0] far_6_6717_0;    relay_conn far_6_6717_0_a(.in(layer_5[894]), .out(far_6_6717_0[0]));    relay_conn far_6_6717_0_b(.in(layer_5[830]), .out(far_6_6717_0[1]));
    wire [1:0] far_6_6717_1;    relay_conn far_6_6717_1_a(.in(far_6_6717_0[0]), .out(far_6_6717_1[0]));    relay_conn far_6_6717_1_b(.in(far_6_6717_0[1]), .out(far_6_6717_1[1]));
    assign layer_6[597] = far_6_6717_1[0] & far_6_6717_1[1]; 
    wire [1:0] far_6_6718_0;    relay_conn far_6_6718_0_a(.in(layer_5[52]), .out(far_6_6718_0[0]));    relay_conn far_6_6718_0_b(.in(layer_5[127]), .out(far_6_6718_0[1]));
    wire [1:0] far_6_6718_1;    relay_conn far_6_6718_1_a(.in(far_6_6718_0[0]), .out(far_6_6718_1[0]));    relay_conn far_6_6718_1_b(.in(far_6_6718_0[1]), .out(far_6_6718_1[1]));
    assign layer_6[598] = ~far_6_6718_1[1]; 
    wire [1:0] far_6_6719_0;    relay_conn far_6_6719_0_a(.in(layer_5[505]), .out(far_6_6719_0[0]));    relay_conn far_6_6719_0_b(.in(layer_5[613]), .out(far_6_6719_0[1]));
    wire [1:0] far_6_6719_1;    relay_conn far_6_6719_1_a(.in(far_6_6719_0[0]), .out(far_6_6719_1[0]));    relay_conn far_6_6719_1_b(.in(far_6_6719_0[1]), .out(far_6_6719_1[1]));
    wire [1:0] far_6_6719_2;    relay_conn far_6_6719_2_a(.in(far_6_6719_1[0]), .out(far_6_6719_2[0]));    relay_conn far_6_6719_2_b(.in(far_6_6719_1[1]), .out(far_6_6719_2[1]));
    assign layer_6[599] = far_6_6719_2[0]; 
    wire [1:0] far_6_6720_0;    relay_conn far_6_6720_0_a(.in(layer_5[740]), .out(far_6_6720_0[0]));    relay_conn far_6_6720_0_b(.in(layer_5[818]), .out(far_6_6720_0[1]));
    wire [1:0] far_6_6720_1;    relay_conn far_6_6720_1_a(.in(far_6_6720_0[0]), .out(far_6_6720_1[0]));    relay_conn far_6_6720_1_b(.in(far_6_6720_0[1]), .out(far_6_6720_1[1]));
    assign layer_6[600] = ~far_6_6720_1[0]; 
    wire [1:0] far_6_6721_0;    relay_conn far_6_6721_0_a(.in(layer_5[903]), .out(far_6_6721_0[0]));    relay_conn far_6_6721_0_b(.in(layer_5[971]), .out(far_6_6721_0[1]));
    wire [1:0] far_6_6721_1;    relay_conn far_6_6721_1_a(.in(far_6_6721_0[0]), .out(far_6_6721_1[0]));    relay_conn far_6_6721_1_b(.in(far_6_6721_0[1]), .out(far_6_6721_1[1]));
    assign layer_6[601] = far_6_6721_1[0]; 
    wire [1:0] far_6_6722_0;    relay_conn far_6_6722_0_a(.in(layer_5[406]), .out(far_6_6722_0[0]));    relay_conn far_6_6722_0_b(.in(layer_5[364]), .out(far_6_6722_0[1]));
    assign layer_6[602] = ~far_6_6722_0[1] | (far_6_6722_0[0] & far_6_6722_0[1]); 
    assign layer_6[603] = layer_5[308]; 
    wire [1:0] far_6_6724_0;    relay_conn far_6_6724_0_a(.in(layer_5[651]), .out(far_6_6724_0[0]));    relay_conn far_6_6724_0_b(.in(layer_5[715]), .out(far_6_6724_0[1]));
    wire [1:0] far_6_6724_1;    relay_conn far_6_6724_1_a(.in(far_6_6724_0[0]), .out(far_6_6724_1[0]));    relay_conn far_6_6724_1_b(.in(far_6_6724_0[1]), .out(far_6_6724_1[1]));
    assign layer_6[604] = ~far_6_6724_1[0]; 
    assign layer_6[605] = layer_5[250]; 
    assign layer_6[606] = layer_5[800] & layer_5[827]; 
    wire [1:0] far_6_6727_0;    relay_conn far_6_6727_0_a(.in(layer_5[879]), .out(far_6_6727_0[0]));    relay_conn far_6_6727_0_b(.in(layer_5[958]), .out(far_6_6727_0[1]));
    wire [1:0] far_6_6727_1;    relay_conn far_6_6727_1_a(.in(far_6_6727_0[0]), .out(far_6_6727_1[0]));    relay_conn far_6_6727_1_b(.in(far_6_6727_0[1]), .out(far_6_6727_1[1]));
    assign layer_6[607] = ~far_6_6727_1[1] | (far_6_6727_1[0] & far_6_6727_1[1]); 
    wire [1:0] far_6_6728_0;    relay_conn far_6_6728_0_a(.in(layer_5[925]), .out(far_6_6728_0[0]));    relay_conn far_6_6728_0_b(.in(layer_5[968]), .out(far_6_6728_0[1]));
    assign layer_6[608] = far_6_6728_0[0] & far_6_6728_0[1]; 
    wire [1:0] far_6_6729_0;    relay_conn far_6_6729_0_a(.in(layer_5[696]), .out(far_6_6729_0[0]));    relay_conn far_6_6729_0_b(.in(layer_5[772]), .out(far_6_6729_0[1]));
    wire [1:0] far_6_6729_1;    relay_conn far_6_6729_1_a(.in(far_6_6729_0[0]), .out(far_6_6729_1[0]));    relay_conn far_6_6729_1_b(.in(far_6_6729_0[1]), .out(far_6_6729_1[1]));
    assign layer_6[609] = ~(far_6_6729_1[0] | far_6_6729_1[1]); 
    wire [1:0] far_6_6730_0;    relay_conn far_6_6730_0_a(.in(layer_5[1001]), .out(far_6_6730_0[0]));    relay_conn far_6_6730_0_b(.in(layer_5[898]), .out(far_6_6730_0[1]));
    wire [1:0] far_6_6730_1;    relay_conn far_6_6730_1_a(.in(far_6_6730_0[0]), .out(far_6_6730_1[0]));    relay_conn far_6_6730_1_b(.in(far_6_6730_0[1]), .out(far_6_6730_1[1]));
    wire [1:0] far_6_6730_2;    relay_conn far_6_6730_2_a(.in(far_6_6730_1[0]), .out(far_6_6730_2[0]));    relay_conn far_6_6730_2_b(.in(far_6_6730_1[1]), .out(far_6_6730_2[1]));
    assign layer_6[610] = ~far_6_6730_2[0] | (far_6_6730_2[0] & far_6_6730_2[1]); 
    wire [1:0] far_6_6731_0;    relay_conn far_6_6731_0_a(.in(layer_5[426]), .out(far_6_6731_0[0]));    relay_conn far_6_6731_0_b(.in(layer_5[492]), .out(far_6_6731_0[1]));
    wire [1:0] far_6_6731_1;    relay_conn far_6_6731_1_a(.in(far_6_6731_0[0]), .out(far_6_6731_1[0]));    relay_conn far_6_6731_1_b(.in(far_6_6731_0[1]), .out(far_6_6731_1[1]));
    assign layer_6[611] = ~(far_6_6731_1[0] ^ far_6_6731_1[1]); 
    wire [1:0] far_6_6732_0;    relay_conn far_6_6732_0_a(.in(layer_5[258]), .out(far_6_6732_0[0]));    relay_conn far_6_6732_0_b(.in(layer_5[182]), .out(far_6_6732_0[1]));
    wire [1:0] far_6_6732_1;    relay_conn far_6_6732_1_a(.in(far_6_6732_0[0]), .out(far_6_6732_1[0]));    relay_conn far_6_6732_1_b(.in(far_6_6732_0[1]), .out(far_6_6732_1[1]));
    assign layer_6[612] = ~(far_6_6732_1[0] | far_6_6732_1[1]); 
    wire [1:0] far_6_6733_0;    relay_conn far_6_6733_0_a(.in(layer_5[950]), .out(far_6_6733_0[0]));    relay_conn far_6_6733_0_b(.in(layer_5[989]), .out(far_6_6733_0[1]));
    assign layer_6[613] = ~far_6_6733_0[0]; 
    assign layer_6[614] = layer_5[670] ^ layer_5[675]; 
    wire [1:0] far_6_6735_0;    relay_conn far_6_6735_0_a(.in(layer_5[167]), .out(far_6_6735_0[0]));    relay_conn far_6_6735_0_b(.in(layer_5[219]), .out(far_6_6735_0[1]));
    assign layer_6[615] = far_6_6735_0[1]; 
    wire [1:0] far_6_6736_0;    relay_conn far_6_6736_0_a(.in(layer_5[555]), .out(far_6_6736_0[0]));    relay_conn far_6_6736_0_b(.in(layer_5[500]), .out(far_6_6736_0[1]));
    assign layer_6[616] = ~(far_6_6736_0[0] & far_6_6736_0[1]); 
    wire [1:0] far_6_6737_0;    relay_conn far_6_6737_0_a(.in(layer_5[288]), .out(far_6_6737_0[0]));    relay_conn far_6_6737_0_b(.in(layer_5[396]), .out(far_6_6737_0[1]));
    wire [1:0] far_6_6737_1;    relay_conn far_6_6737_1_a(.in(far_6_6737_0[0]), .out(far_6_6737_1[0]));    relay_conn far_6_6737_1_b(.in(far_6_6737_0[1]), .out(far_6_6737_1[1]));
    wire [1:0] far_6_6737_2;    relay_conn far_6_6737_2_a(.in(far_6_6737_1[0]), .out(far_6_6737_2[0]));    relay_conn far_6_6737_2_b(.in(far_6_6737_1[1]), .out(far_6_6737_2[1]));
    assign layer_6[617] = ~far_6_6737_2[0] | (far_6_6737_2[0] & far_6_6737_2[1]); 
    assign layer_6[618] = ~(layer_5[1019] ^ layer_5[993]); 
    wire [1:0] far_6_6739_0;    relay_conn far_6_6739_0_a(.in(layer_5[233]), .out(far_6_6739_0[0]));    relay_conn far_6_6739_0_b(.in(layer_5[125]), .out(far_6_6739_0[1]));
    wire [1:0] far_6_6739_1;    relay_conn far_6_6739_1_a(.in(far_6_6739_0[0]), .out(far_6_6739_1[0]));    relay_conn far_6_6739_1_b(.in(far_6_6739_0[1]), .out(far_6_6739_1[1]));
    wire [1:0] far_6_6739_2;    relay_conn far_6_6739_2_a(.in(far_6_6739_1[0]), .out(far_6_6739_2[0]));    relay_conn far_6_6739_2_b(.in(far_6_6739_1[1]), .out(far_6_6739_2[1]));
    assign layer_6[619] = ~(far_6_6739_2[0] ^ far_6_6739_2[1]); 
    wire [1:0] far_6_6740_0;    relay_conn far_6_6740_0_a(.in(layer_5[260]), .out(far_6_6740_0[0]));    relay_conn far_6_6740_0_b(.in(layer_5[378]), .out(far_6_6740_0[1]));
    wire [1:0] far_6_6740_1;    relay_conn far_6_6740_1_a(.in(far_6_6740_0[0]), .out(far_6_6740_1[0]));    relay_conn far_6_6740_1_b(.in(far_6_6740_0[1]), .out(far_6_6740_1[1]));
    wire [1:0] far_6_6740_2;    relay_conn far_6_6740_2_a(.in(far_6_6740_1[0]), .out(far_6_6740_2[0]));    relay_conn far_6_6740_2_b(.in(far_6_6740_1[1]), .out(far_6_6740_2[1]));
    assign layer_6[620] = ~(far_6_6740_2[0] & far_6_6740_2[1]); 
    assign layer_6[621] = layer_5[574] & ~layer_5[556]; 
    wire [1:0] far_6_6742_0;    relay_conn far_6_6742_0_a(.in(layer_5[617]), .out(far_6_6742_0[0]));    relay_conn far_6_6742_0_b(.in(layer_5[653]), .out(far_6_6742_0[1]));
    assign layer_6[622] = ~far_6_6742_0[0] | (far_6_6742_0[0] & far_6_6742_0[1]); 
    wire [1:0] far_6_6743_0;    relay_conn far_6_6743_0_a(.in(layer_5[571]), .out(far_6_6743_0[0]));    relay_conn far_6_6743_0_b(.in(layer_5[513]), .out(far_6_6743_0[1]));
    assign layer_6[623] = far_6_6743_0[0] & far_6_6743_0[1]; 
    wire [1:0] far_6_6744_0;    relay_conn far_6_6744_0_a(.in(layer_5[846]), .out(far_6_6744_0[0]));    relay_conn far_6_6744_0_b(.in(layer_5[729]), .out(far_6_6744_0[1]));
    wire [1:0] far_6_6744_1;    relay_conn far_6_6744_1_a(.in(far_6_6744_0[0]), .out(far_6_6744_1[0]));    relay_conn far_6_6744_1_b(.in(far_6_6744_0[1]), .out(far_6_6744_1[1]));
    wire [1:0] far_6_6744_2;    relay_conn far_6_6744_2_a(.in(far_6_6744_1[0]), .out(far_6_6744_2[0]));    relay_conn far_6_6744_2_b(.in(far_6_6744_1[1]), .out(far_6_6744_2[1]));
    assign layer_6[624] = ~(far_6_6744_2[0] & far_6_6744_2[1]); 
    wire [1:0] far_6_6745_0;    relay_conn far_6_6745_0_a(.in(layer_5[932]), .out(far_6_6745_0[0]));    relay_conn far_6_6745_0_b(.in(layer_5[982]), .out(far_6_6745_0[1]));
    assign layer_6[625] = ~far_6_6745_0[0]; 
    wire [1:0] far_6_6746_0;    relay_conn far_6_6746_0_a(.in(layer_5[275]), .out(far_6_6746_0[0]));    relay_conn far_6_6746_0_b(.in(layer_5[308]), .out(far_6_6746_0[1]));
    assign layer_6[626] = far_6_6746_0[0] & ~far_6_6746_0[1]; 
    wire [1:0] far_6_6747_0;    relay_conn far_6_6747_0_a(.in(layer_5[30]), .out(far_6_6747_0[0]));    relay_conn far_6_6747_0_b(.in(layer_5[67]), .out(far_6_6747_0[1]));
    assign layer_6[627] = ~far_6_6747_0[0] | (far_6_6747_0[0] & far_6_6747_0[1]); 
    wire [1:0] far_6_6748_0;    relay_conn far_6_6748_0_a(.in(layer_5[136]), .out(far_6_6748_0[0]));    relay_conn far_6_6748_0_b(.in(layer_5[234]), .out(far_6_6748_0[1]));
    wire [1:0] far_6_6748_1;    relay_conn far_6_6748_1_a(.in(far_6_6748_0[0]), .out(far_6_6748_1[0]));    relay_conn far_6_6748_1_b(.in(far_6_6748_0[1]), .out(far_6_6748_1[1]));
    wire [1:0] far_6_6748_2;    relay_conn far_6_6748_2_a(.in(far_6_6748_1[0]), .out(far_6_6748_2[0]));    relay_conn far_6_6748_2_b(.in(far_6_6748_1[1]), .out(far_6_6748_2[1]));
    assign layer_6[628] = far_6_6748_2[0] & far_6_6748_2[1]; 
    wire [1:0] far_6_6749_0;    relay_conn far_6_6749_0_a(.in(layer_5[814]), .out(far_6_6749_0[0]));    relay_conn far_6_6749_0_b(.in(layer_5[741]), .out(far_6_6749_0[1]));
    wire [1:0] far_6_6749_1;    relay_conn far_6_6749_1_a(.in(far_6_6749_0[0]), .out(far_6_6749_1[0]));    relay_conn far_6_6749_1_b(.in(far_6_6749_0[1]), .out(far_6_6749_1[1]));
    assign layer_6[629] = ~far_6_6749_1[1]; 
    wire [1:0] far_6_6750_0;    relay_conn far_6_6750_0_a(.in(layer_5[781]), .out(far_6_6750_0[0]));    relay_conn far_6_6750_0_b(.in(layer_5[892]), .out(far_6_6750_0[1]));
    wire [1:0] far_6_6750_1;    relay_conn far_6_6750_1_a(.in(far_6_6750_0[0]), .out(far_6_6750_1[0]));    relay_conn far_6_6750_1_b(.in(far_6_6750_0[1]), .out(far_6_6750_1[1]));
    wire [1:0] far_6_6750_2;    relay_conn far_6_6750_2_a(.in(far_6_6750_1[0]), .out(far_6_6750_2[0]));    relay_conn far_6_6750_2_b(.in(far_6_6750_1[1]), .out(far_6_6750_2[1]));
    assign layer_6[630] = far_6_6750_2[0] | far_6_6750_2[1]; 
    wire [1:0] far_6_6751_0;    relay_conn far_6_6751_0_a(.in(layer_5[138]), .out(far_6_6751_0[0]));    relay_conn far_6_6751_0_b(.in(layer_5[31]), .out(far_6_6751_0[1]));
    wire [1:0] far_6_6751_1;    relay_conn far_6_6751_1_a(.in(far_6_6751_0[0]), .out(far_6_6751_1[0]));    relay_conn far_6_6751_1_b(.in(far_6_6751_0[1]), .out(far_6_6751_1[1]));
    wire [1:0] far_6_6751_2;    relay_conn far_6_6751_2_a(.in(far_6_6751_1[0]), .out(far_6_6751_2[0]));    relay_conn far_6_6751_2_b(.in(far_6_6751_1[1]), .out(far_6_6751_2[1]));
    assign layer_6[631] = far_6_6751_2[0] | far_6_6751_2[1]; 
    assign layer_6[632] = ~(layer_5[477] & layer_5[473]); 
    wire [1:0] far_6_6753_0;    relay_conn far_6_6753_0_a(.in(layer_5[87]), .out(far_6_6753_0[0]));    relay_conn far_6_6753_0_b(.in(layer_5[149]), .out(far_6_6753_0[1]));
    assign layer_6[633] = ~far_6_6753_0[0]; 
    wire [1:0] far_6_6754_0;    relay_conn far_6_6754_0_a(.in(layer_5[722]), .out(far_6_6754_0[0]));    relay_conn far_6_6754_0_b(.in(layer_5[845]), .out(far_6_6754_0[1]));
    wire [1:0] far_6_6754_1;    relay_conn far_6_6754_1_a(.in(far_6_6754_0[0]), .out(far_6_6754_1[0]));    relay_conn far_6_6754_1_b(.in(far_6_6754_0[1]), .out(far_6_6754_1[1]));
    wire [1:0] far_6_6754_2;    relay_conn far_6_6754_2_a(.in(far_6_6754_1[0]), .out(far_6_6754_2[0]));    relay_conn far_6_6754_2_b(.in(far_6_6754_1[1]), .out(far_6_6754_2[1]));
    assign layer_6[634] = far_6_6754_2[1]; 
    wire [1:0] far_6_6755_0;    relay_conn far_6_6755_0_a(.in(layer_5[889]), .out(far_6_6755_0[0]));    relay_conn far_6_6755_0_b(.in(layer_5[955]), .out(far_6_6755_0[1]));
    wire [1:0] far_6_6755_1;    relay_conn far_6_6755_1_a(.in(far_6_6755_0[0]), .out(far_6_6755_1[0]));    relay_conn far_6_6755_1_b(.in(far_6_6755_0[1]), .out(far_6_6755_1[1]));
    assign layer_6[635] = ~far_6_6755_1[0]; 
    wire [1:0] far_6_6756_0;    relay_conn far_6_6756_0_a(.in(layer_5[748]), .out(far_6_6756_0[0]));    relay_conn far_6_6756_0_b(.in(layer_5[847]), .out(far_6_6756_0[1]));
    wire [1:0] far_6_6756_1;    relay_conn far_6_6756_1_a(.in(far_6_6756_0[0]), .out(far_6_6756_1[0]));    relay_conn far_6_6756_1_b(.in(far_6_6756_0[1]), .out(far_6_6756_1[1]));
    wire [1:0] far_6_6756_2;    relay_conn far_6_6756_2_a(.in(far_6_6756_1[0]), .out(far_6_6756_2[0]));    relay_conn far_6_6756_2_b(.in(far_6_6756_1[1]), .out(far_6_6756_2[1]));
    assign layer_6[636] = ~far_6_6756_2[1] | (far_6_6756_2[0] & far_6_6756_2[1]); 
    assign layer_6[637] = layer_5[772] & ~layer_5[746]; 
    assign layer_6[638] = layer_5[834]; 
    assign layer_6[639] = layer_5[149]; 
    wire [1:0] far_6_6760_0;    relay_conn far_6_6760_0_a(.in(layer_5[7]), .out(far_6_6760_0[0]));    relay_conn far_6_6760_0_b(.in(layer_5[127]), .out(far_6_6760_0[1]));
    wire [1:0] far_6_6760_1;    relay_conn far_6_6760_1_a(.in(far_6_6760_0[0]), .out(far_6_6760_1[0]));    relay_conn far_6_6760_1_b(.in(far_6_6760_0[1]), .out(far_6_6760_1[1]));
    wire [1:0] far_6_6760_2;    relay_conn far_6_6760_2_a(.in(far_6_6760_1[0]), .out(far_6_6760_2[0]));    relay_conn far_6_6760_2_b(.in(far_6_6760_1[1]), .out(far_6_6760_2[1]));
    assign layer_6[640] = far_6_6760_2[0] & ~far_6_6760_2[1]; 
    assign layer_6[641] = layer_5[637] & ~layer_5[640]; 
    wire [1:0] far_6_6762_0;    relay_conn far_6_6762_0_a(.in(layer_5[795]), .out(far_6_6762_0[0]));    relay_conn far_6_6762_0_b(.in(layer_5[756]), .out(far_6_6762_0[1]));
    assign layer_6[642] = ~far_6_6762_0[0]; 
    wire [1:0] far_6_6763_0;    relay_conn far_6_6763_0_a(.in(layer_5[290]), .out(far_6_6763_0[0]));    relay_conn far_6_6763_0_b(.in(layer_5[183]), .out(far_6_6763_0[1]));
    wire [1:0] far_6_6763_1;    relay_conn far_6_6763_1_a(.in(far_6_6763_0[0]), .out(far_6_6763_1[0]));    relay_conn far_6_6763_1_b(.in(far_6_6763_0[1]), .out(far_6_6763_1[1]));
    wire [1:0] far_6_6763_2;    relay_conn far_6_6763_2_a(.in(far_6_6763_1[0]), .out(far_6_6763_2[0]));    relay_conn far_6_6763_2_b(.in(far_6_6763_1[1]), .out(far_6_6763_2[1]));
    assign layer_6[643] = ~far_6_6763_2[1]; 
    wire [1:0] far_6_6764_0;    relay_conn far_6_6764_0_a(.in(layer_5[487]), .out(far_6_6764_0[0]));    relay_conn far_6_6764_0_b(.in(layer_5[390]), .out(far_6_6764_0[1]));
    wire [1:0] far_6_6764_1;    relay_conn far_6_6764_1_a(.in(far_6_6764_0[0]), .out(far_6_6764_1[0]));    relay_conn far_6_6764_1_b(.in(far_6_6764_0[1]), .out(far_6_6764_1[1]));
    wire [1:0] far_6_6764_2;    relay_conn far_6_6764_2_a(.in(far_6_6764_1[0]), .out(far_6_6764_2[0]));    relay_conn far_6_6764_2_b(.in(far_6_6764_1[1]), .out(far_6_6764_2[1]));
    assign layer_6[644] = far_6_6764_2[0] ^ far_6_6764_2[1]; 
    wire [1:0] far_6_6765_0;    relay_conn far_6_6765_0_a(.in(layer_5[317]), .out(far_6_6765_0[0]));    relay_conn far_6_6765_0_b(.in(layer_5[215]), .out(far_6_6765_0[1]));
    wire [1:0] far_6_6765_1;    relay_conn far_6_6765_1_a(.in(far_6_6765_0[0]), .out(far_6_6765_1[0]));    relay_conn far_6_6765_1_b(.in(far_6_6765_0[1]), .out(far_6_6765_1[1]));
    wire [1:0] far_6_6765_2;    relay_conn far_6_6765_2_a(.in(far_6_6765_1[0]), .out(far_6_6765_2[0]));    relay_conn far_6_6765_2_b(.in(far_6_6765_1[1]), .out(far_6_6765_2[1]));
    assign layer_6[645] = ~far_6_6765_2[1] | (far_6_6765_2[0] & far_6_6765_2[1]); 
    wire [1:0] far_6_6766_0;    relay_conn far_6_6766_0_a(.in(layer_5[94]), .out(far_6_6766_0[0]));    relay_conn far_6_6766_0_b(.in(layer_5[44]), .out(far_6_6766_0[1]));
    assign layer_6[646] = ~far_6_6766_0[0]; 
    wire [1:0] far_6_6767_0;    relay_conn far_6_6767_0_a(.in(layer_5[725]), .out(far_6_6767_0[0]));    relay_conn far_6_6767_0_b(.in(layer_5[774]), .out(far_6_6767_0[1]));
    assign layer_6[647] = far_6_6767_0[0] & far_6_6767_0[1]; 
    wire [1:0] far_6_6768_0;    relay_conn far_6_6768_0_a(.in(layer_5[296]), .out(far_6_6768_0[0]));    relay_conn far_6_6768_0_b(.in(layer_5[357]), .out(far_6_6768_0[1]));
    assign layer_6[648] = far_6_6768_0[0] | far_6_6768_0[1]; 
    assign layer_6[649] = layer_5[83]; 
    wire [1:0] far_6_6770_0;    relay_conn far_6_6770_0_a(.in(layer_5[233]), .out(far_6_6770_0[0]));    relay_conn far_6_6770_0_b(.in(layer_5[273]), .out(far_6_6770_0[1]));
    assign layer_6[650] = ~far_6_6770_0[1]; 
    wire [1:0] far_6_6771_0;    relay_conn far_6_6771_0_a(.in(layer_5[538]), .out(far_6_6771_0[0]));    relay_conn far_6_6771_0_b(.in(layer_5[413]), .out(far_6_6771_0[1]));
    wire [1:0] far_6_6771_1;    relay_conn far_6_6771_1_a(.in(far_6_6771_0[0]), .out(far_6_6771_1[0]));    relay_conn far_6_6771_1_b(.in(far_6_6771_0[1]), .out(far_6_6771_1[1]));
    wire [1:0] far_6_6771_2;    relay_conn far_6_6771_2_a(.in(far_6_6771_1[0]), .out(far_6_6771_2[0]));    relay_conn far_6_6771_2_b(.in(far_6_6771_1[1]), .out(far_6_6771_2[1]));
    assign layer_6[651] = ~far_6_6771_2[1]; 
    wire [1:0] far_6_6772_0;    relay_conn far_6_6772_0_a(.in(layer_5[854]), .out(far_6_6772_0[0]));    relay_conn far_6_6772_0_b(.in(layer_5[738]), .out(far_6_6772_0[1]));
    wire [1:0] far_6_6772_1;    relay_conn far_6_6772_1_a(.in(far_6_6772_0[0]), .out(far_6_6772_1[0]));    relay_conn far_6_6772_1_b(.in(far_6_6772_0[1]), .out(far_6_6772_1[1]));
    wire [1:0] far_6_6772_2;    relay_conn far_6_6772_2_a(.in(far_6_6772_1[0]), .out(far_6_6772_2[0]));    relay_conn far_6_6772_2_b(.in(far_6_6772_1[1]), .out(far_6_6772_2[1]));
    assign layer_6[652] = ~far_6_6772_2[0]; 
    wire [1:0] far_6_6773_0;    relay_conn far_6_6773_0_a(.in(layer_5[480]), .out(far_6_6773_0[0]));    relay_conn far_6_6773_0_b(.in(layer_5[364]), .out(far_6_6773_0[1]));
    wire [1:0] far_6_6773_1;    relay_conn far_6_6773_1_a(.in(far_6_6773_0[0]), .out(far_6_6773_1[0]));    relay_conn far_6_6773_1_b(.in(far_6_6773_0[1]), .out(far_6_6773_1[1]));
    wire [1:0] far_6_6773_2;    relay_conn far_6_6773_2_a(.in(far_6_6773_1[0]), .out(far_6_6773_2[0]));    relay_conn far_6_6773_2_b(.in(far_6_6773_1[1]), .out(far_6_6773_2[1]));
    assign layer_6[653] = ~far_6_6773_2[0]; 
    wire [1:0] far_6_6774_0;    relay_conn far_6_6774_0_a(.in(layer_5[866]), .out(far_6_6774_0[0]));    relay_conn far_6_6774_0_b(.in(layer_5[817]), .out(far_6_6774_0[1]));
    assign layer_6[654] = far_6_6774_0[0]; 
    assign layer_6[655] = ~layer_5[596] | (layer_5[596] & layer_5[578]); 
    wire [1:0] far_6_6776_0;    relay_conn far_6_6776_0_a(.in(layer_5[620]), .out(far_6_6776_0[0]));    relay_conn far_6_6776_0_b(.in(layer_5[542]), .out(far_6_6776_0[1]));
    wire [1:0] far_6_6776_1;    relay_conn far_6_6776_1_a(.in(far_6_6776_0[0]), .out(far_6_6776_1[0]));    relay_conn far_6_6776_1_b(.in(far_6_6776_0[1]), .out(far_6_6776_1[1]));
    assign layer_6[656] = far_6_6776_1[1] & ~far_6_6776_1[0]; 
    wire [1:0] far_6_6777_0;    relay_conn far_6_6777_0_a(.in(layer_5[613]), .out(far_6_6777_0[0]));    relay_conn far_6_6777_0_b(.in(layer_5[527]), .out(far_6_6777_0[1]));
    wire [1:0] far_6_6777_1;    relay_conn far_6_6777_1_a(.in(far_6_6777_0[0]), .out(far_6_6777_1[0]));    relay_conn far_6_6777_1_b(.in(far_6_6777_0[1]), .out(far_6_6777_1[1]));
    assign layer_6[657] = ~(far_6_6777_1[0] ^ far_6_6777_1[1]); 
    wire [1:0] far_6_6778_0;    relay_conn far_6_6778_0_a(.in(layer_5[706]), .out(far_6_6778_0[0]));    relay_conn far_6_6778_0_b(.in(layer_5[617]), .out(far_6_6778_0[1]));
    wire [1:0] far_6_6778_1;    relay_conn far_6_6778_1_a(.in(far_6_6778_0[0]), .out(far_6_6778_1[0]));    relay_conn far_6_6778_1_b(.in(far_6_6778_0[1]), .out(far_6_6778_1[1]));
    assign layer_6[658] = far_6_6778_1[0]; 
    wire [1:0] far_6_6779_0;    relay_conn far_6_6779_0_a(.in(layer_5[1017]), .out(far_6_6779_0[0]));    relay_conn far_6_6779_0_b(.in(layer_5[985]), .out(far_6_6779_0[1]));
    assign layer_6[659] = far_6_6779_0[0] | far_6_6779_0[1]; 
    wire [1:0] far_6_6780_0;    relay_conn far_6_6780_0_a(.in(layer_5[236]), .out(far_6_6780_0[0]));    relay_conn far_6_6780_0_b(.in(layer_5[177]), .out(far_6_6780_0[1]));
    assign layer_6[660] = ~far_6_6780_0[1]; 
    wire [1:0] far_6_6781_0;    relay_conn far_6_6781_0_a(.in(layer_5[360]), .out(far_6_6781_0[0]));    relay_conn far_6_6781_0_b(.in(layer_5[468]), .out(far_6_6781_0[1]));
    wire [1:0] far_6_6781_1;    relay_conn far_6_6781_1_a(.in(far_6_6781_0[0]), .out(far_6_6781_1[0]));    relay_conn far_6_6781_1_b(.in(far_6_6781_0[1]), .out(far_6_6781_1[1]));
    wire [1:0] far_6_6781_2;    relay_conn far_6_6781_2_a(.in(far_6_6781_1[0]), .out(far_6_6781_2[0]));    relay_conn far_6_6781_2_b(.in(far_6_6781_1[1]), .out(far_6_6781_2[1]));
    assign layer_6[661] = ~(far_6_6781_2[0] & far_6_6781_2[1]); 
    wire [1:0] far_6_6782_0;    relay_conn far_6_6782_0_a(.in(layer_5[584]), .out(far_6_6782_0[0]));    relay_conn far_6_6782_0_b(.in(layer_5[668]), .out(far_6_6782_0[1]));
    wire [1:0] far_6_6782_1;    relay_conn far_6_6782_1_a(.in(far_6_6782_0[0]), .out(far_6_6782_1[0]));    relay_conn far_6_6782_1_b(.in(far_6_6782_0[1]), .out(far_6_6782_1[1]));
    assign layer_6[662] = ~(far_6_6782_1[0] ^ far_6_6782_1[1]); 
    assign layer_6[663] = ~(layer_5[63] & layer_5[79]); 
    wire [1:0] far_6_6784_0;    relay_conn far_6_6784_0_a(.in(layer_5[740]), .out(far_6_6784_0[0]));    relay_conn far_6_6784_0_b(.in(layer_5[692]), .out(far_6_6784_0[1]));
    assign layer_6[664] = far_6_6784_0[0] & far_6_6784_0[1]; 
    wire [1:0] far_6_6785_0;    relay_conn far_6_6785_0_a(.in(layer_5[430]), .out(far_6_6785_0[0]));    relay_conn far_6_6785_0_b(.in(layer_5[525]), .out(far_6_6785_0[1]));
    wire [1:0] far_6_6785_1;    relay_conn far_6_6785_1_a(.in(far_6_6785_0[0]), .out(far_6_6785_1[0]));    relay_conn far_6_6785_1_b(.in(far_6_6785_0[1]), .out(far_6_6785_1[1]));
    assign layer_6[665] = far_6_6785_1[1] & ~far_6_6785_1[0]; 
    assign layer_6[666] = layer_5[556]; 
    wire [1:0] far_6_6787_0;    relay_conn far_6_6787_0_a(.in(layer_5[7]), .out(far_6_6787_0[0]));    relay_conn far_6_6787_0_b(.in(layer_5[79]), .out(far_6_6787_0[1]));
    wire [1:0] far_6_6787_1;    relay_conn far_6_6787_1_a(.in(far_6_6787_0[0]), .out(far_6_6787_1[0]));    relay_conn far_6_6787_1_b(.in(far_6_6787_0[1]), .out(far_6_6787_1[1]));
    assign layer_6[667] = far_6_6787_1[1] & ~far_6_6787_1[0]; 
    assign layer_6[668] = layer_5[972] & layer_5[948]; 
    wire [1:0] far_6_6789_0;    relay_conn far_6_6789_0_a(.in(layer_5[328]), .out(far_6_6789_0[0]));    relay_conn far_6_6789_0_b(.in(layer_5[440]), .out(far_6_6789_0[1]));
    wire [1:0] far_6_6789_1;    relay_conn far_6_6789_1_a(.in(far_6_6789_0[0]), .out(far_6_6789_1[0]));    relay_conn far_6_6789_1_b(.in(far_6_6789_0[1]), .out(far_6_6789_1[1]));
    wire [1:0] far_6_6789_2;    relay_conn far_6_6789_2_a(.in(far_6_6789_1[0]), .out(far_6_6789_2[0]));    relay_conn far_6_6789_2_b(.in(far_6_6789_1[1]), .out(far_6_6789_2[1]));
    assign layer_6[669] = far_6_6789_2[0]; 
    wire [1:0] far_6_6790_0;    relay_conn far_6_6790_0_a(.in(layer_5[139]), .out(far_6_6790_0[0]));    relay_conn far_6_6790_0_b(.in(layer_5[216]), .out(far_6_6790_0[1]));
    wire [1:0] far_6_6790_1;    relay_conn far_6_6790_1_a(.in(far_6_6790_0[0]), .out(far_6_6790_1[0]));    relay_conn far_6_6790_1_b(.in(far_6_6790_0[1]), .out(far_6_6790_1[1]));
    assign layer_6[670] = ~far_6_6790_1[0] | (far_6_6790_1[0] & far_6_6790_1[1]); 
    wire [1:0] far_6_6791_0;    relay_conn far_6_6791_0_a(.in(layer_5[782]), .out(far_6_6791_0[0]));    relay_conn far_6_6791_0_b(.in(layer_5[876]), .out(far_6_6791_0[1]));
    wire [1:0] far_6_6791_1;    relay_conn far_6_6791_1_a(.in(far_6_6791_0[0]), .out(far_6_6791_1[0]));    relay_conn far_6_6791_1_b(.in(far_6_6791_0[1]), .out(far_6_6791_1[1]));
    assign layer_6[671] = far_6_6791_1[1] & ~far_6_6791_1[0]; 
    wire [1:0] far_6_6792_0;    relay_conn far_6_6792_0_a(.in(layer_5[743]), .out(far_6_6792_0[0]));    relay_conn far_6_6792_0_b(.in(layer_5[849]), .out(far_6_6792_0[1]));
    wire [1:0] far_6_6792_1;    relay_conn far_6_6792_1_a(.in(far_6_6792_0[0]), .out(far_6_6792_1[0]));    relay_conn far_6_6792_1_b(.in(far_6_6792_0[1]), .out(far_6_6792_1[1]));
    wire [1:0] far_6_6792_2;    relay_conn far_6_6792_2_a(.in(far_6_6792_1[0]), .out(far_6_6792_2[0]));    relay_conn far_6_6792_2_b(.in(far_6_6792_1[1]), .out(far_6_6792_2[1]));
    assign layer_6[672] = far_6_6792_2[0] ^ far_6_6792_2[1]; 
    wire [1:0] far_6_6793_0;    relay_conn far_6_6793_0_a(.in(layer_5[593]), .out(far_6_6793_0[0]));    relay_conn far_6_6793_0_b(.in(layer_5[630]), .out(far_6_6793_0[1]));
    assign layer_6[673] = far_6_6793_0[1]; 
    wire [1:0] far_6_6794_0;    relay_conn far_6_6794_0_a(.in(layer_5[731]), .out(far_6_6794_0[0]));    relay_conn far_6_6794_0_b(.in(layer_5[656]), .out(far_6_6794_0[1]));
    wire [1:0] far_6_6794_1;    relay_conn far_6_6794_1_a(.in(far_6_6794_0[0]), .out(far_6_6794_1[0]));    relay_conn far_6_6794_1_b(.in(far_6_6794_0[1]), .out(far_6_6794_1[1]));
    assign layer_6[674] = far_6_6794_1[0] & far_6_6794_1[1]; 
    wire [1:0] far_6_6795_0;    relay_conn far_6_6795_0_a(.in(layer_5[244]), .out(far_6_6795_0[0]));    relay_conn far_6_6795_0_b(.in(layer_5[283]), .out(far_6_6795_0[1]));
    assign layer_6[675] = ~far_6_6795_0[0] | (far_6_6795_0[0] & far_6_6795_0[1]); 
    assign layer_6[676] = layer_5[464] ^ layer_5[439]; 
    wire [1:0] far_6_6797_0;    relay_conn far_6_6797_0_a(.in(layer_5[314]), .out(far_6_6797_0[0]));    relay_conn far_6_6797_0_b(.in(layer_5[258]), .out(far_6_6797_0[1]));
    assign layer_6[677] = ~far_6_6797_0[1]; 
    wire [1:0] far_6_6798_0;    relay_conn far_6_6798_0_a(.in(layer_5[911]), .out(far_6_6798_0[0]));    relay_conn far_6_6798_0_b(.in(layer_5[943]), .out(far_6_6798_0[1]));
    assign layer_6[678] = ~far_6_6798_0[1] | (far_6_6798_0[0] & far_6_6798_0[1]); 
    wire [1:0] far_6_6799_0;    relay_conn far_6_6799_0_a(.in(layer_5[758]), .out(far_6_6799_0[0]));    relay_conn far_6_6799_0_b(.in(layer_5[653]), .out(far_6_6799_0[1]));
    wire [1:0] far_6_6799_1;    relay_conn far_6_6799_1_a(.in(far_6_6799_0[0]), .out(far_6_6799_1[0]));    relay_conn far_6_6799_1_b(.in(far_6_6799_0[1]), .out(far_6_6799_1[1]));
    wire [1:0] far_6_6799_2;    relay_conn far_6_6799_2_a(.in(far_6_6799_1[0]), .out(far_6_6799_2[0]));    relay_conn far_6_6799_2_b(.in(far_6_6799_1[1]), .out(far_6_6799_2[1]));
    assign layer_6[679] = far_6_6799_2[0] & far_6_6799_2[1]; 
    assign layer_6[680] = layer_5[94] & ~layer_5[87]; 
    assign layer_6[681] = ~layer_5[124]; 
    wire [1:0] far_6_6802_0;    relay_conn far_6_6802_0_a(.in(layer_5[885]), .out(far_6_6802_0[0]));    relay_conn far_6_6802_0_b(.in(layer_5[972]), .out(far_6_6802_0[1]));
    wire [1:0] far_6_6802_1;    relay_conn far_6_6802_1_a(.in(far_6_6802_0[0]), .out(far_6_6802_1[0]));    relay_conn far_6_6802_1_b(.in(far_6_6802_0[1]), .out(far_6_6802_1[1]));
    assign layer_6[682] = far_6_6802_1[0] | far_6_6802_1[1]; 
    wire [1:0] far_6_6803_0;    relay_conn far_6_6803_0_a(.in(layer_5[948]), .out(far_6_6803_0[0]));    relay_conn far_6_6803_0_b(.in(layer_5[1019]), .out(far_6_6803_0[1]));
    wire [1:0] far_6_6803_1;    relay_conn far_6_6803_1_a(.in(far_6_6803_0[0]), .out(far_6_6803_1[0]));    relay_conn far_6_6803_1_b(.in(far_6_6803_0[1]), .out(far_6_6803_1[1]));
    assign layer_6[683] = far_6_6803_1[0] & far_6_6803_1[1]; 
    wire [1:0] far_6_6804_0;    relay_conn far_6_6804_0_a(.in(layer_5[598]), .out(far_6_6804_0[0]));    relay_conn far_6_6804_0_b(.in(layer_5[710]), .out(far_6_6804_0[1]));
    wire [1:0] far_6_6804_1;    relay_conn far_6_6804_1_a(.in(far_6_6804_0[0]), .out(far_6_6804_1[0]));    relay_conn far_6_6804_1_b(.in(far_6_6804_0[1]), .out(far_6_6804_1[1]));
    wire [1:0] far_6_6804_2;    relay_conn far_6_6804_2_a(.in(far_6_6804_1[0]), .out(far_6_6804_2[0]));    relay_conn far_6_6804_2_b(.in(far_6_6804_1[1]), .out(far_6_6804_2[1]));
    assign layer_6[684] = ~far_6_6804_2[0]; 
    wire [1:0] far_6_6805_0;    relay_conn far_6_6805_0_a(.in(layer_5[96]), .out(far_6_6805_0[0]));    relay_conn far_6_6805_0_b(.in(layer_5[44]), .out(far_6_6805_0[1]));
    assign layer_6[685] = ~(far_6_6805_0[0] | far_6_6805_0[1]); 
    assign layer_6[686] = ~layer_5[263]; 
    wire [1:0] far_6_6807_0;    relay_conn far_6_6807_0_a(.in(layer_5[209]), .out(far_6_6807_0[0]));    relay_conn far_6_6807_0_b(.in(layer_5[290]), .out(far_6_6807_0[1]));
    wire [1:0] far_6_6807_1;    relay_conn far_6_6807_1_a(.in(far_6_6807_0[0]), .out(far_6_6807_1[0]));    relay_conn far_6_6807_1_b(.in(far_6_6807_0[1]), .out(far_6_6807_1[1]));
    assign layer_6[687] = far_6_6807_1[0]; 
    wire [1:0] far_6_6808_0;    relay_conn far_6_6808_0_a(.in(layer_5[857]), .out(far_6_6808_0[0]));    relay_conn far_6_6808_0_b(.in(layer_5[741]), .out(far_6_6808_0[1]));
    wire [1:0] far_6_6808_1;    relay_conn far_6_6808_1_a(.in(far_6_6808_0[0]), .out(far_6_6808_1[0]));    relay_conn far_6_6808_1_b(.in(far_6_6808_0[1]), .out(far_6_6808_1[1]));
    wire [1:0] far_6_6808_2;    relay_conn far_6_6808_2_a(.in(far_6_6808_1[0]), .out(far_6_6808_2[0]));    relay_conn far_6_6808_2_b(.in(far_6_6808_1[1]), .out(far_6_6808_2[1]));
    assign layer_6[688] = far_6_6808_2[1]; 
    assign layer_6[689] = ~(layer_5[758] & layer_5[773]); 
    wire [1:0] far_6_6810_0;    relay_conn far_6_6810_0_a(.in(layer_5[758]), .out(far_6_6810_0[0]));    relay_conn far_6_6810_0_b(.in(layer_5[865]), .out(far_6_6810_0[1]));
    wire [1:0] far_6_6810_1;    relay_conn far_6_6810_1_a(.in(far_6_6810_0[0]), .out(far_6_6810_1[0]));    relay_conn far_6_6810_1_b(.in(far_6_6810_0[1]), .out(far_6_6810_1[1]));
    wire [1:0] far_6_6810_2;    relay_conn far_6_6810_2_a(.in(far_6_6810_1[0]), .out(far_6_6810_2[0]));    relay_conn far_6_6810_2_b(.in(far_6_6810_1[1]), .out(far_6_6810_2[1]));
    assign layer_6[690] = ~(far_6_6810_2[0] & far_6_6810_2[1]); 
    wire [1:0] far_6_6811_0;    relay_conn far_6_6811_0_a(.in(layer_5[886]), .out(far_6_6811_0[0]));    relay_conn far_6_6811_0_b(.in(layer_5[765]), .out(far_6_6811_0[1]));
    wire [1:0] far_6_6811_1;    relay_conn far_6_6811_1_a(.in(far_6_6811_0[0]), .out(far_6_6811_1[0]));    relay_conn far_6_6811_1_b(.in(far_6_6811_0[1]), .out(far_6_6811_1[1]));
    wire [1:0] far_6_6811_2;    relay_conn far_6_6811_2_a(.in(far_6_6811_1[0]), .out(far_6_6811_2[0]));    relay_conn far_6_6811_2_b(.in(far_6_6811_1[1]), .out(far_6_6811_2[1]));
    assign layer_6[691] = far_6_6811_2[0] | far_6_6811_2[1]; 
    wire [1:0] far_6_6812_0;    relay_conn far_6_6812_0_a(.in(layer_5[783]), .out(far_6_6812_0[0]));    relay_conn far_6_6812_0_b(.in(layer_5[704]), .out(far_6_6812_0[1]));
    wire [1:0] far_6_6812_1;    relay_conn far_6_6812_1_a(.in(far_6_6812_0[0]), .out(far_6_6812_1[0]));    relay_conn far_6_6812_1_b(.in(far_6_6812_0[1]), .out(far_6_6812_1[1]));
    assign layer_6[692] = ~(far_6_6812_1[0] | far_6_6812_1[1]); 
    wire [1:0] far_6_6813_0;    relay_conn far_6_6813_0_a(.in(layer_5[746]), .out(far_6_6813_0[0]));    relay_conn far_6_6813_0_b(.in(layer_5[872]), .out(far_6_6813_0[1]));
    wire [1:0] far_6_6813_1;    relay_conn far_6_6813_1_a(.in(far_6_6813_0[0]), .out(far_6_6813_1[0]));    relay_conn far_6_6813_1_b(.in(far_6_6813_0[1]), .out(far_6_6813_1[1]));
    wire [1:0] far_6_6813_2;    relay_conn far_6_6813_2_a(.in(far_6_6813_1[0]), .out(far_6_6813_2[0]));    relay_conn far_6_6813_2_b(.in(far_6_6813_1[1]), .out(far_6_6813_2[1]));
    assign layer_6[693] = ~far_6_6813_2[0]; 
    wire [1:0] far_6_6814_0;    relay_conn far_6_6814_0_a(.in(layer_5[509]), .out(far_6_6814_0[0]));    relay_conn far_6_6814_0_b(.in(layer_5[611]), .out(far_6_6814_0[1]));
    wire [1:0] far_6_6814_1;    relay_conn far_6_6814_1_a(.in(far_6_6814_0[0]), .out(far_6_6814_1[0]));    relay_conn far_6_6814_1_b(.in(far_6_6814_0[1]), .out(far_6_6814_1[1]));
    wire [1:0] far_6_6814_2;    relay_conn far_6_6814_2_a(.in(far_6_6814_1[0]), .out(far_6_6814_2[0]));    relay_conn far_6_6814_2_b(.in(far_6_6814_1[1]), .out(far_6_6814_2[1]));
    assign layer_6[694] = far_6_6814_2[0] & ~far_6_6814_2[1]; 
    wire [1:0] far_6_6815_0;    relay_conn far_6_6815_0_a(.in(layer_5[934]), .out(far_6_6815_0[0]));    relay_conn far_6_6815_0_b(.in(layer_5[867]), .out(far_6_6815_0[1]));
    wire [1:0] far_6_6815_1;    relay_conn far_6_6815_1_a(.in(far_6_6815_0[0]), .out(far_6_6815_1[0]));    relay_conn far_6_6815_1_b(.in(far_6_6815_0[1]), .out(far_6_6815_1[1]));
    assign layer_6[695] = far_6_6815_1[0]; 
    wire [1:0] far_6_6816_0;    relay_conn far_6_6816_0_a(.in(layer_5[879]), .out(far_6_6816_0[0]));    relay_conn far_6_6816_0_b(.in(layer_5[840]), .out(far_6_6816_0[1]));
    assign layer_6[696] = far_6_6816_0[1] & ~far_6_6816_0[0]; 
    wire [1:0] far_6_6817_0;    relay_conn far_6_6817_0_a(.in(layer_5[550]), .out(far_6_6817_0[0]));    relay_conn far_6_6817_0_b(.in(layer_5[613]), .out(far_6_6817_0[1]));
    assign layer_6[697] = ~(far_6_6817_0[0] & far_6_6817_0[1]); 
    wire [1:0] far_6_6818_0;    relay_conn far_6_6818_0_a(.in(layer_5[760]), .out(far_6_6818_0[0]));    relay_conn far_6_6818_0_b(.in(layer_5[885]), .out(far_6_6818_0[1]));
    wire [1:0] far_6_6818_1;    relay_conn far_6_6818_1_a(.in(far_6_6818_0[0]), .out(far_6_6818_1[0]));    relay_conn far_6_6818_1_b(.in(far_6_6818_0[1]), .out(far_6_6818_1[1]));
    wire [1:0] far_6_6818_2;    relay_conn far_6_6818_2_a(.in(far_6_6818_1[0]), .out(far_6_6818_2[0]));    relay_conn far_6_6818_2_b(.in(far_6_6818_1[1]), .out(far_6_6818_2[1]));
    assign layer_6[698] = ~far_6_6818_2[0]; 
    wire [1:0] far_6_6819_0;    relay_conn far_6_6819_0_a(.in(layer_5[550]), .out(far_6_6819_0[0]));    relay_conn far_6_6819_0_b(.in(layer_5[439]), .out(far_6_6819_0[1]));
    wire [1:0] far_6_6819_1;    relay_conn far_6_6819_1_a(.in(far_6_6819_0[0]), .out(far_6_6819_1[0]));    relay_conn far_6_6819_1_b(.in(far_6_6819_0[1]), .out(far_6_6819_1[1]));
    wire [1:0] far_6_6819_2;    relay_conn far_6_6819_2_a(.in(far_6_6819_1[0]), .out(far_6_6819_2[0]));    relay_conn far_6_6819_2_b(.in(far_6_6819_1[1]), .out(far_6_6819_2[1]));
    assign layer_6[699] = ~far_6_6819_2[0]; 
    wire [1:0] far_6_6820_0;    relay_conn far_6_6820_0_a(.in(layer_5[147]), .out(far_6_6820_0[0]));    relay_conn far_6_6820_0_b(.in(layer_5[182]), .out(far_6_6820_0[1]));
    assign layer_6[700] = far_6_6820_0[0] | far_6_6820_0[1]; 
    assign layer_6[701] = ~(layer_5[825] ^ layer_5[814]); 
    assign layer_6[702] = ~layer_5[706]; 
    wire [1:0] far_6_6823_0;    relay_conn far_6_6823_0_a(.in(layer_5[250]), .out(far_6_6823_0[0]));    relay_conn far_6_6823_0_b(.in(layer_5[203]), .out(far_6_6823_0[1]));
    assign layer_6[703] = far_6_6823_0[0] & ~far_6_6823_0[1]; 
    wire [1:0] far_6_6824_0;    relay_conn far_6_6824_0_a(.in(layer_5[477]), .out(far_6_6824_0[0]));    relay_conn far_6_6824_0_b(.in(layer_5[596]), .out(far_6_6824_0[1]));
    wire [1:0] far_6_6824_1;    relay_conn far_6_6824_1_a(.in(far_6_6824_0[0]), .out(far_6_6824_1[0]));    relay_conn far_6_6824_1_b(.in(far_6_6824_0[1]), .out(far_6_6824_1[1]));
    wire [1:0] far_6_6824_2;    relay_conn far_6_6824_2_a(.in(far_6_6824_1[0]), .out(far_6_6824_2[0]));    relay_conn far_6_6824_2_b(.in(far_6_6824_1[1]), .out(far_6_6824_2[1]));
    assign layer_6[704] = far_6_6824_2[1]; 
    assign layer_6[705] = ~layer_5[480] | (layer_5[480] & layer_5[487]); 
    wire [1:0] far_6_6826_0;    relay_conn far_6_6826_0_a(.in(layer_5[512]), .out(far_6_6826_0[0]));    relay_conn far_6_6826_0_b(.in(layer_5[598]), .out(far_6_6826_0[1]));
    wire [1:0] far_6_6826_1;    relay_conn far_6_6826_1_a(.in(far_6_6826_0[0]), .out(far_6_6826_1[0]));    relay_conn far_6_6826_1_b(.in(far_6_6826_0[1]), .out(far_6_6826_1[1]));
    assign layer_6[706] = far_6_6826_1[0] | far_6_6826_1[1]; 
    wire [1:0] far_6_6827_0;    relay_conn far_6_6827_0_a(.in(layer_5[306]), .out(far_6_6827_0[0]));    relay_conn far_6_6827_0_b(.in(layer_5[219]), .out(far_6_6827_0[1]));
    wire [1:0] far_6_6827_1;    relay_conn far_6_6827_1_a(.in(far_6_6827_0[0]), .out(far_6_6827_1[0]));    relay_conn far_6_6827_1_b(.in(far_6_6827_0[1]), .out(far_6_6827_1[1]));
    assign layer_6[707] = far_6_6827_1[0] | far_6_6827_1[1]; 
    wire [1:0] far_6_6828_0;    relay_conn far_6_6828_0_a(.in(layer_5[351]), .out(far_6_6828_0[0]));    relay_conn far_6_6828_0_b(.in(layer_5[312]), .out(far_6_6828_0[1]));
    assign layer_6[708] = far_6_6828_0[1]; 
    assign layer_6[709] = ~(layer_5[519] ^ layer_5[501]); 
    wire [1:0] far_6_6830_0;    relay_conn far_6_6830_0_a(.in(layer_5[26]), .out(far_6_6830_0[0]));    relay_conn far_6_6830_0_b(.in(layer_5[150]), .out(far_6_6830_0[1]));
    wire [1:0] far_6_6830_1;    relay_conn far_6_6830_1_a(.in(far_6_6830_0[0]), .out(far_6_6830_1[0]));    relay_conn far_6_6830_1_b(.in(far_6_6830_0[1]), .out(far_6_6830_1[1]));
    wire [1:0] far_6_6830_2;    relay_conn far_6_6830_2_a(.in(far_6_6830_1[0]), .out(far_6_6830_2[0]));    relay_conn far_6_6830_2_b(.in(far_6_6830_1[1]), .out(far_6_6830_2[1]));
    assign layer_6[710] = far_6_6830_2[0] & ~far_6_6830_2[1]; 
    wire [1:0] far_6_6831_0;    relay_conn far_6_6831_0_a(.in(layer_5[222]), .out(far_6_6831_0[0]));    relay_conn far_6_6831_0_b(.in(layer_5[159]), .out(far_6_6831_0[1]));
    assign layer_6[711] = ~(far_6_6831_0[0] | far_6_6831_0[1]); 
    wire [1:0] far_6_6832_0;    relay_conn far_6_6832_0_a(.in(layer_5[527]), .out(far_6_6832_0[0]));    relay_conn far_6_6832_0_b(.in(layer_5[605]), .out(far_6_6832_0[1]));
    wire [1:0] far_6_6832_1;    relay_conn far_6_6832_1_a(.in(far_6_6832_0[0]), .out(far_6_6832_1[0]));    relay_conn far_6_6832_1_b(.in(far_6_6832_0[1]), .out(far_6_6832_1[1]));
    assign layer_6[712] = far_6_6832_1[0] & far_6_6832_1[1]; 
    assign layer_6[713] = ~(layer_5[424] ^ layer_5[445]); 
    wire [1:0] far_6_6834_0;    relay_conn far_6_6834_0_a(.in(layer_5[374]), .out(far_6_6834_0[0]));    relay_conn far_6_6834_0_b(.in(layer_5[424]), .out(far_6_6834_0[1]));
    assign layer_6[714] = far_6_6834_0[0] & ~far_6_6834_0[1]; 
    assign layer_6[715] = ~(layer_5[370] & layer_5[394]); 
    wire [1:0] far_6_6836_0;    relay_conn far_6_6836_0_a(.in(layer_5[405]), .out(far_6_6836_0[0]));    relay_conn far_6_6836_0_b(.in(layer_5[308]), .out(far_6_6836_0[1]));
    wire [1:0] far_6_6836_1;    relay_conn far_6_6836_1_a(.in(far_6_6836_0[0]), .out(far_6_6836_1[0]));    relay_conn far_6_6836_1_b(.in(far_6_6836_0[1]), .out(far_6_6836_1[1]));
    wire [1:0] far_6_6836_2;    relay_conn far_6_6836_2_a(.in(far_6_6836_1[0]), .out(far_6_6836_2[0]));    relay_conn far_6_6836_2_b(.in(far_6_6836_1[1]), .out(far_6_6836_2[1]));
    assign layer_6[716] = far_6_6836_2[0] | far_6_6836_2[1]; 
    assign layer_6[717] = layer_5[106] & ~layer_5[115]; 
    assign layer_6[718] = layer_5[751] & ~layer_5[746]; 
    assign layer_6[719] = layer_5[841] & layer_5[845]; 
    wire [1:0] far_6_6840_0;    relay_conn far_6_6840_0_a(.in(layer_5[3]), .out(far_6_6840_0[0]));    relay_conn far_6_6840_0_b(.in(layer_5[99]), .out(far_6_6840_0[1]));
    wire [1:0] far_6_6840_1;    relay_conn far_6_6840_1_a(.in(far_6_6840_0[0]), .out(far_6_6840_1[0]));    relay_conn far_6_6840_1_b(.in(far_6_6840_0[1]), .out(far_6_6840_1[1]));
    wire [1:0] far_6_6840_2;    relay_conn far_6_6840_2_a(.in(far_6_6840_1[0]), .out(far_6_6840_2[0]));    relay_conn far_6_6840_2_b(.in(far_6_6840_1[1]), .out(far_6_6840_2[1]));
    assign layer_6[720] = ~far_6_6840_2[0] | (far_6_6840_2[0] & far_6_6840_2[1]); 
    wire [1:0] far_6_6841_0;    relay_conn far_6_6841_0_a(.in(layer_5[471]), .out(far_6_6841_0[0]));    relay_conn far_6_6841_0_b(.in(layer_5[405]), .out(far_6_6841_0[1]));
    wire [1:0] far_6_6841_1;    relay_conn far_6_6841_1_a(.in(far_6_6841_0[0]), .out(far_6_6841_1[0]));    relay_conn far_6_6841_1_b(.in(far_6_6841_0[1]), .out(far_6_6841_1[1]));
    assign layer_6[721] = far_6_6841_1[0] | far_6_6841_1[1]; 
    wire [1:0] far_6_6842_0;    relay_conn far_6_6842_0_a(.in(layer_5[742]), .out(far_6_6842_0[0]));    relay_conn far_6_6842_0_b(.in(layer_5[651]), .out(far_6_6842_0[1]));
    wire [1:0] far_6_6842_1;    relay_conn far_6_6842_1_a(.in(far_6_6842_0[0]), .out(far_6_6842_1[0]));    relay_conn far_6_6842_1_b(.in(far_6_6842_0[1]), .out(far_6_6842_1[1]));
    assign layer_6[722] = far_6_6842_1[0] & ~far_6_6842_1[1]; 
    assign layer_6[723] = ~layer_5[25]; 
    wire [1:0] far_6_6844_0;    relay_conn far_6_6844_0_a(.in(layer_5[23]), .out(far_6_6844_0[0]));    relay_conn far_6_6844_0_b(.in(layer_5[95]), .out(far_6_6844_0[1]));
    wire [1:0] far_6_6844_1;    relay_conn far_6_6844_1_a(.in(far_6_6844_0[0]), .out(far_6_6844_1[0]));    relay_conn far_6_6844_1_b(.in(far_6_6844_0[1]), .out(far_6_6844_1[1]));
    assign layer_6[724] = ~far_6_6844_1[0]; 
    wire [1:0] far_6_6845_0;    relay_conn far_6_6845_0_a(.in(layer_5[559]), .out(far_6_6845_0[0]));    relay_conn far_6_6845_0_b(.in(layer_5[623]), .out(far_6_6845_0[1]));
    wire [1:0] far_6_6845_1;    relay_conn far_6_6845_1_a(.in(far_6_6845_0[0]), .out(far_6_6845_1[0]));    relay_conn far_6_6845_1_b(.in(far_6_6845_0[1]), .out(far_6_6845_1[1]));
    assign layer_6[725] = ~far_6_6845_1[1]; 
    assign layer_6[726] = ~layer_5[215]; 
    assign layer_6[727] = layer_5[795] & ~layer_5[802]; 
    wire [1:0] far_6_6848_0;    relay_conn far_6_6848_0_a(.in(layer_5[111]), .out(far_6_6848_0[0]));    relay_conn far_6_6848_0_b(.in(layer_5[78]), .out(far_6_6848_0[1]));
    assign layer_6[728] = ~far_6_6848_0[1]; 
    wire [1:0] far_6_6849_0;    relay_conn far_6_6849_0_a(.in(layer_5[432]), .out(far_6_6849_0[0]));    relay_conn far_6_6849_0_b(.in(layer_5[315]), .out(far_6_6849_0[1]));
    wire [1:0] far_6_6849_1;    relay_conn far_6_6849_1_a(.in(far_6_6849_0[0]), .out(far_6_6849_1[0]));    relay_conn far_6_6849_1_b(.in(far_6_6849_0[1]), .out(far_6_6849_1[1]));
    wire [1:0] far_6_6849_2;    relay_conn far_6_6849_2_a(.in(far_6_6849_1[0]), .out(far_6_6849_2[0]));    relay_conn far_6_6849_2_b(.in(far_6_6849_1[1]), .out(far_6_6849_2[1]));
    assign layer_6[729] = far_6_6849_2[0] | far_6_6849_2[1]; 
    wire [1:0] far_6_6850_0;    relay_conn far_6_6850_0_a(.in(layer_5[845]), .out(far_6_6850_0[0]));    relay_conn far_6_6850_0_b(.in(layer_5[910]), .out(far_6_6850_0[1]));
    wire [1:0] far_6_6850_1;    relay_conn far_6_6850_1_a(.in(far_6_6850_0[0]), .out(far_6_6850_1[0]));    relay_conn far_6_6850_1_b(.in(far_6_6850_0[1]), .out(far_6_6850_1[1]));
    assign layer_6[730] = far_6_6850_1[0]; 
    assign layer_6[731] = layer_5[261] & layer_5[274]; 
    wire [1:0] far_6_6852_0;    relay_conn far_6_6852_0_a(.in(layer_5[98]), .out(far_6_6852_0[0]));    relay_conn far_6_6852_0_b(.in(layer_5[190]), .out(far_6_6852_0[1]));
    wire [1:0] far_6_6852_1;    relay_conn far_6_6852_1_a(.in(far_6_6852_0[0]), .out(far_6_6852_1[0]));    relay_conn far_6_6852_1_b(.in(far_6_6852_0[1]), .out(far_6_6852_1[1]));
    assign layer_6[732] = ~(far_6_6852_1[0] ^ far_6_6852_1[1]); 
    assign layer_6[733] = layer_5[25] & layer_5[8]; 
    wire [1:0] far_6_6854_0;    relay_conn far_6_6854_0_a(.in(layer_5[258]), .out(far_6_6854_0[0]));    relay_conn far_6_6854_0_b(.in(layer_5[290]), .out(far_6_6854_0[1]));
    assign layer_6[734] = ~far_6_6854_0[0]; 
    assign layer_6[735] = ~layer_5[63] | (layer_5[63] & layer_5[92]); 
    assign layer_6[736] = layer_5[185] & ~layer_5[209]; 
    wire [1:0] far_6_6857_0;    relay_conn far_6_6857_0_a(.in(layer_5[791]), .out(far_6_6857_0[0]));    relay_conn far_6_6857_0_b(.in(layer_5[753]), .out(far_6_6857_0[1]));
    assign layer_6[737] = ~far_6_6857_0[1]; 
    wire [1:0] far_6_6858_0;    relay_conn far_6_6858_0_a(.in(layer_5[197]), .out(far_6_6858_0[0]));    relay_conn far_6_6858_0_b(.in(layer_5[139]), .out(far_6_6858_0[1]));
    assign layer_6[738] = ~far_6_6858_0[0] | (far_6_6858_0[0] & far_6_6858_0[1]); 
    wire [1:0] far_6_6859_0;    relay_conn far_6_6859_0_a(.in(layer_5[231]), .out(far_6_6859_0[0]));    relay_conn far_6_6859_0_b(.in(layer_5[185]), .out(far_6_6859_0[1]));
    assign layer_6[739] = ~far_6_6859_0[0]; 
    assign layer_6[740] = layer_5[186]; 
    wire [1:0] far_6_6861_0;    relay_conn far_6_6861_0_a(.in(layer_5[305]), .out(far_6_6861_0[0]));    relay_conn far_6_6861_0_b(.in(layer_5[430]), .out(far_6_6861_0[1]));
    wire [1:0] far_6_6861_1;    relay_conn far_6_6861_1_a(.in(far_6_6861_0[0]), .out(far_6_6861_1[0]));    relay_conn far_6_6861_1_b(.in(far_6_6861_0[1]), .out(far_6_6861_1[1]));
    wire [1:0] far_6_6861_2;    relay_conn far_6_6861_2_a(.in(far_6_6861_1[0]), .out(far_6_6861_2[0]));    relay_conn far_6_6861_2_b(.in(far_6_6861_1[1]), .out(far_6_6861_2[1]));
    assign layer_6[741] = ~far_6_6861_2[1]; 
    wire [1:0] far_6_6862_0;    relay_conn far_6_6862_0_a(.in(layer_5[483]), .out(far_6_6862_0[0]));    relay_conn far_6_6862_0_b(.in(layer_5[432]), .out(far_6_6862_0[1]));
    assign layer_6[742] = ~(far_6_6862_0[0] & far_6_6862_0[1]); 
    wire [1:0] far_6_6863_0;    relay_conn far_6_6863_0_a(.in(layer_5[368]), .out(far_6_6863_0[0]));    relay_conn far_6_6863_0_b(.in(layer_5[487]), .out(far_6_6863_0[1]));
    wire [1:0] far_6_6863_1;    relay_conn far_6_6863_1_a(.in(far_6_6863_0[0]), .out(far_6_6863_1[0]));    relay_conn far_6_6863_1_b(.in(far_6_6863_0[1]), .out(far_6_6863_1[1]));
    wire [1:0] far_6_6863_2;    relay_conn far_6_6863_2_a(.in(far_6_6863_1[0]), .out(far_6_6863_2[0]));    relay_conn far_6_6863_2_b(.in(far_6_6863_1[1]), .out(far_6_6863_2[1]));
    assign layer_6[743] = far_6_6863_2[0] | far_6_6863_2[1]; 
    wire [1:0] far_6_6864_0;    relay_conn far_6_6864_0_a(.in(layer_5[746]), .out(far_6_6864_0[0]));    relay_conn far_6_6864_0_b(.in(layer_5[847]), .out(far_6_6864_0[1]));
    wire [1:0] far_6_6864_1;    relay_conn far_6_6864_1_a(.in(far_6_6864_0[0]), .out(far_6_6864_1[0]));    relay_conn far_6_6864_1_b(.in(far_6_6864_0[1]), .out(far_6_6864_1[1]));
    wire [1:0] far_6_6864_2;    relay_conn far_6_6864_2_a(.in(far_6_6864_1[0]), .out(far_6_6864_2[0]));    relay_conn far_6_6864_2_b(.in(far_6_6864_1[1]), .out(far_6_6864_2[1]));
    assign layer_6[744] = ~far_6_6864_2[0]; 
    assign layer_6[745] = layer_5[217]; 
    wire [1:0] far_6_6866_0;    relay_conn far_6_6866_0_a(.in(layer_5[423]), .out(far_6_6866_0[0]));    relay_conn far_6_6866_0_b(.in(layer_5[498]), .out(far_6_6866_0[1]));
    wire [1:0] far_6_6866_1;    relay_conn far_6_6866_1_a(.in(far_6_6866_0[0]), .out(far_6_6866_1[0]));    relay_conn far_6_6866_1_b(.in(far_6_6866_0[1]), .out(far_6_6866_1[1]));
    assign layer_6[746] = far_6_6866_1[0]; 
    assign layer_6[747] = layer_5[851]; 
    assign layer_6[748] = ~(layer_5[795] | layer_5[797]); 
    wire [1:0] far_6_6869_0;    relay_conn far_6_6869_0_a(.in(layer_5[659]), .out(far_6_6869_0[0]));    relay_conn far_6_6869_0_b(.in(layer_5[774]), .out(far_6_6869_0[1]));
    wire [1:0] far_6_6869_1;    relay_conn far_6_6869_1_a(.in(far_6_6869_0[0]), .out(far_6_6869_1[0]));    relay_conn far_6_6869_1_b(.in(far_6_6869_0[1]), .out(far_6_6869_1[1]));
    wire [1:0] far_6_6869_2;    relay_conn far_6_6869_2_a(.in(far_6_6869_1[0]), .out(far_6_6869_2[0]));    relay_conn far_6_6869_2_b(.in(far_6_6869_1[1]), .out(far_6_6869_2[1]));
    assign layer_6[749] = ~far_6_6869_2[0]; 
    wire [1:0] far_6_6870_0;    relay_conn far_6_6870_0_a(.in(layer_5[565]), .out(far_6_6870_0[0]));    relay_conn far_6_6870_0_b(.in(layer_5[643]), .out(far_6_6870_0[1]));
    wire [1:0] far_6_6870_1;    relay_conn far_6_6870_1_a(.in(far_6_6870_0[0]), .out(far_6_6870_1[0]));    relay_conn far_6_6870_1_b(.in(far_6_6870_0[1]), .out(far_6_6870_1[1]));
    assign layer_6[750] = far_6_6870_1[0]; 
    wire [1:0] far_6_6871_0;    relay_conn far_6_6871_0_a(.in(layer_5[673]), .out(far_6_6871_0[0]));    relay_conn far_6_6871_0_b(.in(layer_5[722]), .out(far_6_6871_0[1]));
    assign layer_6[751] = ~far_6_6871_0[1]; 
    wire [1:0] far_6_6872_0;    relay_conn far_6_6872_0_a(.in(layer_5[439]), .out(far_6_6872_0[0]));    relay_conn far_6_6872_0_b(.in(layer_5[394]), .out(far_6_6872_0[1]));
    assign layer_6[752] = ~(far_6_6872_0[0] | far_6_6872_0[1]); 
    wire [1:0] far_6_6873_0;    relay_conn far_6_6873_0_a(.in(layer_5[231]), .out(far_6_6873_0[0]));    relay_conn far_6_6873_0_b(.in(layer_5[326]), .out(far_6_6873_0[1]));
    wire [1:0] far_6_6873_1;    relay_conn far_6_6873_1_a(.in(far_6_6873_0[0]), .out(far_6_6873_1[0]));    relay_conn far_6_6873_1_b(.in(far_6_6873_0[1]), .out(far_6_6873_1[1]));
    assign layer_6[753] = ~far_6_6873_1[1]; 
    wire [1:0] far_6_6874_0;    relay_conn far_6_6874_0_a(.in(layer_5[644]), .out(far_6_6874_0[0]));    relay_conn far_6_6874_0_b(.in(layer_5[752]), .out(far_6_6874_0[1]));
    wire [1:0] far_6_6874_1;    relay_conn far_6_6874_1_a(.in(far_6_6874_0[0]), .out(far_6_6874_1[0]));    relay_conn far_6_6874_1_b(.in(far_6_6874_0[1]), .out(far_6_6874_1[1]));
    wire [1:0] far_6_6874_2;    relay_conn far_6_6874_2_a(.in(far_6_6874_1[0]), .out(far_6_6874_2[0]));    relay_conn far_6_6874_2_b(.in(far_6_6874_1[1]), .out(far_6_6874_2[1]));
    assign layer_6[754] = ~far_6_6874_2[1] | (far_6_6874_2[0] & far_6_6874_2[1]); 
    wire [1:0] far_6_6875_0;    relay_conn far_6_6875_0_a(.in(layer_5[653]), .out(far_6_6875_0[0]));    relay_conn far_6_6875_0_b(.in(layer_5[769]), .out(far_6_6875_0[1]));
    wire [1:0] far_6_6875_1;    relay_conn far_6_6875_1_a(.in(far_6_6875_0[0]), .out(far_6_6875_1[0]));    relay_conn far_6_6875_1_b(.in(far_6_6875_0[1]), .out(far_6_6875_1[1]));
    wire [1:0] far_6_6875_2;    relay_conn far_6_6875_2_a(.in(far_6_6875_1[0]), .out(far_6_6875_2[0]));    relay_conn far_6_6875_2_b(.in(far_6_6875_1[1]), .out(far_6_6875_2[1]));
    assign layer_6[755] = ~(far_6_6875_2[0] | far_6_6875_2[1]); 
    wire [1:0] far_6_6876_0;    relay_conn far_6_6876_0_a(.in(layer_5[216]), .out(far_6_6876_0[0]));    relay_conn far_6_6876_0_b(.in(layer_5[309]), .out(far_6_6876_0[1]));
    wire [1:0] far_6_6876_1;    relay_conn far_6_6876_1_a(.in(far_6_6876_0[0]), .out(far_6_6876_1[0]));    relay_conn far_6_6876_1_b(.in(far_6_6876_0[1]), .out(far_6_6876_1[1]));
    assign layer_6[756] = ~far_6_6876_1[0]; 
    wire [1:0] far_6_6877_0;    relay_conn far_6_6877_0_a(.in(layer_5[206]), .out(far_6_6877_0[0]));    relay_conn far_6_6877_0_b(.in(layer_5[286]), .out(far_6_6877_0[1]));
    wire [1:0] far_6_6877_1;    relay_conn far_6_6877_1_a(.in(far_6_6877_0[0]), .out(far_6_6877_1[0]));    relay_conn far_6_6877_1_b(.in(far_6_6877_0[1]), .out(far_6_6877_1[1]));
    assign layer_6[757] = far_6_6877_1[0] & ~far_6_6877_1[1]; 
    assign layer_6[758] = ~layer_5[834]; 
    wire [1:0] far_6_6879_0;    relay_conn far_6_6879_0_a(.in(layer_5[489]), .out(far_6_6879_0[0]));    relay_conn far_6_6879_0_b(.in(layer_5[602]), .out(far_6_6879_0[1]));
    wire [1:0] far_6_6879_1;    relay_conn far_6_6879_1_a(.in(far_6_6879_0[0]), .out(far_6_6879_1[0]));    relay_conn far_6_6879_1_b(.in(far_6_6879_0[1]), .out(far_6_6879_1[1]));
    wire [1:0] far_6_6879_2;    relay_conn far_6_6879_2_a(.in(far_6_6879_1[0]), .out(far_6_6879_2[0]));    relay_conn far_6_6879_2_b(.in(far_6_6879_1[1]), .out(far_6_6879_2[1]));
    assign layer_6[759] = ~(far_6_6879_2[0] & far_6_6879_2[1]); 
    wire [1:0] far_6_6880_0;    relay_conn far_6_6880_0_a(.in(layer_5[152]), .out(far_6_6880_0[0]));    relay_conn far_6_6880_0_b(.in(layer_5[250]), .out(far_6_6880_0[1]));
    wire [1:0] far_6_6880_1;    relay_conn far_6_6880_1_a(.in(far_6_6880_0[0]), .out(far_6_6880_1[0]));    relay_conn far_6_6880_1_b(.in(far_6_6880_0[1]), .out(far_6_6880_1[1]));
    wire [1:0] far_6_6880_2;    relay_conn far_6_6880_2_a(.in(far_6_6880_1[0]), .out(far_6_6880_2[0]));    relay_conn far_6_6880_2_b(.in(far_6_6880_1[1]), .out(far_6_6880_2[1]));
    assign layer_6[760] = far_6_6880_2[1]; 
    wire [1:0] far_6_6881_0;    relay_conn far_6_6881_0_a(.in(layer_5[58]), .out(far_6_6881_0[0]));    relay_conn far_6_6881_0_b(.in(layer_5[106]), .out(far_6_6881_0[1]));
    assign layer_6[761] = far_6_6881_0[1] & ~far_6_6881_0[0]; 
    wire [1:0] far_6_6882_0;    relay_conn far_6_6882_0_a(.in(layer_5[203]), .out(far_6_6882_0[0]));    relay_conn far_6_6882_0_b(.in(layer_5[258]), .out(far_6_6882_0[1]));
    assign layer_6[762] = far_6_6882_0[0]; 
    assign layer_6[763] = layer_5[282]; 
    wire [1:0] far_6_6884_0;    relay_conn far_6_6884_0_a(.in(layer_5[845]), .out(far_6_6884_0[0]));    relay_conn far_6_6884_0_b(.in(layer_5[797]), .out(far_6_6884_0[1]));
    assign layer_6[764] = far_6_6884_0[0] & ~far_6_6884_0[1]; 
    wire [1:0] far_6_6885_0;    relay_conn far_6_6885_0_a(.in(layer_5[512]), .out(far_6_6885_0[0]));    relay_conn far_6_6885_0_b(.in(layer_5[578]), .out(far_6_6885_0[1]));
    wire [1:0] far_6_6885_1;    relay_conn far_6_6885_1_a(.in(far_6_6885_0[0]), .out(far_6_6885_1[0]));    relay_conn far_6_6885_1_b(.in(far_6_6885_0[1]), .out(far_6_6885_1[1]));
    assign layer_6[765] = ~far_6_6885_1[1] | (far_6_6885_1[0] & far_6_6885_1[1]); 
    wire [1:0] far_6_6886_0;    relay_conn far_6_6886_0_a(.in(layer_5[972]), .out(far_6_6886_0[0]));    relay_conn far_6_6886_0_b(.in(layer_5[875]), .out(far_6_6886_0[1]));
    wire [1:0] far_6_6886_1;    relay_conn far_6_6886_1_a(.in(far_6_6886_0[0]), .out(far_6_6886_1[0]));    relay_conn far_6_6886_1_b(.in(far_6_6886_0[1]), .out(far_6_6886_1[1]));
    wire [1:0] far_6_6886_2;    relay_conn far_6_6886_2_a(.in(far_6_6886_1[0]), .out(far_6_6886_2[0]));    relay_conn far_6_6886_2_b(.in(far_6_6886_1[1]), .out(far_6_6886_2[1]));
    assign layer_6[766] = far_6_6886_2[0]; 
    assign layer_6[767] = ~layer_5[639]; 
    assign layer_6[768] = ~(layer_5[121] | layer_5[152]); 
    wire [1:0] far_6_6889_0;    relay_conn far_6_6889_0_a(.in(layer_5[572]), .out(far_6_6889_0[0]));    relay_conn far_6_6889_0_b(.in(layer_5[688]), .out(far_6_6889_0[1]));
    wire [1:0] far_6_6889_1;    relay_conn far_6_6889_1_a(.in(far_6_6889_0[0]), .out(far_6_6889_1[0]));    relay_conn far_6_6889_1_b(.in(far_6_6889_0[1]), .out(far_6_6889_1[1]));
    wire [1:0] far_6_6889_2;    relay_conn far_6_6889_2_a(.in(far_6_6889_1[0]), .out(far_6_6889_2[0]));    relay_conn far_6_6889_2_b(.in(far_6_6889_1[1]), .out(far_6_6889_2[1]));
    assign layer_6[769] = ~(far_6_6889_2[0] & far_6_6889_2[1]); 
    wire [1:0] far_6_6890_0;    relay_conn far_6_6890_0_a(.in(layer_5[890]), .out(far_6_6890_0[0]));    relay_conn far_6_6890_0_b(.in(layer_5[765]), .out(far_6_6890_0[1]));
    wire [1:0] far_6_6890_1;    relay_conn far_6_6890_1_a(.in(far_6_6890_0[0]), .out(far_6_6890_1[0]));    relay_conn far_6_6890_1_b(.in(far_6_6890_0[1]), .out(far_6_6890_1[1]));
    wire [1:0] far_6_6890_2;    relay_conn far_6_6890_2_a(.in(far_6_6890_1[0]), .out(far_6_6890_2[0]));    relay_conn far_6_6890_2_b(.in(far_6_6890_1[1]), .out(far_6_6890_2[1]));
    assign layer_6[770] = far_6_6890_2[0] ^ far_6_6890_2[1]; 
    wire [1:0] far_6_6891_0;    relay_conn far_6_6891_0_a(.in(layer_5[157]), .out(far_6_6891_0[0]));    relay_conn far_6_6891_0_b(.in(layer_5[90]), .out(far_6_6891_0[1]));
    wire [1:0] far_6_6891_1;    relay_conn far_6_6891_1_a(.in(far_6_6891_0[0]), .out(far_6_6891_1[0]));    relay_conn far_6_6891_1_b(.in(far_6_6891_0[1]), .out(far_6_6891_1[1]));
    assign layer_6[771] = ~far_6_6891_1[1] | (far_6_6891_1[0] & far_6_6891_1[1]); 
    wire [1:0] far_6_6892_0;    relay_conn far_6_6892_0_a(.in(layer_5[230]), .out(far_6_6892_0[0]));    relay_conn far_6_6892_0_b(.in(layer_5[296]), .out(far_6_6892_0[1]));
    wire [1:0] far_6_6892_1;    relay_conn far_6_6892_1_a(.in(far_6_6892_0[0]), .out(far_6_6892_1[0]));    relay_conn far_6_6892_1_b(.in(far_6_6892_0[1]), .out(far_6_6892_1[1]));
    assign layer_6[772] = far_6_6892_1[0]; 
    wire [1:0] far_6_6893_0;    relay_conn far_6_6893_0_a(.in(layer_5[720]), .out(far_6_6893_0[0]));    relay_conn far_6_6893_0_b(.in(layer_5[653]), .out(far_6_6893_0[1]));
    wire [1:0] far_6_6893_1;    relay_conn far_6_6893_1_a(.in(far_6_6893_0[0]), .out(far_6_6893_1[0]));    relay_conn far_6_6893_1_b(.in(far_6_6893_0[1]), .out(far_6_6893_1[1]));
    assign layer_6[773] = far_6_6893_1[0] & ~far_6_6893_1[1]; 
    wire [1:0] far_6_6894_0;    relay_conn far_6_6894_0_a(.in(layer_5[939]), .out(far_6_6894_0[0]));    relay_conn far_6_6894_0_b(.in(layer_5[840]), .out(far_6_6894_0[1]));
    wire [1:0] far_6_6894_1;    relay_conn far_6_6894_1_a(.in(far_6_6894_0[0]), .out(far_6_6894_1[0]));    relay_conn far_6_6894_1_b(.in(far_6_6894_0[1]), .out(far_6_6894_1[1]));
    wire [1:0] far_6_6894_2;    relay_conn far_6_6894_2_a(.in(far_6_6894_1[0]), .out(far_6_6894_2[0]));    relay_conn far_6_6894_2_b(.in(far_6_6894_1[1]), .out(far_6_6894_2[1]));
    assign layer_6[774] = far_6_6894_2[0] ^ far_6_6894_2[1]; 
    wire [1:0] far_6_6895_0;    relay_conn far_6_6895_0_a(.in(layer_5[394]), .out(far_6_6895_0[0]));    relay_conn far_6_6895_0_b(.in(layer_5[431]), .out(far_6_6895_0[1]));
    assign layer_6[775] = ~far_6_6895_0[0]; 
    wire [1:0] far_6_6896_0;    relay_conn far_6_6896_0_a(.in(layer_5[122]), .out(far_6_6896_0[0]));    relay_conn far_6_6896_0_b(.in(layer_5[209]), .out(far_6_6896_0[1]));
    wire [1:0] far_6_6896_1;    relay_conn far_6_6896_1_a(.in(far_6_6896_0[0]), .out(far_6_6896_1[0]));    relay_conn far_6_6896_1_b(.in(far_6_6896_0[1]), .out(far_6_6896_1[1]));
    assign layer_6[776] = ~far_6_6896_1[1] | (far_6_6896_1[0] & far_6_6896_1[1]); 
    wire [1:0] far_6_6897_0;    relay_conn far_6_6897_0_a(.in(layer_5[470]), .out(far_6_6897_0[0]));    relay_conn far_6_6897_0_b(.in(layer_5[555]), .out(far_6_6897_0[1]));
    wire [1:0] far_6_6897_1;    relay_conn far_6_6897_1_a(.in(far_6_6897_0[0]), .out(far_6_6897_1[0]));    relay_conn far_6_6897_1_b(.in(far_6_6897_0[1]), .out(far_6_6897_1[1]));
    assign layer_6[777] = ~(far_6_6897_1[0] & far_6_6897_1[1]); 
    wire [1:0] far_6_6898_0;    relay_conn far_6_6898_0_a(.in(layer_5[104]), .out(far_6_6898_0[0]));    relay_conn far_6_6898_0_b(.in(layer_5[69]), .out(far_6_6898_0[1]));
    assign layer_6[778] = far_6_6898_0[1] & ~far_6_6898_0[0]; 
    wire [1:0] far_6_6899_0;    relay_conn far_6_6899_0_a(.in(layer_5[393]), .out(far_6_6899_0[0]));    relay_conn far_6_6899_0_b(.in(layer_5[275]), .out(far_6_6899_0[1]));
    wire [1:0] far_6_6899_1;    relay_conn far_6_6899_1_a(.in(far_6_6899_0[0]), .out(far_6_6899_1[0]));    relay_conn far_6_6899_1_b(.in(far_6_6899_0[1]), .out(far_6_6899_1[1]));
    wire [1:0] far_6_6899_2;    relay_conn far_6_6899_2_a(.in(far_6_6899_1[0]), .out(far_6_6899_2[0]));    relay_conn far_6_6899_2_b(.in(far_6_6899_1[1]), .out(far_6_6899_2[1]));
    assign layer_6[779] = ~far_6_6899_2[0]; 
    wire [1:0] far_6_6900_0;    relay_conn far_6_6900_0_a(.in(layer_5[832]), .out(far_6_6900_0[0]));    relay_conn far_6_6900_0_b(.in(layer_5[761]), .out(far_6_6900_0[1]));
    wire [1:0] far_6_6900_1;    relay_conn far_6_6900_1_a(.in(far_6_6900_0[0]), .out(far_6_6900_1[0]));    relay_conn far_6_6900_1_b(.in(far_6_6900_0[1]), .out(far_6_6900_1[1]));
    assign layer_6[780] = far_6_6900_1[0] & far_6_6900_1[1]; 
    wire [1:0] far_6_6901_0;    relay_conn far_6_6901_0_a(.in(layer_5[452]), .out(far_6_6901_0[0]));    relay_conn far_6_6901_0_b(.in(layer_5[515]), .out(far_6_6901_0[1]));
    assign layer_6[781] = ~far_6_6901_0[0] | (far_6_6901_0[0] & far_6_6901_0[1]); 
    assign layer_6[782] = ~(layer_5[925] | layer_5[956]); 
    assign layer_6[783] = layer_5[161] & layer_5[147]; 
    wire [1:0] far_6_6904_0;    relay_conn far_6_6904_0_a(.in(layer_5[69]), .out(far_6_6904_0[0]));    relay_conn far_6_6904_0_b(.in(layer_5[193]), .out(far_6_6904_0[1]));
    wire [1:0] far_6_6904_1;    relay_conn far_6_6904_1_a(.in(far_6_6904_0[0]), .out(far_6_6904_1[0]));    relay_conn far_6_6904_1_b(.in(far_6_6904_0[1]), .out(far_6_6904_1[1]));
    wire [1:0] far_6_6904_2;    relay_conn far_6_6904_2_a(.in(far_6_6904_1[0]), .out(far_6_6904_2[0]));    relay_conn far_6_6904_2_b(.in(far_6_6904_1[1]), .out(far_6_6904_2[1]));
    assign layer_6[784] = ~far_6_6904_2[1] | (far_6_6904_2[0] & far_6_6904_2[1]); 
    wire [1:0] far_6_6905_0;    relay_conn far_6_6905_0_a(.in(layer_5[685]), .out(far_6_6905_0[0]));    relay_conn far_6_6905_0_b(.in(layer_5[761]), .out(far_6_6905_0[1]));
    wire [1:0] far_6_6905_1;    relay_conn far_6_6905_1_a(.in(far_6_6905_0[0]), .out(far_6_6905_1[0]));    relay_conn far_6_6905_1_b(.in(far_6_6905_0[1]), .out(far_6_6905_1[1]));
    assign layer_6[785] = ~far_6_6905_1[1] | (far_6_6905_1[0] & far_6_6905_1[1]); 
    wire [1:0] far_6_6906_0;    relay_conn far_6_6906_0_a(.in(layer_5[228]), .out(far_6_6906_0[0]));    relay_conn far_6_6906_0_b(.in(layer_5[311]), .out(far_6_6906_0[1]));
    wire [1:0] far_6_6906_1;    relay_conn far_6_6906_1_a(.in(far_6_6906_0[0]), .out(far_6_6906_1[0]));    relay_conn far_6_6906_1_b(.in(far_6_6906_0[1]), .out(far_6_6906_1[1]));
    assign layer_6[786] = far_6_6906_1[0] | far_6_6906_1[1]; 
    wire [1:0] far_6_6907_0;    relay_conn far_6_6907_0_a(.in(layer_5[875]), .out(far_6_6907_0[0]));    relay_conn far_6_6907_0_b(.in(layer_5[837]), .out(far_6_6907_0[1]));
    assign layer_6[787] = ~far_6_6907_0[1] | (far_6_6907_0[0] & far_6_6907_0[1]); 
    wire [1:0] far_6_6908_0;    relay_conn far_6_6908_0_a(.in(layer_5[39]), .out(far_6_6908_0[0]));    relay_conn far_6_6908_0_b(.in(layer_5[3]), .out(far_6_6908_0[1]));
    assign layer_6[788] = far_6_6908_0[1]; 
    assign layer_6[789] = layer_5[746] & ~layer_5[774]; 
    wire [1:0] far_6_6910_0;    relay_conn far_6_6910_0_a(.in(layer_5[51]), .out(far_6_6910_0[0]));    relay_conn far_6_6910_0_b(.in(layer_5[11]), .out(far_6_6910_0[1]));
    assign layer_6[790] = ~far_6_6910_0[0]; 
    wire [1:0] far_6_6911_0;    relay_conn far_6_6911_0_a(.in(layer_5[813]), .out(far_6_6911_0[0]));    relay_conn far_6_6911_0_b(.in(layer_5[919]), .out(far_6_6911_0[1]));
    wire [1:0] far_6_6911_1;    relay_conn far_6_6911_1_a(.in(far_6_6911_0[0]), .out(far_6_6911_1[0]));    relay_conn far_6_6911_1_b(.in(far_6_6911_0[1]), .out(far_6_6911_1[1]));
    wire [1:0] far_6_6911_2;    relay_conn far_6_6911_2_a(.in(far_6_6911_1[0]), .out(far_6_6911_2[0]));    relay_conn far_6_6911_2_b(.in(far_6_6911_1[1]), .out(far_6_6911_2[1]));
    assign layer_6[791] = far_6_6911_2[0]; 
    wire [1:0] far_6_6912_0;    relay_conn far_6_6912_0_a(.in(layer_5[437]), .out(far_6_6912_0[0]));    relay_conn far_6_6912_0_b(.in(layer_5[328]), .out(far_6_6912_0[1]));
    wire [1:0] far_6_6912_1;    relay_conn far_6_6912_1_a(.in(far_6_6912_0[0]), .out(far_6_6912_1[0]));    relay_conn far_6_6912_1_b(.in(far_6_6912_0[1]), .out(far_6_6912_1[1]));
    wire [1:0] far_6_6912_2;    relay_conn far_6_6912_2_a(.in(far_6_6912_1[0]), .out(far_6_6912_2[0]));    relay_conn far_6_6912_2_b(.in(far_6_6912_1[1]), .out(far_6_6912_2[1]));
    assign layer_6[792] = ~far_6_6912_2[0]; 
    assign layer_6[793] = ~(layer_5[569] ^ layer_5[592]); 
    assign layer_6[794] = ~(layer_5[961] ^ layer_5[968]); 
    wire [1:0] far_6_6915_0;    relay_conn far_6_6915_0_a(.in(layer_5[209]), .out(far_6_6915_0[0]));    relay_conn far_6_6915_0_b(.in(layer_5[102]), .out(far_6_6915_0[1]));
    wire [1:0] far_6_6915_1;    relay_conn far_6_6915_1_a(.in(far_6_6915_0[0]), .out(far_6_6915_1[0]));    relay_conn far_6_6915_1_b(.in(far_6_6915_0[1]), .out(far_6_6915_1[1]));
    wire [1:0] far_6_6915_2;    relay_conn far_6_6915_2_a(.in(far_6_6915_1[0]), .out(far_6_6915_2[0]));    relay_conn far_6_6915_2_b(.in(far_6_6915_1[1]), .out(far_6_6915_2[1]));
    assign layer_6[795] = ~(far_6_6915_2[0] ^ far_6_6915_2[1]); 
    assign layer_6[796] = ~layer_5[57]; 
    wire [1:0] far_6_6917_0;    relay_conn far_6_6917_0_a(.in(layer_5[330]), .out(far_6_6917_0[0]));    relay_conn far_6_6917_0_b(.in(layer_5[455]), .out(far_6_6917_0[1]));
    wire [1:0] far_6_6917_1;    relay_conn far_6_6917_1_a(.in(far_6_6917_0[0]), .out(far_6_6917_1[0]));    relay_conn far_6_6917_1_b(.in(far_6_6917_0[1]), .out(far_6_6917_1[1]));
    wire [1:0] far_6_6917_2;    relay_conn far_6_6917_2_a(.in(far_6_6917_1[0]), .out(far_6_6917_2[0]));    relay_conn far_6_6917_2_b(.in(far_6_6917_1[1]), .out(far_6_6917_2[1]));
    assign layer_6[797] = ~(far_6_6917_2[0] & far_6_6917_2[1]); 
    assign layer_6[798] = layer_5[968] & layer_5[971]; 
    assign layer_6[799] = ~(layer_5[414] & layer_5[398]); 
    wire [1:0] far_6_6920_0;    relay_conn far_6_6920_0_a(.in(layer_5[400]), .out(far_6_6920_0[0]));    relay_conn far_6_6920_0_b(.in(layer_5[513]), .out(far_6_6920_0[1]));
    wire [1:0] far_6_6920_1;    relay_conn far_6_6920_1_a(.in(far_6_6920_0[0]), .out(far_6_6920_1[0]));    relay_conn far_6_6920_1_b(.in(far_6_6920_0[1]), .out(far_6_6920_1[1]));
    wire [1:0] far_6_6920_2;    relay_conn far_6_6920_2_a(.in(far_6_6920_1[0]), .out(far_6_6920_2[0]));    relay_conn far_6_6920_2_b(.in(far_6_6920_1[1]), .out(far_6_6920_2[1]));
    assign layer_6[800] = ~(far_6_6920_2[0] | far_6_6920_2[1]); 
    wire [1:0] far_6_6921_0;    relay_conn far_6_6921_0_a(.in(layer_5[125]), .out(far_6_6921_0[0]));    relay_conn far_6_6921_0_b(.in(layer_5[196]), .out(far_6_6921_0[1]));
    wire [1:0] far_6_6921_1;    relay_conn far_6_6921_1_a(.in(far_6_6921_0[0]), .out(far_6_6921_1[0]));    relay_conn far_6_6921_1_b(.in(far_6_6921_0[1]), .out(far_6_6921_1[1]));
    assign layer_6[801] = far_6_6921_1[0] & ~far_6_6921_1[1]; 
    wire [1:0] far_6_6922_0;    relay_conn far_6_6922_0_a(.in(layer_5[673]), .out(far_6_6922_0[0]));    relay_conn far_6_6922_0_b(.in(layer_5[758]), .out(far_6_6922_0[1]));
    wire [1:0] far_6_6922_1;    relay_conn far_6_6922_1_a(.in(far_6_6922_0[0]), .out(far_6_6922_1[0]));    relay_conn far_6_6922_1_b(.in(far_6_6922_0[1]), .out(far_6_6922_1[1]));
    assign layer_6[802] = far_6_6922_1[0] & far_6_6922_1[1]; 
    wire [1:0] far_6_6923_0;    relay_conn far_6_6923_0_a(.in(layer_5[791]), .out(far_6_6923_0[0]));    relay_conn far_6_6923_0_b(.in(layer_5[746]), .out(far_6_6923_0[1]));
    assign layer_6[803] = far_6_6923_0[1] & ~far_6_6923_0[0]; 
    wire [1:0] far_6_6924_0;    relay_conn far_6_6924_0_a(.in(layer_5[773]), .out(far_6_6924_0[0]));    relay_conn far_6_6924_0_b(.in(layer_5[865]), .out(far_6_6924_0[1]));
    wire [1:0] far_6_6924_1;    relay_conn far_6_6924_1_a(.in(far_6_6924_0[0]), .out(far_6_6924_1[0]));    relay_conn far_6_6924_1_b(.in(far_6_6924_0[1]), .out(far_6_6924_1[1]));
    assign layer_6[804] = ~(far_6_6924_1[0] ^ far_6_6924_1[1]); 
    assign layer_6[805] = ~layer_5[89]; 
    wire [1:0] far_6_6926_0;    relay_conn far_6_6926_0_a(.in(layer_5[706]), .out(far_6_6926_0[0]));    relay_conn far_6_6926_0_b(.in(layer_5[596]), .out(far_6_6926_0[1]));
    wire [1:0] far_6_6926_1;    relay_conn far_6_6926_1_a(.in(far_6_6926_0[0]), .out(far_6_6926_1[0]));    relay_conn far_6_6926_1_b(.in(far_6_6926_0[1]), .out(far_6_6926_1[1]));
    wire [1:0] far_6_6926_2;    relay_conn far_6_6926_2_a(.in(far_6_6926_1[0]), .out(far_6_6926_2[0]));    relay_conn far_6_6926_2_b(.in(far_6_6926_1[1]), .out(far_6_6926_2[1]));
    assign layer_6[806] = far_6_6926_2[0] & ~far_6_6926_2[1]; 
    wire [1:0] far_6_6927_0;    relay_conn far_6_6927_0_a(.in(layer_5[962]), .out(far_6_6927_0[0]));    relay_conn far_6_6927_0_b(.in(layer_5[921]), .out(far_6_6927_0[1]));
    assign layer_6[807] = far_6_6927_0[0]; 
    wire [1:0] far_6_6928_0;    relay_conn far_6_6928_0_a(.in(layer_5[422]), .out(far_6_6928_0[0]));    relay_conn far_6_6928_0_b(.in(layer_5[480]), .out(far_6_6928_0[1]));
    assign layer_6[808] = far_6_6928_0[0]; 
    assign layer_6[809] = ~(layer_5[945] ^ layer_5[922]); 
    wire [1:0] far_6_6930_0;    relay_conn far_6_6930_0_a(.in(layer_5[209]), .out(far_6_6930_0[0]));    relay_conn far_6_6930_0_b(.in(layer_5[263]), .out(far_6_6930_0[1]));
    assign layer_6[810] = far_6_6930_0[1] & ~far_6_6930_0[0]; 
    wire [1:0] far_6_6931_0;    relay_conn far_6_6931_0_a(.in(layer_5[390]), .out(far_6_6931_0[0]));    relay_conn far_6_6931_0_b(.in(layer_5[296]), .out(far_6_6931_0[1]));
    wire [1:0] far_6_6931_1;    relay_conn far_6_6931_1_a(.in(far_6_6931_0[0]), .out(far_6_6931_1[0]));    relay_conn far_6_6931_1_b(.in(far_6_6931_0[1]), .out(far_6_6931_1[1]));
    assign layer_6[811] = far_6_6931_1[1]; 
    wire [1:0] far_6_6932_0;    relay_conn far_6_6932_0_a(.in(layer_5[533]), .out(far_6_6932_0[0]));    relay_conn far_6_6932_0_b(.in(layer_5[467]), .out(far_6_6932_0[1]));
    wire [1:0] far_6_6932_1;    relay_conn far_6_6932_1_a(.in(far_6_6932_0[0]), .out(far_6_6932_1[0]));    relay_conn far_6_6932_1_b(.in(far_6_6932_0[1]), .out(far_6_6932_1[1]));
    assign layer_6[812] = ~far_6_6932_1[0]; 
    wire [1:0] far_6_6933_0;    relay_conn far_6_6933_0_a(.in(layer_5[756]), .out(far_6_6933_0[0]));    relay_conn far_6_6933_0_b(.in(layer_5[791]), .out(far_6_6933_0[1]));
    assign layer_6[813] = far_6_6933_0[0] & far_6_6933_0[1]; 
    assign layer_6[814] = ~layer_5[962] | (layer_5[962] & layer_5[968]); 
    wire [1:0] far_6_6935_0;    relay_conn far_6_6935_0_a(.in(layer_5[706]), .out(far_6_6935_0[0]));    relay_conn far_6_6935_0_b(.in(layer_5[617]), .out(far_6_6935_0[1]));
    wire [1:0] far_6_6935_1;    relay_conn far_6_6935_1_a(.in(far_6_6935_0[0]), .out(far_6_6935_1[0]));    relay_conn far_6_6935_1_b(.in(far_6_6935_0[1]), .out(far_6_6935_1[1]));
    assign layer_6[815] = far_6_6935_1[0] & far_6_6935_1[1]; 
    wire [1:0] far_6_6936_0;    relay_conn far_6_6936_0_a(.in(layer_5[636]), .out(far_6_6936_0[0]));    relay_conn far_6_6936_0_b(.in(layer_5[737]), .out(far_6_6936_0[1]));
    wire [1:0] far_6_6936_1;    relay_conn far_6_6936_1_a(.in(far_6_6936_0[0]), .out(far_6_6936_1[0]));    relay_conn far_6_6936_1_b(.in(far_6_6936_0[1]), .out(far_6_6936_1[1]));
    wire [1:0] far_6_6936_2;    relay_conn far_6_6936_2_a(.in(far_6_6936_1[0]), .out(far_6_6936_2[0]));    relay_conn far_6_6936_2_b(.in(far_6_6936_1[1]), .out(far_6_6936_2[1]));
    assign layer_6[816] = ~(far_6_6936_2[0] ^ far_6_6936_2[1]); 
    assign layer_6[817] = ~layer_5[746]; 
    wire [1:0] far_6_6938_0;    relay_conn far_6_6938_0_a(.in(layer_5[559]), .out(far_6_6938_0[0]));    relay_conn far_6_6938_0_b(.in(layer_5[644]), .out(far_6_6938_0[1]));
    wire [1:0] far_6_6938_1;    relay_conn far_6_6938_1_a(.in(far_6_6938_0[0]), .out(far_6_6938_1[0]));    relay_conn far_6_6938_1_b(.in(far_6_6938_0[1]), .out(far_6_6938_1[1]));
    assign layer_6[818] = far_6_6938_1[0] & ~far_6_6938_1[1]; 
    assign layer_6[819] = ~layer_5[774]; 
    wire [1:0] far_6_6940_0;    relay_conn far_6_6940_0_a(.in(layer_5[748]), .out(far_6_6940_0[0]));    relay_conn far_6_6940_0_b(.in(layer_5[654]), .out(far_6_6940_0[1]));
    wire [1:0] far_6_6940_1;    relay_conn far_6_6940_1_a(.in(far_6_6940_0[0]), .out(far_6_6940_1[0]));    relay_conn far_6_6940_1_b(.in(far_6_6940_0[1]), .out(far_6_6940_1[1]));
    assign layer_6[820] = ~far_6_6940_1[1] | (far_6_6940_1[0] & far_6_6940_1[1]); 
    wire [1:0] far_6_6941_0;    relay_conn far_6_6941_0_a(.in(layer_5[527]), .out(far_6_6941_0[0]));    relay_conn far_6_6941_0_b(.in(layer_5[487]), .out(far_6_6941_0[1]));
    assign layer_6[821] = far_6_6941_0[0] ^ far_6_6941_0[1]; 
    wire [1:0] far_6_6942_0;    relay_conn far_6_6942_0_a(.in(layer_5[175]), .out(far_6_6942_0[0]));    relay_conn far_6_6942_0_b(.in(layer_5[128]), .out(far_6_6942_0[1]));
    assign layer_6[822] = ~(far_6_6942_0[0] | far_6_6942_0[1]); 
    wire [1:0] far_6_6943_0;    relay_conn far_6_6943_0_a(.in(layer_5[613]), .out(far_6_6943_0[0]));    relay_conn far_6_6943_0_b(.in(layer_5[550]), .out(far_6_6943_0[1]));
    assign layer_6[823] = ~(far_6_6943_0[0] & far_6_6943_0[1]); 
    wire [1:0] far_6_6944_0;    relay_conn far_6_6944_0_a(.in(layer_5[430]), .out(far_6_6944_0[0]));    relay_conn far_6_6944_0_b(.in(layer_5[493]), .out(far_6_6944_0[1]));
    assign layer_6[824] = ~far_6_6944_0[0]; 
    wire [1:0] far_6_6945_0;    relay_conn far_6_6945_0_a(.in(layer_5[48]), .out(far_6_6945_0[0]));    relay_conn far_6_6945_0_b(.in(layer_5[156]), .out(far_6_6945_0[1]));
    wire [1:0] far_6_6945_1;    relay_conn far_6_6945_1_a(.in(far_6_6945_0[0]), .out(far_6_6945_1[0]));    relay_conn far_6_6945_1_b(.in(far_6_6945_0[1]), .out(far_6_6945_1[1]));
    wire [1:0] far_6_6945_2;    relay_conn far_6_6945_2_a(.in(far_6_6945_1[0]), .out(far_6_6945_2[0]));    relay_conn far_6_6945_2_b(.in(far_6_6945_1[1]), .out(far_6_6945_2[1]));
    assign layer_6[825] = ~(far_6_6945_2[0] | far_6_6945_2[1]); 
    wire [1:0] far_6_6946_0;    relay_conn far_6_6946_0_a(.in(layer_5[553]), .out(far_6_6946_0[0]));    relay_conn far_6_6946_0_b(.in(layer_5[602]), .out(far_6_6946_0[1]));
    assign layer_6[826] = far_6_6946_0[0] | far_6_6946_0[1]; 
    wire [1:0] far_6_6947_0;    relay_conn far_6_6947_0_a(.in(layer_5[384]), .out(far_6_6947_0[0]));    relay_conn far_6_6947_0_b(.in(layer_5[432]), .out(far_6_6947_0[1]));
    assign layer_6[827] = far_6_6947_0[1]; 
    assign layer_6[828] = ~(layer_5[606] | layer_5[599]); 
    wire [1:0] far_6_6949_0;    relay_conn far_6_6949_0_a(.in(layer_5[888]), .out(far_6_6949_0[0]));    relay_conn far_6_6949_0_b(.in(layer_5[983]), .out(far_6_6949_0[1]));
    wire [1:0] far_6_6949_1;    relay_conn far_6_6949_1_a(.in(far_6_6949_0[0]), .out(far_6_6949_1[0]));    relay_conn far_6_6949_1_b(.in(far_6_6949_0[1]), .out(far_6_6949_1[1]));
    assign layer_6[829] = ~far_6_6949_1[0]; 
    wire [1:0] far_6_6950_0;    relay_conn far_6_6950_0_a(.in(layer_5[454]), .out(far_6_6950_0[0]));    relay_conn far_6_6950_0_b(.in(layer_5[557]), .out(far_6_6950_0[1]));
    wire [1:0] far_6_6950_1;    relay_conn far_6_6950_1_a(.in(far_6_6950_0[0]), .out(far_6_6950_1[0]));    relay_conn far_6_6950_1_b(.in(far_6_6950_0[1]), .out(far_6_6950_1[1]));
    wire [1:0] far_6_6950_2;    relay_conn far_6_6950_2_a(.in(far_6_6950_1[0]), .out(far_6_6950_2[0]));    relay_conn far_6_6950_2_b(.in(far_6_6950_1[1]), .out(far_6_6950_2[1]));
    assign layer_6[830] = ~(far_6_6950_2[0] | far_6_6950_2[1]); 
    wire [1:0] far_6_6951_0;    relay_conn far_6_6951_0_a(.in(layer_5[233]), .out(far_6_6951_0[0]));    relay_conn far_6_6951_0_b(.in(layer_5[122]), .out(far_6_6951_0[1]));
    wire [1:0] far_6_6951_1;    relay_conn far_6_6951_1_a(.in(far_6_6951_0[0]), .out(far_6_6951_1[0]));    relay_conn far_6_6951_1_b(.in(far_6_6951_0[1]), .out(far_6_6951_1[1]));
    wire [1:0] far_6_6951_2;    relay_conn far_6_6951_2_a(.in(far_6_6951_1[0]), .out(far_6_6951_2[0]));    relay_conn far_6_6951_2_b(.in(far_6_6951_1[1]), .out(far_6_6951_2[1]));
    assign layer_6[831] = far_6_6951_2[1]; 
    wire [1:0] far_6_6952_0;    relay_conn far_6_6952_0_a(.in(layer_5[60]), .out(far_6_6952_0[0]));    relay_conn far_6_6952_0_b(.in(layer_5[141]), .out(far_6_6952_0[1]));
    wire [1:0] far_6_6952_1;    relay_conn far_6_6952_1_a(.in(far_6_6952_0[0]), .out(far_6_6952_1[0]));    relay_conn far_6_6952_1_b(.in(far_6_6952_0[1]), .out(far_6_6952_1[1]));
    assign layer_6[832] = ~(far_6_6952_1[0] | far_6_6952_1[1]); 
    wire [1:0] far_6_6953_0;    relay_conn far_6_6953_0_a(.in(layer_5[218]), .out(far_6_6953_0[0]));    relay_conn far_6_6953_0_b(.in(layer_5[258]), .out(far_6_6953_0[1]));
    assign layer_6[833] = ~(far_6_6953_0[0] | far_6_6953_0[1]); 
    assign layer_6[834] = ~layer_5[450]; 
    assign layer_6[835] = layer_5[128] ^ layer_5[115]; 
    wire [1:0] far_6_6956_0;    relay_conn far_6_6956_0_a(.in(layer_5[304]), .out(far_6_6956_0[0]));    relay_conn far_6_6956_0_b(.in(layer_5[205]), .out(far_6_6956_0[1]));
    wire [1:0] far_6_6956_1;    relay_conn far_6_6956_1_a(.in(far_6_6956_0[0]), .out(far_6_6956_1[0]));    relay_conn far_6_6956_1_b(.in(far_6_6956_0[1]), .out(far_6_6956_1[1]));
    wire [1:0] far_6_6956_2;    relay_conn far_6_6956_2_a(.in(far_6_6956_1[0]), .out(far_6_6956_2[0]));    relay_conn far_6_6956_2_b(.in(far_6_6956_1[1]), .out(far_6_6956_2[1]));
    assign layer_6[836] = ~far_6_6956_2[1] | (far_6_6956_2[0] & far_6_6956_2[1]); 
    wire [1:0] far_6_6957_0;    relay_conn far_6_6957_0_a(.in(layer_5[850]), .out(far_6_6957_0[0]));    relay_conn far_6_6957_0_b(.in(layer_5[736]), .out(far_6_6957_0[1]));
    wire [1:0] far_6_6957_1;    relay_conn far_6_6957_1_a(.in(far_6_6957_0[0]), .out(far_6_6957_1[0]));    relay_conn far_6_6957_1_b(.in(far_6_6957_0[1]), .out(far_6_6957_1[1]));
    wire [1:0] far_6_6957_2;    relay_conn far_6_6957_2_a(.in(far_6_6957_1[0]), .out(far_6_6957_2[0]));    relay_conn far_6_6957_2_b(.in(far_6_6957_1[1]), .out(far_6_6957_2[1]));
    assign layer_6[837] = far_6_6957_2[1]; 
    assign layer_6[838] = ~(layer_5[944] & layer_5[938]); 
    assign layer_6[839] = layer_5[748] ^ layer_5[759]; 
    wire [1:0] far_6_6960_0;    relay_conn far_6_6960_0_a(.in(layer_5[927]), .out(far_6_6960_0[0]));    relay_conn far_6_6960_0_b(.in(layer_5[889]), .out(far_6_6960_0[1]));
    assign layer_6[840] = far_6_6960_0[0] & ~far_6_6960_0[1]; 
    assign layer_6[841] = layer_5[585] & ~layer_5[604]; 
    wire [1:0] far_6_6962_0;    relay_conn far_6_6962_0_a(.in(layer_5[688]), .out(far_6_6962_0[0]));    relay_conn far_6_6962_0_b(.in(layer_5[743]), .out(far_6_6962_0[1]));
    assign layer_6[842] = ~(far_6_6962_0[0] | far_6_6962_0[1]); 
    wire [1:0] far_6_6963_0;    relay_conn far_6_6963_0_a(.in(layer_5[159]), .out(far_6_6963_0[0]));    relay_conn far_6_6963_0_b(.in(layer_5[111]), .out(far_6_6963_0[1]));
    assign layer_6[843] = far_6_6963_0[0] | far_6_6963_0[1]; 
    wire [1:0] far_6_6964_0;    relay_conn far_6_6964_0_a(.in(layer_5[194]), .out(far_6_6964_0[0]));    relay_conn far_6_6964_0_b(.in(layer_5[229]), .out(far_6_6964_0[1]));
    assign layer_6[844] = ~far_6_6964_0[0]; 
    wire [1:0] far_6_6965_0;    relay_conn far_6_6965_0_a(.in(layer_5[0]), .out(far_6_6965_0[0]));    relay_conn far_6_6965_0_b(.in(layer_5[50]), .out(far_6_6965_0[1]));
    assign layer_6[845] = ~far_6_6965_0[1]; 
    wire [1:0] far_6_6966_0;    relay_conn far_6_6966_0_a(.in(layer_5[369]), .out(far_6_6966_0[0]));    relay_conn far_6_6966_0_b(.in(layer_5[439]), .out(far_6_6966_0[1]));
    wire [1:0] far_6_6966_1;    relay_conn far_6_6966_1_a(.in(far_6_6966_0[0]), .out(far_6_6966_1[0]));    relay_conn far_6_6966_1_b(.in(far_6_6966_0[1]), .out(far_6_6966_1[1]));
    assign layer_6[846] = ~far_6_6966_1[0] | (far_6_6966_1[0] & far_6_6966_1[1]); 
    wire [1:0] far_6_6967_0;    relay_conn far_6_6967_0_a(.in(layer_5[773]), .out(far_6_6967_0[0]));    relay_conn far_6_6967_0_b(.in(layer_5[886]), .out(far_6_6967_0[1]));
    wire [1:0] far_6_6967_1;    relay_conn far_6_6967_1_a(.in(far_6_6967_0[0]), .out(far_6_6967_1[0]));    relay_conn far_6_6967_1_b(.in(far_6_6967_0[1]), .out(far_6_6967_1[1]));
    wire [1:0] far_6_6967_2;    relay_conn far_6_6967_2_a(.in(far_6_6967_1[0]), .out(far_6_6967_2[0]));    relay_conn far_6_6967_2_b(.in(far_6_6967_1[1]), .out(far_6_6967_2[1]));
    assign layer_6[847] = far_6_6967_2[0] | far_6_6967_2[1]; 
    wire [1:0] far_6_6968_0;    relay_conn far_6_6968_0_a(.in(layer_5[369]), .out(far_6_6968_0[0]));    relay_conn far_6_6968_0_b(.in(layer_5[250]), .out(far_6_6968_0[1]));
    wire [1:0] far_6_6968_1;    relay_conn far_6_6968_1_a(.in(far_6_6968_0[0]), .out(far_6_6968_1[0]));    relay_conn far_6_6968_1_b(.in(far_6_6968_0[1]), .out(far_6_6968_1[1]));
    wire [1:0] far_6_6968_2;    relay_conn far_6_6968_2_a(.in(far_6_6968_1[0]), .out(far_6_6968_2[0]));    relay_conn far_6_6968_2_b(.in(far_6_6968_1[1]), .out(far_6_6968_2[1]));
    assign layer_6[848] = far_6_6968_2[0]; 
    wire [1:0] far_6_6969_0;    relay_conn far_6_6969_0_a(.in(layer_5[96]), .out(far_6_6969_0[0]));    relay_conn far_6_6969_0_b(.in(layer_5[16]), .out(far_6_6969_0[1]));
    wire [1:0] far_6_6969_1;    relay_conn far_6_6969_1_a(.in(far_6_6969_0[0]), .out(far_6_6969_1[0]));    relay_conn far_6_6969_1_b(.in(far_6_6969_0[1]), .out(far_6_6969_1[1]));
    assign layer_6[849] = far_6_6969_1[0] & far_6_6969_1[1]; 
    wire [1:0] far_6_6970_0;    relay_conn far_6_6970_0_a(.in(layer_5[436]), .out(far_6_6970_0[0]));    relay_conn far_6_6970_0_b(.in(layer_5[384]), .out(far_6_6970_0[1]));
    assign layer_6[850] = far_6_6970_0[0]; 
    wire [1:0] far_6_6971_0;    relay_conn far_6_6971_0_a(.in(layer_5[85]), .out(far_6_6971_0[0]));    relay_conn far_6_6971_0_b(.in(layer_5[203]), .out(far_6_6971_0[1]));
    wire [1:0] far_6_6971_1;    relay_conn far_6_6971_1_a(.in(far_6_6971_0[0]), .out(far_6_6971_1[0]));    relay_conn far_6_6971_1_b(.in(far_6_6971_0[1]), .out(far_6_6971_1[1]));
    wire [1:0] far_6_6971_2;    relay_conn far_6_6971_2_a(.in(far_6_6971_1[0]), .out(far_6_6971_2[0]));    relay_conn far_6_6971_2_b(.in(far_6_6971_1[1]), .out(far_6_6971_2[1]));
    assign layer_6[851] = far_6_6971_2[0]; 
    wire [1:0] far_6_6972_0;    relay_conn far_6_6972_0_a(.in(layer_5[254]), .out(far_6_6972_0[0]));    relay_conn far_6_6972_0_b(.in(layer_5[222]), .out(far_6_6972_0[1]));
    assign layer_6[852] = ~far_6_6972_0[0]; 
    wire [1:0] far_6_6973_0;    relay_conn far_6_6973_0_a(.in(layer_5[286]), .out(far_6_6973_0[0]));    relay_conn far_6_6973_0_b(.in(layer_5[221]), .out(far_6_6973_0[1]));
    wire [1:0] far_6_6973_1;    relay_conn far_6_6973_1_a(.in(far_6_6973_0[0]), .out(far_6_6973_1[0]));    relay_conn far_6_6973_1_b(.in(far_6_6973_0[1]), .out(far_6_6973_1[1]));
    assign layer_6[853] = far_6_6973_1[1]; 
    assign layer_6[854] = layer_5[436] & ~layer_5[438]; 
    wire [1:0] far_6_6975_0;    relay_conn far_6_6975_0_a(.in(layer_5[769]), .out(far_6_6975_0[0]));    relay_conn far_6_6975_0_b(.in(layer_5[860]), .out(far_6_6975_0[1]));
    wire [1:0] far_6_6975_1;    relay_conn far_6_6975_1_a(.in(far_6_6975_0[0]), .out(far_6_6975_1[0]));    relay_conn far_6_6975_1_b(.in(far_6_6975_0[1]), .out(far_6_6975_1[1]));
    assign layer_6[855] = far_6_6975_1[0]; 
    wire [1:0] far_6_6976_0;    relay_conn far_6_6976_0_a(.in(layer_5[654]), .out(far_6_6976_0[0]));    relay_conn far_6_6976_0_b(.in(layer_5[777]), .out(far_6_6976_0[1]));
    wire [1:0] far_6_6976_1;    relay_conn far_6_6976_1_a(.in(far_6_6976_0[0]), .out(far_6_6976_1[0]));    relay_conn far_6_6976_1_b(.in(far_6_6976_0[1]), .out(far_6_6976_1[1]));
    wire [1:0] far_6_6976_2;    relay_conn far_6_6976_2_a(.in(far_6_6976_1[0]), .out(far_6_6976_2[0]));    relay_conn far_6_6976_2_b(.in(far_6_6976_1[1]), .out(far_6_6976_2[1]));
    assign layer_6[856] = ~(far_6_6976_2[0] | far_6_6976_2[1]); 
    assign layer_6[857] = layer_5[452] & ~layer_5[477]; 
    wire [1:0] far_6_6978_0;    relay_conn far_6_6978_0_a(.in(layer_5[691]), .out(far_6_6978_0[0]));    relay_conn far_6_6978_0_b(.in(layer_5[596]), .out(far_6_6978_0[1]));
    wire [1:0] far_6_6978_1;    relay_conn far_6_6978_1_a(.in(far_6_6978_0[0]), .out(far_6_6978_1[0]));    relay_conn far_6_6978_1_b(.in(far_6_6978_0[1]), .out(far_6_6978_1[1]));
    assign layer_6[858] = ~far_6_6978_1[1]; 
    wire [1:0] far_6_6979_0;    relay_conn far_6_6979_0_a(.in(layer_5[225]), .out(far_6_6979_0[0]));    relay_conn far_6_6979_0_b(.in(layer_5[115]), .out(far_6_6979_0[1]));
    wire [1:0] far_6_6979_1;    relay_conn far_6_6979_1_a(.in(far_6_6979_0[0]), .out(far_6_6979_1[0]));    relay_conn far_6_6979_1_b(.in(far_6_6979_0[1]), .out(far_6_6979_1[1]));
    wire [1:0] far_6_6979_2;    relay_conn far_6_6979_2_a(.in(far_6_6979_1[0]), .out(far_6_6979_2[0]));    relay_conn far_6_6979_2_b(.in(far_6_6979_1[1]), .out(far_6_6979_2[1]));
    assign layer_6[859] = ~far_6_6979_2[0]; 
    assign layer_6[860] = layer_5[430] & ~layer_5[400]; 
    wire [1:0] far_6_6981_0;    relay_conn far_6_6981_0_a(.in(layer_5[921]), .out(far_6_6981_0[0]));    relay_conn far_6_6981_0_b(.in(layer_5[1015]), .out(far_6_6981_0[1]));
    wire [1:0] far_6_6981_1;    relay_conn far_6_6981_1_a(.in(far_6_6981_0[0]), .out(far_6_6981_1[0]));    relay_conn far_6_6981_1_b(.in(far_6_6981_0[1]), .out(far_6_6981_1[1]));
    assign layer_6[861] = far_6_6981_1[1]; 
    wire [1:0] far_6_6982_0;    relay_conn far_6_6982_0_a(.in(layer_5[424]), .out(far_6_6982_0[0]));    relay_conn far_6_6982_0_b(.in(layer_5[356]), .out(far_6_6982_0[1]));
    wire [1:0] far_6_6982_1;    relay_conn far_6_6982_1_a(.in(far_6_6982_0[0]), .out(far_6_6982_1[0]));    relay_conn far_6_6982_1_b(.in(far_6_6982_0[1]), .out(far_6_6982_1[1]));
    assign layer_6[862] = far_6_6982_1[0] & ~far_6_6982_1[1]; 
    wire [1:0] far_6_6983_0;    relay_conn far_6_6983_0_a(.in(layer_5[19]), .out(far_6_6983_0[0]));    relay_conn far_6_6983_0_b(.in(layer_5[115]), .out(far_6_6983_0[1]));
    wire [1:0] far_6_6983_1;    relay_conn far_6_6983_1_a(.in(far_6_6983_0[0]), .out(far_6_6983_1[0]));    relay_conn far_6_6983_1_b(.in(far_6_6983_0[1]), .out(far_6_6983_1[1]));
    wire [1:0] far_6_6983_2;    relay_conn far_6_6983_2_a(.in(far_6_6983_1[0]), .out(far_6_6983_2[0]));    relay_conn far_6_6983_2_b(.in(far_6_6983_1[1]), .out(far_6_6983_2[1]));
    assign layer_6[863] = ~(far_6_6983_2[0] ^ far_6_6983_2[1]); 
    assign layer_6[864] = ~(layer_5[761] | layer_5[734]); 
    assign layer_6[865] = ~layer_5[915]; 
    wire [1:0] far_6_6986_0;    relay_conn far_6_6986_0_a(.in(layer_5[512]), .out(far_6_6986_0[0]));    relay_conn far_6_6986_0_b(.in(layer_5[473]), .out(far_6_6986_0[1]));
    assign layer_6[866] = ~far_6_6986_0[0]; 
    wire [1:0] far_6_6987_0;    relay_conn far_6_6987_0_a(.in(layer_5[339]), .out(far_6_6987_0[0]));    relay_conn far_6_6987_0_b(.in(layer_5[304]), .out(far_6_6987_0[1]));
    assign layer_6[867] = far_6_6987_0[0] & ~far_6_6987_0[1]; 
    wire [1:0] far_6_6988_0;    relay_conn far_6_6988_0_a(.in(layer_5[924]), .out(far_6_6988_0[0]));    relay_conn far_6_6988_0_b(.in(layer_5[886]), .out(far_6_6988_0[1]));
    assign layer_6[868] = far_6_6988_0[0] ^ far_6_6988_0[1]; 
    assign layer_6[869] = ~layer_5[396]; 
    wire [1:0] far_6_6990_0;    relay_conn far_6_6990_0_a(.in(layer_5[581]), .out(far_6_6990_0[0]));    relay_conn far_6_6990_0_b(.in(layer_5[656]), .out(far_6_6990_0[1]));
    wire [1:0] far_6_6990_1;    relay_conn far_6_6990_1_a(.in(far_6_6990_0[0]), .out(far_6_6990_1[0]));    relay_conn far_6_6990_1_b(.in(far_6_6990_0[1]), .out(far_6_6990_1[1]));
    assign layer_6[870] = ~far_6_6990_1[0] | (far_6_6990_1[0] & far_6_6990_1[1]); 
    wire [1:0] far_6_6991_0;    relay_conn far_6_6991_0_a(.in(layer_5[837]), .out(far_6_6991_0[0]));    relay_conn far_6_6991_0_b(.in(layer_5[751]), .out(far_6_6991_0[1]));
    wire [1:0] far_6_6991_1;    relay_conn far_6_6991_1_a(.in(far_6_6991_0[0]), .out(far_6_6991_1[0]));    relay_conn far_6_6991_1_b(.in(far_6_6991_0[1]), .out(far_6_6991_1[1]));
    assign layer_6[871] = far_6_6991_1[0] ^ far_6_6991_1[1]; 
    wire [1:0] far_6_6992_0;    relay_conn far_6_6992_0_a(.in(layer_5[271]), .out(far_6_6992_0[0]));    relay_conn far_6_6992_0_b(.in(layer_5[211]), .out(far_6_6992_0[1]));
    assign layer_6[872] = far_6_6992_0[0] ^ far_6_6992_0[1]; 
    assign layer_6[873] = layer_5[234] & layer_5[218]; 
    wire [1:0] far_6_6994_0;    relay_conn far_6_6994_0_a(.in(layer_5[467]), .out(far_6_6994_0[0]));    relay_conn far_6_6994_0_b(.in(layer_5[561]), .out(far_6_6994_0[1]));
    wire [1:0] far_6_6994_1;    relay_conn far_6_6994_1_a(.in(far_6_6994_0[0]), .out(far_6_6994_1[0]));    relay_conn far_6_6994_1_b(.in(far_6_6994_0[1]), .out(far_6_6994_1[1]));
    assign layer_6[874] = ~far_6_6994_1[1] | (far_6_6994_1[0] & far_6_6994_1[1]); 
    wire [1:0] far_6_6995_0;    relay_conn far_6_6995_0_a(.in(layer_5[832]), .out(far_6_6995_0[0]));    relay_conn far_6_6995_0_b(.in(layer_5[751]), .out(far_6_6995_0[1]));
    wire [1:0] far_6_6995_1;    relay_conn far_6_6995_1_a(.in(far_6_6995_0[0]), .out(far_6_6995_1[0]));    relay_conn far_6_6995_1_b(.in(far_6_6995_0[1]), .out(far_6_6995_1[1]));
    assign layer_6[875] = far_6_6995_1[0] & far_6_6995_1[1]; 
    assign layer_6[876] = ~(layer_5[956] & layer_5[980]); 
    wire [1:0] far_6_6997_0;    relay_conn far_6_6997_0_a(.in(layer_5[149]), .out(far_6_6997_0[0]));    relay_conn far_6_6997_0_b(.in(layer_5[32]), .out(far_6_6997_0[1]));
    wire [1:0] far_6_6997_1;    relay_conn far_6_6997_1_a(.in(far_6_6997_0[0]), .out(far_6_6997_1[0]));    relay_conn far_6_6997_1_b(.in(far_6_6997_0[1]), .out(far_6_6997_1[1]));
    wire [1:0] far_6_6997_2;    relay_conn far_6_6997_2_a(.in(far_6_6997_1[0]), .out(far_6_6997_2[0]));    relay_conn far_6_6997_2_b(.in(far_6_6997_1[1]), .out(far_6_6997_2[1]));
    assign layer_6[877] = ~far_6_6997_2[1] | (far_6_6997_2[0] & far_6_6997_2[1]); 
    wire [1:0] far_6_6998_0;    relay_conn far_6_6998_0_a(.in(layer_5[657]), .out(far_6_6998_0[0]));    relay_conn far_6_6998_0_b(.in(layer_5[773]), .out(far_6_6998_0[1]));
    wire [1:0] far_6_6998_1;    relay_conn far_6_6998_1_a(.in(far_6_6998_0[0]), .out(far_6_6998_1[0]));    relay_conn far_6_6998_1_b(.in(far_6_6998_0[1]), .out(far_6_6998_1[1]));
    wire [1:0] far_6_6998_2;    relay_conn far_6_6998_2_a(.in(far_6_6998_1[0]), .out(far_6_6998_2[0]));    relay_conn far_6_6998_2_b(.in(far_6_6998_1[1]), .out(far_6_6998_2[1]));
    assign layer_6[878] = far_6_6998_2[1]; 
    assign layer_6[879] = ~(layer_5[864] | layer_5[869]); 
    assign layer_6[880] = ~(layer_5[127] & layer_5[121]); 
    wire [1:0] far_6_7001_0;    relay_conn far_6_7001_0_a(.in(layer_5[430]), .out(far_6_7001_0[0]));    relay_conn far_6_7001_0_b(.in(layer_5[357]), .out(far_6_7001_0[1]));
    wire [1:0] far_6_7001_1;    relay_conn far_6_7001_1_a(.in(far_6_7001_0[0]), .out(far_6_7001_1[0]));    relay_conn far_6_7001_1_b(.in(far_6_7001_0[1]), .out(far_6_7001_1[1]));
    assign layer_6[881] = ~far_6_7001_1[0]; 
    wire [1:0] far_6_7002_0;    relay_conn far_6_7002_0_a(.in(layer_5[430]), .out(far_6_7002_0[0]));    relay_conn far_6_7002_0_b(.in(layer_5[315]), .out(far_6_7002_0[1]));
    wire [1:0] far_6_7002_1;    relay_conn far_6_7002_1_a(.in(far_6_7002_0[0]), .out(far_6_7002_1[0]));    relay_conn far_6_7002_1_b(.in(far_6_7002_0[1]), .out(far_6_7002_1[1]));
    wire [1:0] far_6_7002_2;    relay_conn far_6_7002_2_a(.in(far_6_7002_1[0]), .out(far_6_7002_2[0]));    relay_conn far_6_7002_2_b(.in(far_6_7002_1[1]), .out(far_6_7002_2[1]));
    assign layer_6[882] = far_6_7002_2[0]; 
    wire [1:0] far_6_7003_0;    relay_conn far_6_7003_0_a(.in(layer_5[57]), .out(far_6_7003_0[0]));    relay_conn far_6_7003_0_b(.in(layer_5[128]), .out(far_6_7003_0[1]));
    wire [1:0] far_6_7003_1;    relay_conn far_6_7003_1_a(.in(far_6_7003_0[0]), .out(far_6_7003_1[0]));    relay_conn far_6_7003_1_b(.in(far_6_7003_0[1]), .out(far_6_7003_1[1]));
    assign layer_6[883] = ~far_6_7003_1[0] | (far_6_7003_1[0] & far_6_7003_1[1]); 
    wire [1:0] far_6_7004_0;    relay_conn far_6_7004_0_a(.in(layer_5[390]), .out(far_6_7004_0[0]));    relay_conn far_6_7004_0_b(.in(layer_5[487]), .out(far_6_7004_0[1]));
    wire [1:0] far_6_7004_1;    relay_conn far_6_7004_1_a(.in(far_6_7004_0[0]), .out(far_6_7004_1[0]));    relay_conn far_6_7004_1_b(.in(far_6_7004_0[1]), .out(far_6_7004_1[1]));
    wire [1:0] far_6_7004_2;    relay_conn far_6_7004_2_a(.in(far_6_7004_1[0]), .out(far_6_7004_2[0]));    relay_conn far_6_7004_2_b(.in(far_6_7004_1[1]), .out(far_6_7004_2[1]));
    assign layer_6[884] = ~far_6_7004_2[0] | (far_6_7004_2[0] & far_6_7004_2[1]); 
    assign layer_6[885] = ~layer_5[151]; 
    assign layer_6[886] = ~layer_5[111] | (layer_5[83] & layer_5[111]); 
    assign layer_6[887] = layer_5[152]; 
    wire [1:0] far_6_7008_0;    relay_conn far_6_7008_0_a(.in(layer_5[434]), .out(far_6_7008_0[0]));    relay_conn far_6_7008_0_b(.in(layer_5[346]), .out(far_6_7008_0[1]));
    wire [1:0] far_6_7008_1;    relay_conn far_6_7008_1_a(.in(far_6_7008_0[0]), .out(far_6_7008_1[0]));    relay_conn far_6_7008_1_b(.in(far_6_7008_0[1]), .out(far_6_7008_1[1]));
    assign layer_6[888] = far_6_7008_1[0] & far_6_7008_1[1]; 
    wire [1:0] far_6_7009_0;    relay_conn far_6_7009_0_a(.in(layer_5[894]), .out(far_6_7009_0[0]));    relay_conn far_6_7009_0_b(.in(layer_5[977]), .out(far_6_7009_0[1]));
    wire [1:0] far_6_7009_1;    relay_conn far_6_7009_1_a(.in(far_6_7009_0[0]), .out(far_6_7009_1[0]));    relay_conn far_6_7009_1_b(.in(far_6_7009_0[1]), .out(far_6_7009_1[1]));
    assign layer_6[889] = far_6_7009_1[1]; 
    wire [1:0] far_6_7010_0;    relay_conn far_6_7010_0_a(.in(layer_5[690]), .out(far_6_7010_0[0]));    relay_conn far_6_7010_0_b(.in(layer_5[741]), .out(far_6_7010_0[1]));
    assign layer_6[890] = ~(far_6_7010_0[0] | far_6_7010_0[1]); 
    assign layer_6[891] = ~(layer_5[185] & layer_5[156]); 
    wire [1:0] far_6_7012_0;    relay_conn far_6_7012_0_a(.in(layer_5[1001]), .out(far_6_7012_0[0]));    relay_conn far_6_7012_0_b(.in(layer_5[915]), .out(far_6_7012_0[1]));
    wire [1:0] far_6_7012_1;    relay_conn far_6_7012_1_a(.in(far_6_7012_0[0]), .out(far_6_7012_1[0]));    relay_conn far_6_7012_1_b(.in(far_6_7012_0[1]), .out(far_6_7012_1[1]));
    assign layer_6[892] = far_6_7012_1[1]; 
    assign layer_6[893] = ~(layer_5[839] ^ layer_5[849]); 
    wire [1:0] far_6_7014_0;    relay_conn far_6_7014_0_a(.in(layer_5[832]), .out(far_6_7014_0[0]));    relay_conn far_6_7014_0_b(.in(layer_5[766]), .out(far_6_7014_0[1]));
    wire [1:0] far_6_7014_1;    relay_conn far_6_7014_1_a(.in(far_6_7014_0[0]), .out(far_6_7014_1[0]));    relay_conn far_6_7014_1_b(.in(far_6_7014_0[1]), .out(far_6_7014_1[1]));
    assign layer_6[894] = ~(far_6_7014_1[0] & far_6_7014_1[1]); 
    wire [1:0] far_6_7015_0;    relay_conn far_6_7015_0_a(.in(layer_5[732]), .out(far_6_7015_0[0]));    relay_conn far_6_7015_0_b(.in(layer_5[773]), .out(far_6_7015_0[1]));
    assign layer_6[895] = far_6_7015_0[0] & far_6_7015_0[1]; 
    wire [1:0] far_6_7016_0;    relay_conn far_6_7016_0_a(.in(layer_5[820]), .out(far_6_7016_0[0]));    relay_conn far_6_7016_0_b(.in(layer_5[694]), .out(far_6_7016_0[1]));
    wire [1:0] far_6_7016_1;    relay_conn far_6_7016_1_a(.in(far_6_7016_0[0]), .out(far_6_7016_1[0]));    relay_conn far_6_7016_1_b(.in(far_6_7016_0[1]), .out(far_6_7016_1[1]));
    wire [1:0] far_6_7016_2;    relay_conn far_6_7016_2_a(.in(far_6_7016_1[0]), .out(far_6_7016_2[0]));    relay_conn far_6_7016_2_b(.in(far_6_7016_1[1]), .out(far_6_7016_2[1]));
    assign layer_6[896] = far_6_7016_2[0] & far_6_7016_2[1]; 
    assign layer_6[897] = layer_5[788] & layer_5[786]; 
    assign layer_6[898] = ~layer_5[19] | (layer_5[19] & layer_5[6]); 
    wire [1:0] far_6_7019_0;    relay_conn far_6_7019_0_a(.in(layer_5[581]), .out(far_6_7019_0[0]));    relay_conn far_6_7019_0_b(.in(layer_5[518]), .out(far_6_7019_0[1]));
    assign layer_6[899] = far_6_7019_0[1] & ~far_6_7019_0[0]; 
    assign layer_6[900] = ~(layer_5[871] ^ layer_5[873]); 
    wire [1:0] far_6_7021_0;    relay_conn far_6_7021_0_a(.in(layer_5[791]), .out(far_6_7021_0[0]));    relay_conn far_6_7021_0_b(.in(layer_5[891]), .out(far_6_7021_0[1]));
    wire [1:0] far_6_7021_1;    relay_conn far_6_7021_1_a(.in(far_6_7021_0[0]), .out(far_6_7021_1[0]));    relay_conn far_6_7021_1_b(.in(far_6_7021_0[1]), .out(far_6_7021_1[1]));
    wire [1:0] far_6_7021_2;    relay_conn far_6_7021_2_a(.in(far_6_7021_1[0]), .out(far_6_7021_2[0]));    relay_conn far_6_7021_2_b(.in(far_6_7021_1[1]), .out(far_6_7021_2[1]));
    assign layer_6[901] = ~far_6_7021_2[0] | (far_6_7021_2[0] & far_6_7021_2[1]); 
    wire [1:0] far_6_7022_0;    relay_conn far_6_7022_0_a(.in(layer_5[529]), .out(far_6_7022_0[0]));    relay_conn far_6_7022_0_b(.in(layer_5[636]), .out(far_6_7022_0[1]));
    wire [1:0] far_6_7022_1;    relay_conn far_6_7022_1_a(.in(far_6_7022_0[0]), .out(far_6_7022_1[0]));    relay_conn far_6_7022_1_b(.in(far_6_7022_0[1]), .out(far_6_7022_1[1]));
    wire [1:0] far_6_7022_2;    relay_conn far_6_7022_2_a(.in(far_6_7022_1[0]), .out(far_6_7022_2[0]));    relay_conn far_6_7022_2_b(.in(far_6_7022_1[1]), .out(far_6_7022_2[1]));
    assign layer_6[902] = far_6_7022_2[0] | far_6_7022_2[1]; 
    assign layer_6[903] = ~layer_5[950]; 
    wire [1:0] far_6_7024_0;    relay_conn far_6_7024_0_a(.in(layer_5[815]), .out(far_6_7024_0[0]));    relay_conn far_6_7024_0_b(.in(layer_5[932]), .out(far_6_7024_0[1]));
    wire [1:0] far_6_7024_1;    relay_conn far_6_7024_1_a(.in(far_6_7024_0[0]), .out(far_6_7024_1[0]));    relay_conn far_6_7024_1_b(.in(far_6_7024_0[1]), .out(far_6_7024_1[1]));
    wire [1:0] far_6_7024_2;    relay_conn far_6_7024_2_a(.in(far_6_7024_1[0]), .out(far_6_7024_2[0]));    relay_conn far_6_7024_2_b(.in(far_6_7024_1[1]), .out(far_6_7024_2[1]));
    assign layer_6[904] = far_6_7024_2[0] & far_6_7024_2[1]; 
    wire [1:0] far_6_7025_0;    relay_conn far_6_7025_0_a(.in(layer_5[840]), .out(far_6_7025_0[0]));    relay_conn far_6_7025_0_b(.in(layer_5[930]), .out(far_6_7025_0[1]));
    wire [1:0] far_6_7025_1;    relay_conn far_6_7025_1_a(.in(far_6_7025_0[0]), .out(far_6_7025_1[0]));    relay_conn far_6_7025_1_b(.in(far_6_7025_0[1]), .out(far_6_7025_1[1]));
    assign layer_6[905] = ~far_6_7025_1[0] | (far_6_7025_1[0] & far_6_7025_1[1]); 
    wire [1:0] far_6_7026_0;    relay_conn far_6_7026_0_a(.in(layer_5[111]), .out(far_6_7026_0[0]));    relay_conn far_6_7026_0_b(.in(layer_5[229]), .out(far_6_7026_0[1]));
    wire [1:0] far_6_7026_1;    relay_conn far_6_7026_1_a(.in(far_6_7026_0[0]), .out(far_6_7026_1[0]));    relay_conn far_6_7026_1_b(.in(far_6_7026_0[1]), .out(far_6_7026_1[1]));
    wire [1:0] far_6_7026_2;    relay_conn far_6_7026_2_a(.in(far_6_7026_1[0]), .out(far_6_7026_2[0]));    relay_conn far_6_7026_2_b(.in(far_6_7026_1[1]), .out(far_6_7026_2[1]));
    assign layer_6[906] = ~(far_6_7026_2[0] ^ far_6_7026_2[1]); 
    wire [1:0] far_6_7027_0;    relay_conn far_6_7027_0_a(.in(layer_5[505]), .out(far_6_7027_0[0]));    relay_conn far_6_7027_0_b(.in(layer_5[443]), .out(far_6_7027_0[1]));
    assign layer_6[907] = far_6_7027_0[0] & ~far_6_7027_0[1]; 
    assign layer_6[908] = layer_5[199]; 
    wire [1:0] far_6_7029_0;    relay_conn far_6_7029_0_a(.in(layer_5[328]), .out(far_6_7029_0[0]));    relay_conn far_6_7029_0_b(.in(layer_5[261]), .out(far_6_7029_0[1]));
    wire [1:0] far_6_7029_1;    relay_conn far_6_7029_1_a(.in(far_6_7029_0[0]), .out(far_6_7029_1[0]));    relay_conn far_6_7029_1_b(.in(far_6_7029_0[1]), .out(far_6_7029_1[1]));
    assign layer_6[909] = far_6_7029_1[1]; 
    wire [1:0] far_6_7030_0;    relay_conn far_6_7030_0_a(.in(layer_5[214]), .out(far_6_7030_0[0]));    relay_conn far_6_7030_0_b(.in(layer_5[94]), .out(far_6_7030_0[1]));
    wire [1:0] far_6_7030_1;    relay_conn far_6_7030_1_a(.in(far_6_7030_0[0]), .out(far_6_7030_1[0]));    relay_conn far_6_7030_1_b(.in(far_6_7030_0[1]), .out(far_6_7030_1[1]));
    wire [1:0] far_6_7030_2;    relay_conn far_6_7030_2_a(.in(far_6_7030_1[0]), .out(far_6_7030_2[0]));    relay_conn far_6_7030_2_b(.in(far_6_7030_1[1]), .out(far_6_7030_2[1]));
    assign layer_6[910] = far_6_7030_2[1]; 
    wire [1:0] far_6_7031_0;    relay_conn far_6_7031_0_a(.in(layer_5[469]), .out(far_6_7031_0[0]));    relay_conn far_6_7031_0_b(.in(layer_5[389]), .out(far_6_7031_0[1]));
    wire [1:0] far_6_7031_1;    relay_conn far_6_7031_1_a(.in(far_6_7031_0[0]), .out(far_6_7031_1[0]));    relay_conn far_6_7031_1_b(.in(far_6_7031_0[1]), .out(far_6_7031_1[1]));
    assign layer_6[911] = far_6_7031_1[1]; 
    wire [1:0] far_6_7032_0;    relay_conn far_6_7032_0_a(.in(layer_5[653]), .out(far_6_7032_0[0]));    relay_conn far_6_7032_0_b(.in(layer_5[737]), .out(far_6_7032_0[1]));
    wire [1:0] far_6_7032_1;    relay_conn far_6_7032_1_a(.in(far_6_7032_0[0]), .out(far_6_7032_1[0]));    relay_conn far_6_7032_1_b(.in(far_6_7032_0[1]), .out(far_6_7032_1[1]));
    assign layer_6[912] = far_6_7032_1[1] & ~far_6_7032_1[0]; 
    assign layer_6[913] = layer_5[682] & ~layer_5[688]; 
    assign layer_6[914] = layer_5[980] & layer_5[976]; 
    wire [1:0] far_6_7035_0;    relay_conn far_6_7035_0_a(.in(layer_5[721]), .out(far_6_7035_0[0]));    relay_conn far_6_7035_0_b(.in(layer_5[668]), .out(far_6_7035_0[1]));
    assign layer_6[915] = far_6_7035_0[0] & ~far_6_7035_0[1]; 
    wire [1:0] far_6_7036_0;    relay_conn far_6_7036_0_a(.in(layer_5[939]), .out(far_6_7036_0[0]));    relay_conn far_6_7036_0_b(.in(layer_5[847]), .out(far_6_7036_0[1]));
    wire [1:0] far_6_7036_1;    relay_conn far_6_7036_1_a(.in(far_6_7036_0[0]), .out(far_6_7036_1[0]));    relay_conn far_6_7036_1_b(.in(far_6_7036_0[1]), .out(far_6_7036_1[1]));
    assign layer_6[916] = ~far_6_7036_1[1]; 
    wire [1:0] far_6_7037_0;    relay_conn far_6_7037_0_a(.in(layer_5[452]), .out(far_6_7037_0[0]));    relay_conn far_6_7037_0_b(.in(layer_5[402]), .out(far_6_7037_0[1]));
    assign layer_6[917] = far_6_7037_0[0] ^ far_6_7037_0[1]; 
    wire [1:0] far_6_7038_0;    relay_conn far_6_7038_0_a(.in(layer_5[643]), .out(far_6_7038_0[0]));    relay_conn far_6_7038_0_b(.in(layer_5[595]), .out(far_6_7038_0[1]));
    assign layer_6[918] = ~far_6_7038_0[1] | (far_6_7038_0[0] & far_6_7038_0[1]); 
    wire [1:0] far_6_7039_0;    relay_conn far_6_7039_0_a(.in(layer_5[870]), .out(far_6_7039_0[0]));    relay_conn far_6_7039_0_b(.in(layer_5[832]), .out(far_6_7039_0[1]));
    assign layer_6[919] = ~far_6_7039_0[1] | (far_6_7039_0[0] & far_6_7039_0[1]); 
    assign layer_6[920] = ~(layer_5[968] ^ layer_5[949]); 
    wire [1:0] far_6_7041_0;    relay_conn far_6_7041_0_a(.in(layer_5[576]), .out(far_6_7041_0[0]));    relay_conn far_6_7041_0_b(.in(layer_5[474]), .out(far_6_7041_0[1]));
    wire [1:0] far_6_7041_1;    relay_conn far_6_7041_1_a(.in(far_6_7041_0[0]), .out(far_6_7041_1[0]));    relay_conn far_6_7041_1_b(.in(far_6_7041_0[1]), .out(far_6_7041_1[1]));
    wire [1:0] far_6_7041_2;    relay_conn far_6_7041_2_a(.in(far_6_7041_1[0]), .out(far_6_7041_2[0]));    relay_conn far_6_7041_2_b(.in(far_6_7041_1[1]), .out(far_6_7041_2[1]));
    assign layer_6[921] = ~(far_6_7041_2[0] ^ far_6_7041_2[1]); 
    wire [1:0] far_6_7042_0;    relay_conn far_6_7042_0_a(.in(layer_5[875]), .out(far_6_7042_0[0]));    relay_conn far_6_7042_0_b(.in(layer_5[777]), .out(far_6_7042_0[1]));
    wire [1:0] far_6_7042_1;    relay_conn far_6_7042_1_a(.in(far_6_7042_0[0]), .out(far_6_7042_1[0]));    relay_conn far_6_7042_1_b(.in(far_6_7042_0[1]), .out(far_6_7042_1[1]));
    wire [1:0] far_6_7042_2;    relay_conn far_6_7042_2_a(.in(far_6_7042_1[0]), .out(far_6_7042_2[0]));    relay_conn far_6_7042_2_b(.in(far_6_7042_1[1]), .out(far_6_7042_2[1]));
    assign layer_6[922] = ~(far_6_7042_2[0] ^ far_6_7042_2[1]); 
    wire [1:0] far_6_7043_0;    relay_conn far_6_7043_0_a(.in(layer_5[746]), .out(far_6_7043_0[0]));    relay_conn far_6_7043_0_b(.in(layer_5[706]), .out(far_6_7043_0[1]));
    assign layer_6[923] = ~far_6_7043_0[0] | (far_6_7043_0[0] & far_6_7043_0[1]); 
    assign layer_6[924] = ~(layer_5[756] & layer_5[763]); 
    assign layer_6[925] = layer_5[891] & ~layer_5[893]; 
    assign layer_6[926] = ~layer_5[369] | (layer_5[396] & layer_5[369]); 
    wire [1:0] far_6_7047_0;    relay_conn far_6_7047_0_a(.in(layer_5[976]), .out(far_6_7047_0[0]));    relay_conn far_6_7047_0_b(.in(layer_5[906]), .out(far_6_7047_0[1]));
    wire [1:0] far_6_7047_1;    relay_conn far_6_7047_1_a(.in(far_6_7047_0[0]), .out(far_6_7047_1[0]));    relay_conn far_6_7047_1_b(.in(far_6_7047_0[1]), .out(far_6_7047_1[1]));
    assign layer_6[927] = ~far_6_7047_1[0]; 
    wire [1:0] far_6_7048_0;    relay_conn far_6_7048_0_a(.in(layer_5[79]), .out(far_6_7048_0[0]));    relay_conn far_6_7048_0_b(.in(layer_5[169]), .out(far_6_7048_0[1]));
    wire [1:0] far_6_7048_1;    relay_conn far_6_7048_1_a(.in(far_6_7048_0[0]), .out(far_6_7048_1[0]));    relay_conn far_6_7048_1_b(.in(far_6_7048_0[1]), .out(far_6_7048_1[1]));
    assign layer_6[928] = far_6_7048_1[1]; 
    wire [1:0] far_6_7049_0;    relay_conn far_6_7049_0_a(.in(layer_5[782]), .out(far_6_7049_0[0]));    relay_conn far_6_7049_0_b(.in(layer_5[860]), .out(far_6_7049_0[1]));
    wire [1:0] far_6_7049_1;    relay_conn far_6_7049_1_a(.in(far_6_7049_0[0]), .out(far_6_7049_1[0]));    relay_conn far_6_7049_1_b(.in(far_6_7049_0[1]), .out(far_6_7049_1[1]));
    assign layer_6[929] = far_6_7049_1[1]; 
    assign layer_6[930] = ~(layer_5[745] & layer_5[750]); 
    wire [1:0] far_6_7051_0;    relay_conn far_6_7051_0_a(.in(layer_5[106]), .out(far_6_7051_0[0]));    relay_conn far_6_7051_0_b(.in(layer_5[234]), .out(far_6_7051_0[1]));
    wire [1:0] far_6_7051_1;    relay_conn far_6_7051_1_a(.in(far_6_7051_0[0]), .out(far_6_7051_1[0]));    relay_conn far_6_7051_1_b(.in(far_6_7051_0[1]), .out(far_6_7051_1[1]));
    wire [1:0] far_6_7051_2;    relay_conn far_6_7051_2_a(.in(far_6_7051_1[0]), .out(far_6_7051_2[0]));    relay_conn far_6_7051_2_b(.in(far_6_7051_1[1]), .out(far_6_7051_2[1]));
    wire [1:0] far_6_7051_3;    relay_conn far_6_7051_3_a(.in(far_6_7051_2[0]), .out(far_6_7051_3[0]));    relay_conn far_6_7051_3_b(.in(far_6_7051_2[1]), .out(far_6_7051_3[1]));
    assign layer_6[931] = far_6_7051_3[0] & far_6_7051_3[1]; 
    wire [1:0] far_6_7052_0;    relay_conn far_6_7052_0_a(.in(layer_5[366]), .out(far_6_7052_0[0]));    relay_conn far_6_7052_0_b(.in(layer_5[401]), .out(far_6_7052_0[1]));
    assign layer_6[932] = ~(far_6_7052_0[0] & far_6_7052_0[1]); 
    wire [1:0] far_6_7053_0;    relay_conn far_6_7053_0_a(.in(layer_5[63]), .out(far_6_7053_0[0]));    relay_conn far_6_7053_0_b(.in(layer_5[185]), .out(far_6_7053_0[1]));
    wire [1:0] far_6_7053_1;    relay_conn far_6_7053_1_a(.in(far_6_7053_0[0]), .out(far_6_7053_1[0]));    relay_conn far_6_7053_1_b(.in(far_6_7053_0[1]), .out(far_6_7053_1[1]));
    wire [1:0] far_6_7053_2;    relay_conn far_6_7053_2_a(.in(far_6_7053_1[0]), .out(far_6_7053_2[0]));    relay_conn far_6_7053_2_b(.in(far_6_7053_1[1]), .out(far_6_7053_2[1]));
    assign layer_6[933] = far_6_7053_2[0] & ~far_6_7053_2[1]; 
    assign layer_6[934] = layer_5[95]; 
    wire [1:0] far_6_7055_0;    relay_conn far_6_7055_0_a(.in(layer_5[912]), .out(far_6_7055_0[0]));    relay_conn far_6_7055_0_b(.in(layer_5[826]), .out(far_6_7055_0[1]));
    wire [1:0] far_6_7055_1;    relay_conn far_6_7055_1_a(.in(far_6_7055_0[0]), .out(far_6_7055_1[0]));    relay_conn far_6_7055_1_b(.in(far_6_7055_0[1]), .out(far_6_7055_1[1]));
    assign layer_6[935] = ~(far_6_7055_1[0] & far_6_7055_1[1]); 
    wire [1:0] far_6_7056_0;    relay_conn far_6_7056_0_a(.in(layer_5[697]), .out(far_6_7056_0[0]));    relay_conn far_6_7056_0_b(.in(layer_5[595]), .out(far_6_7056_0[1]));
    wire [1:0] far_6_7056_1;    relay_conn far_6_7056_1_a(.in(far_6_7056_0[0]), .out(far_6_7056_1[0]));    relay_conn far_6_7056_1_b(.in(far_6_7056_0[1]), .out(far_6_7056_1[1]));
    wire [1:0] far_6_7056_2;    relay_conn far_6_7056_2_a(.in(far_6_7056_1[0]), .out(far_6_7056_2[0]));    relay_conn far_6_7056_2_b(.in(far_6_7056_1[1]), .out(far_6_7056_2[1]));
    assign layer_6[936] = ~far_6_7056_2[1]; 
    wire [1:0] far_6_7057_0;    relay_conn far_6_7057_0_a(.in(layer_5[127]), .out(far_6_7057_0[0]));    relay_conn far_6_7057_0_b(.in(layer_5[179]), .out(far_6_7057_0[1]));
    assign layer_6[937] = ~far_6_7057_0[1] | (far_6_7057_0[0] & far_6_7057_0[1]); 
    wire [1:0] far_6_7058_0;    relay_conn far_6_7058_0_a(.in(layer_5[742]), .out(far_6_7058_0[0]));    relay_conn far_6_7058_0_b(.in(layer_5[774]), .out(far_6_7058_0[1]));
    assign layer_6[938] = far_6_7058_0[0] & far_6_7058_0[1]; 
    wire [1:0] far_6_7059_0;    relay_conn far_6_7059_0_a(.in(layer_5[92]), .out(far_6_7059_0[0]));    relay_conn far_6_7059_0_b(.in(layer_5[156]), .out(far_6_7059_0[1]));
    wire [1:0] far_6_7059_1;    relay_conn far_6_7059_1_a(.in(far_6_7059_0[0]), .out(far_6_7059_1[0]));    relay_conn far_6_7059_1_b(.in(far_6_7059_0[1]), .out(far_6_7059_1[1]));
    assign layer_6[939] = far_6_7059_1[1]; 
    wire [1:0] far_6_7060_0;    relay_conn far_6_7060_0_a(.in(layer_5[623]), .out(far_6_7060_0[0]));    relay_conn far_6_7060_0_b(.in(layer_5[562]), .out(far_6_7060_0[1]));
    assign layer_6[940] = far_6_7060_0[0] & ~far_6_7060_0[1]; 
    assign layer_6[941] = layer_5[717] & layer_5[734]; 
    wire [1:0] far_6_7062_0;    relay_conn far_6_7062_0_a(.in(layer_5[615]), .out(far_6_7062_0[0]));    relay_conn far_6_7062_0_b(.in(layer_5[648]), .out(far_6_7062_0[1]));
    assign layer_6[942] = ~far_6_7062_0[1]; 
    wire [1:0] far_6_7063_0;    relay_conn far_6_7063_0_a(.in(layer_5[972]), .out(far_6_7063_0[0]));    relay_conn far_6_7063_0_b(.in(layer_5[864]), .out(far_6_7063_0[1]));
    wire [1:0] far_6_7063_1;    relay_conn far_6_7063_1_a(.in(far_6_7063_0[0]), .out(far_6_7063_1[0]));    relay_conn far_6_7063_1_b(.in(far_6_7063_0[1]), .out(far_6_7063_1[1]));
    wire [1:0] far_6_7063_2;    relay_conn far_6_7063_2_a(.in(far_6_7063_1[0]), .out(far_6_7063_2[0]));    relay_conn far_6_7063_2_b(.in(far_6_7063_1[1]), .out(far_6_7063_2[1]));
    assign layer_6[943] = far_6_7063_2[0] | far_6_7063_2[1]; 
    wire [1:0] far_6_7064_0;    relay_conn far_6_7064_0_a(.in(layer_5[983]), .out(far_6_7064_0[0]));    relay_conn far_6_7064_0_b(.in(layer_5[900]), .out(far_6_7064_0[1]));
    wire [1:0] far_6_7064_1;    relay_conn far_6_7064_1_a(.in(far_6_7064_0[0]), .out(far_6_7064_1[0]));    relay_conn far_6_7064_1_b(.in(far_6_7064_0[1]), .out(far_6_7064_1[1]));
    assign layer_6[944] = ~far_6_7064_1[1] | (far_6_7064_1[0] & far_6_7064_1[1]); 
    wire [1:0] far_6_7065_0;    relay_conn far_6_7065_0_a(.in(layer_5[996]), .out(far_6_7065_0[0]));    relay_conn far_6_7065_0_b(.in(layer_5[939]), .out(far_6_7065_0[1]));
    assign layer_6[945] = ~(far_6_7065_0[0] & far_6_7065_0[1]); 
    wire [1:0] far_6_7066_0;    relay_conn far_6_7066_0_a(.in(layer_5[715]), .out(far_6_7066_0[0]));    relay_conn far_6_7066_0_b(.in(layer_5[660]), .out(far_6_7066_0[1]));
    assign layer_6[946] = far_6_7066_0[0] & far_6_7066_0[1]; 
    assign layer_6[947] = ~layer_5[863] | (layer_5[891] & layer_5[863]); 
    wire [1:0] far_6_7068_0;    relay_conn far_6_7068_0_a(.in(layer_5[860]), .out(far_6_7068_0[0]));    relay_conn far_6_7068_0_b(.in(layer_5[791]), .out(far_6_7068_0[1]));
    wire [1:0] far_6_7068_1;    relay_conn far_6_7068_1_a(.in(far_6_7068_0[0]), .out(far_6_7068_1[0]));    relay_conn far_6_7068_1_b(.in(far_6_7068_0[1]), .out(far_6_7068_1[1]));
    assign layer_6[948] = ~far_6_7068_1[0] | (far_6_7068_1[0] & far_6_7068_1[1]); 
    assign layer_6[949] = ~layer_5[69]; 
    wire [1:0] far_6_7070_0;    relay_conn far_6_7070_0_a(.in(layer_5[448]), .out(far_6_7070_0[0]));    relay_conn far_6_7070_0_b(.in(layer_5[489]), .out(far_6_7070_0[1]));
    assign layer_6[950] = ~far_6_7070_0[1]; 
    wire [1:0] far_6_7071_0;    relay_conn far_6_7071_0_a(.in(layer_5[364]), .out(far_6_7071_0[0]));    relay_conn far_6_7071_0_b(.in(layer_5[476]), .out(far_6_7071_0[1]));
    wire [1:0] far_6_7071_1;    relay_conn far_6_7071_1_a(.in(far_6_7071_0[0]), .out(far_6_7071_1[0]));    relay_conn far_6_7071_1_b(.in(far_6_7071_0[1]), .out(far_6_7071_1[1]));
    wire [1:0] far_6_7071_2;    relay_conn far_6_7071_2_a(.in(far_6_7071_1[0]), .out(far_6_7071_2[0]));    relay_conn far_6_7071_2_b(.in(far_6_7071_1[1]), .out(far_6_7071_2[1]));
    assign layer_6[951] = ~(far_6_7071_2[0] & far_6_7071_2[1]); 
    wire [1:0] far_6_7072_0;    relay_conn far_6_7072_0_a(.in(layer_5[433]), .out(far_6_7072_0[0]));    relay_conn far_6_7072_0_b(.in(layer_5[550]), .out(far_6_7072_0[1]));
    wire [1:0] far_6_7072_1;    relay_conn far_6_7072_1_a(.in(far_6_7072_0[0]), .out(far_6_7072_1[0]));    relay_conn far_6_7072_1_b(.in(far_6_7072_0[1]), .out(far_6_7072_1[1]));
    wire [1:0] far_6_7072_2;    relay_conn far_6_7072_2_a(.in(far_6_7072_1[0]), .out(far_6_7072_2[0]));    relay_conn far_6_7072_2_b(.in(far_6_7072_1[1]), .out(far_6_7072_2[1]));
    assign layer_6[952] = ~far_6_7072_2[0]; 
    wire [1:0] far_6_7073_0;    relay_conn far_6_7073_0_a(.in(layer_5[761]), .out(far_6_7073_0[0]));    relay_conn far_6_7073_0_b(.in(layer_5[801]), .out(far_6_7073_0[1]));
    assign layer_6[953] = ~far_6_7073_0[1]; 
    assign layer_6[954] = layer_5[791]; 
    wire [1:0] far_6_7075_0;    relay_conn far_6_7075_0_a(.in(layer_5[693]), .out(far_6_7075_0[0]));    relay_conn far_6_7075_0_b(.in(layer_5[766]), .out(far_6_7075_0[1]));
    wire [1:0] far_6_7075_1;    relay_conn far_6_7075_1_a(.in(far_6_7075_0[0]), .out(far_6_7075_1[0]));    relay_conn far_6_7075_1_b(.in(far_6_7075_0[1]), .out(far_6_7075_1[1]));
    assign layer_6[955] = ~far_6_7075_1[1] | (far_6_7075_1[0] & far_6_7075_1[1]); 
    assign layer_6[956] = ~(layer_5[613] | layer_5[639]); 
    wire [1:0] far_6_7077_0;    relay_conn far_6_7077_0_a(.in(layer_5[136]), .out(far_6_7077_0[0]));    relay_conn far_6_7077_0_b(.in(layer_5[35]), .out(far_6_7077_0[1]));
    wire [1:0] far_6_7077_1;    relay_conn far_6_7077_1_a(.in(far_6_7077_0[0]), .out(far_6_7077_1[0]));    relay_conn far_6_7077_1_b(.in(far_6_7077_0[1]), .out(far_6_7077_1[1]));
    wire [1:0] far_6_7077_2;    relay_conn far_6_7077_2_a(.in(far_6_7077_1[0]), .out(far_6_7077_2[0]));    relay_conn far_6_7077_2_b(.in(far_6_7077_1[1]), .out(far_6_7077_2[1]));
    assign layer_6[957] = far_6_7077_2[0] ^ far_6_7077_2[1]; 
    wire [1:0] far_6_7078_0;    relay_conn far_6_7078_0_a(.in(layer_5[612]), .out(far_6_7078_0[0]));    relay_conn far_6_7078_0_b(.in(layer_5[495]), .out(far_6_7078_0[1]));
    wire [1:0] far_6_7078_1;    relay_conn far_6_7078_1_a(.in(far_6_7078_0[0]), .out(far_6_7078_1[0]));    relay_conn far_6_7078_1_b(.in(far_6_7078_0[1]), .out(far_6_7078_1[1]));
    wire [1:0] far_6_7078_2;    relay_conn far_6_7078_2_a(.in(far_6_7078_1[0]), .out(far_6_7078_2[0]));    relay_conn far_6_7078_2_b(.in(far_6_7078_1[1]), .out(far_6_7078_2[1]));
    assign layer_6[958] = ~(far_6_7078_2[0] ^ far_6_7078_2[1]); 
    assign layer_6[959] = layer_5[455] & ~layer_5[449]; 
    wire [1:0] far_6_7080_0;    relay_conn far_6_7080_0_a(.in(layer_5[330]), .out(far_6_7080_0[0]));    relay_conn far_6_7080_0_b(.in(layer_5[391]), .out(far_6_7080_0[1]));
    assign layer_6[960] = ~(far_6_7080_0[0] | far_6_7080_0[1]); 
    wire [1:0] far_6_7081_0;    relay_conn far_6_7081_0_a(.in(layer_5[238]), .out(far_6_7081_0[0]));    relay_conn far_6_7081_0_b(.in(layer_5[111]), .out(far_6_7081_0[1]));
    wire [1:0] far_6_7081_1;    relay_conn far_6_7081_1_a(.in(far_6_7081_0[0]), .out(far_6_7081_1[0]));    relay_conn far_6_7081_1_b(.in(far_6_7081_0[1]), .out(far_6_7081_1[1]));
    wire [1:0] far_6_7081_2;    relay_conn far_6_7081_2_a(.in(far_6_7081_1[0]), .out(far_6_7081_2[0]));    relay_conn far_6_7081_2_b(.in(far_6_7081_1[1]), .out(far_6_7081_2[1]));
    assign layer_6[961] = ~far_6_7081_2[1]; 
    wire [1:0] far_6_7082_0;    relay_conn far_6_7082_0_a(.in(layer_5[256]), .out(far_6_7082_0[0]));    relay_conn far_6_7082_0_b(.in(layer_5[129]), .out(far_6_7082_0[1]));
    wire [1:0] far_6_7082_1;    relay_conn far_6_7082_1_a(.in(far_6_7082_0[0]), .out(far_6_7082_1[0]));    relay_conn far_6_7082_1_b(.in(far_6_7082_0[1]), .out(far_6_7082_1[1]));
    wire [1:0] far_6_7082_2;    relay_conn far_6_7082_2_a(.in(far_6_7082_1[0]), .out(far_6_7082_2[0]));    relay_conn far_6_7082_2_b(.in(far_6_7082_1[1]), .out(far_6_7082_2[1]));
    assign layer_6[962] = far_6_7082_2[0] & far_6_7082_2[1]; 
    wire [1:0] far_6_7083_0;    relay_conn far_6_7083_0_a(.in(layer_5[684]), .out(far_6_7083_0[0]));    relay_conn far_6_7083_0_b(.in(layer_5[801]), .out(far_6_7083_0[1]));
    wire [1:0] far_6_7083_1;    relay_conn far_6_7083_1_a(.in(far_6_7083_0[0]), .out(far_6_7083_1[0]));    relay_conn far_6_7083_1_b(.in(far_6_7083_0[1]), .out(far_6_7083_1[1]));
    wire [1:0] far_6_7083_2;    relay_conn far_6_7083_2_a(.in(far_6_7083_1[0]), .out(far_6_7083_2[0]));    relay_conn far_6_7083_2_b(.in(far_6_7083_1[1]), .out(far_6_7083_2[1]));
    assign layer_6[963] = ~far_6_7083_2[1] | (far_6_7083_2[0] & far_6_7083_2[1]); 
    wire [1:0] far_6_7084_0;    relay_conn far_6_7084_0_a(.in(layer_5[640]), .out(far_6_7084_0[0]));    relay_conn far_6_7084_0_b(.in(layer_5[689]), .out(far_6_7084_0[1]));
    assign layer_6[964] = ~(far_6_7084_0[0] & far_6_7084_0[1]); 
    wire [1:0] far_6_7085_0;    relay_conn far_6_7085_0_a(.in(layer_5[481]), .out(far_6_7085_0[0]));    relay_conn far_6_7085_0_b(.in(layer_5[368]), .out(far_6_7085_0[1]));
    wire [1:0] far_6_7085_1;    relay_conn far_6_7085_1_a(.in(far_6_7085_0[0]), .out(far_6_7085_1[0]));    relay_conn far_6_7085_1_b(.in(far_6_7085_0[1]), .out(far_6_7085_1[1]));
    wire [1:0] far_6_7085_2;    relay_conn far_6_7085_2_a(.in(far_6_7085_1[0]), .out(far_6_7085_2[0]));    relay_conn far_6_7085_2_b(.in(far_6_7085_1[1]), .out(far_6_7085_2[1]));
    assign layer_6[965] = far_6_7085_2[1]; 
    wire [1:0] far_6_7086_0;    relay_conn far_6_7086_0_a(.in(layer_5[720]), .out(far_6_7086_0[0]));    relay_conn far_6_7086_0_b(.in(layer_5[678]), .out(far_6_7086_0[1]));
    assign layer_6[966] = far_6_7086_0[0] ^ far_6_7086_0[1]; 
    assign layer_6[967] = layer_5[556] | layer_5[537]; 
    wire [1:0] far_6_7088_0;    relay_conn far_6_7088_0_a(.in(layer_5[310]), .out(far_6_7088_0[0]));    relay_conn far_6_7088_0_b(.in(layer_5[361]), .out(far_6_7088_0[1]));
    assign layer_6[968] = far_6_7088_0[1]; 
    wire [1:0] far_6_7089_0;    relay_conn far_6_7089_0_a(.in(layer_5[1005]), .out(far_6_7089_0[0]));    relay_conn far_6_7089_0_b(.in(layer_5[945]), .out(far_6_7089_0[1]));
    assign layer_6[969] = ~far_6_7089_0[1] | (far_6_7089_0[0] & far_6_7089_0[1]); 
    wire [1:0] far_6_7090_0;    relay_conn far_6_7090_0_a(.in(layer_5[613]), .out(far_6_7090_0[0]));    relay_conn far_6_7090_0_b(.in(layer_5[670]), .out(far_6_7090_0[1]));
    assign layer_6[970] = ~(far_6_7090_0[0] & far_6_7090_0[1]); 
    wire [1:0] far_6_7091_0;    relay_conn far_6_7091_0_a(.in(layer_5[885]), .out(far_6_7091_0[0]));    relay_conn far_6_7091_0_b(.in(layer_5[967]), .out(far_6_7091_0[1]));
    wire [1:0] far_6_7091_1;    relay_conn far_6_7091_1_a(.in(far_6_7091_0[0]), .out(far_6_7091_1[0]));    relay_conn far_6_7091_1_b(.in(far_6_7091_0[1]), .out(far_6_7091_1[1]));
    assign layer_6[971] = ~far_6_7091_1[1]; 
    wire [1:0] far_6_7092_0;    relay_conn far_6_7092_0_a(.in(layer_5[926]), .out(far_6_7092_0[0]));    relay_conn far_6_7092_0_b(.in(layer_5[845]), .out(far_6_7092_0[1]));
    wire [1:0] far_6_7092_1;    relay_conn far_6_7092_1_a(.in(far_6_7092_0[0]), .out(far_6_7092_1[0]));    relay_conn far_6_7092_1_b(.in(far_6_7092_0[1]), .out(far_6_7092_1[1]));
    assign layer_6[972] = far_6_7092_1[0]; 
    wire [1:0] far_6_7093_0;    relay_conn far_6_7093_0_a(.in(layer_5[83]), .out(far_6_7093_0[0]));    relay_conn far_6_7093_0_b(.in(layer_5[121]), .out(far_6_7093_0[1]));
    assign layer_6[973] = far_6_7093_0[0] ^ far_6_7093_0[1]; 
    wire [1:0] far_6_7094_0;    relay_conn far_6_7094_0_a(.in(layer_5[86]), .out(far_6_7094_0[0]));    relay_conn far_6_7094_0_b(.in(layer_5[196]), .out(far_6_7094_0[1]));
    wire [1:0] far_6_7094_1;    relay_conn far_6_7094_1_a(.in(far_6_7094_0[0]), .out(far_6_7094_1[0]));    relay_conn far_6_7094_1_b(.in(far_6_7094_0[1]), .out(far_6_7094_1[1]));
    wire [1:0] far_6_7094_2;    relay_conn far_6_7094_2_a(.in(far_6_7094_1[0]), .out(far_6_7094_2[0]));    relay_conn far_6_7094_2_b(.in(far_6_7094_1[1]), .out(far_6_7094_2[1]));
    assign layer_6[974] = far_6_7094_2[0] | far_6_7094_2[1]; 
    wire [1:0] far_6_7095_0;    relay_conn far_6_7095_0_a(.in(layer_5[761]), .out(far_6_7095_0[0]));    relay_conn far_6_7095_0_b(.in(layer_5[846]), .out(far_6_7095_0[1]));
    wire [1:0] far_6_7095_1;    relay_conn far_6_7095_1_a(.in(far_6_7095_0[0]), .out(far_6_7095_1[0]));    relay_conn far_6_7095_1_b(.in(far_6_7095_0[1]), .out(far_6_7095_1[1]));
    assign layer_6[975] = far_6_7095_1[1] & ~far_6_7095_1[0]; 
    wire [1:0] far_6_7096_0;    relay_conn far_6_7096_0_a(.in(layer_5[471]), .out(far_6_7096_0[0]));    relay_conn far_6_7096_0_b(.in(layer_5[364]), .out(far_6_7096_0[1]));
    wire [1:0] far_6_7096_1;    relay_conn far_6_7096_1_a(.in(far_6_7096_0[0]), .out(far_6_7096_1[0]));    relay_conn far_6_7096_1_b(.in(far_6_7096_0[1]), .out(far_6_7096_1[1]));
    wire [1:0] far_6_7096_2;    relay_conn far_6_7096_2_a(.in(far_6_7096_1[0]), .out(far_6_7096_2[0]));    relay_conn far_6_7096_2_b(.in(far_6_7096_1[1]), .out(far_6_7096_2[1]));
    assign layer_6[976] = far_6_7096_2[0] & far_6_7096_2[1]; 
    assign layer_6[977] = layer_5[216] & ~layer_5[238]; 
    wire [1:0] far_6_7098_0;    relay_conn far_6_7098_0_a(.in(layer_5[308]), .out(far_6_7098_0[0]));    relay_conn far_6_7098_0_b(.in(layer_5[430]), .out(far_6_7098_0[1]));
    wire [1:0] far_6_7098_1;    relay_conn far_6_7098_1_a(.in(far_6_7098_0[0]), .out(far_6_7098_1[0]));    relay_conn far_6_7098_1_b(.in(far_6_7098_0[1]), .out(far_6_7098_1[1]));
    wire [1:0] far_6_7098_2;    relay_conn far_6_7098_2_a(.in(far_6_7098_1[0]), .out(far_6_7098_2[0]));    relay_conn far_6_7098_2_b(.in(far_6_7098_1[1]), .out(far_6_7098_2[1]));
    assign layer_6[978] = far_6_7098_2[0] ^ far_6_7098_2[1]; 
    wire [1:0] far_6_7099_0;    relay_conn far_6_7099_0_a(.in(layer_5[949]), .out(far_6_7099_0[0]));    relay_conn far_6_7099_0_b(.in(layer_5[837]), .out(far_6_7099_0[1]));
    wire [1:0] far_6_7099_1;    relay_conn far_6_7099_1_a(.in(far_6_7099_0[0]), .out(far_6_7099_1[0]));    relay_conn far_6_7099_1_b(.in(far_6_7099_0[1]), .out(far_6_7099_1[1]));
    wire [1:0] far_6_7099_2;    relay_conn far_6_7099_2_a(.in(far_6_7099_1[0]), .out(far_6_7099_2[0]));    relay_conn far_6_7099_2_b(.in(far_6_7099_1[1]), .out(far_6_7099_2[1]));
    assign layer_6[979] = far_6_7099_2[0] & far_6_7099_2[1]; 
    wire [1:0] far_6_7100_0;    relay_conn far_6_7100_0_a(.in(layer_5[922]), .out(far_6_7100_0[0]));    relay_conn far_6_7100_0_b(.in(layer_5[886]), .out(far_6_7100_0[1]));
    assign layer_6[980] = ~far_6_7100_0[1] | (far_6_7100_0[0] & far_6_7100_0[1]); 
    wire [1:0] far_6_7101_0;    relay_conn far_6_7101_0_a(.in(layer_5[426]), .out(far_6_7101_0[0]));    relay_conn far_6_7101_0_b(.in(layer_5[504]), .out(far_6_7101_0[1]));
    wire [1:0] far_6_7101_1;    relay_conn far_6_7101_1_a(.in(far_6_7101_0[0]), .out(far_6_7101_1[0]));    relay_conn far_6_7101_1_b(.in(far_6_7101_0[1]), .out(far_6_7101_1[1]));
    assign layer_6[981] = ~far_6_7101_1[1] | (far_6_7101_1[0] & far_6_7101_1[1]); 
    wire [1:0] far_6_7102_0;    relay_conn far_6_7102_0_a(.in(layer_5[153]), .out(far_6_7102_0[0]));    relay_conn far_6_7102_0_b(.in(layer_5[115]), .out(far_6_7102_0[1]));
    assign layer_6[982] = far_6_7102_0[1] & ~far_6_7102_0[0]; 
    wire [1:0] far_6_7103_0;    relay_conn far_6_7103_0_a(.in(layer_5[194]), .out(far_6_7103_0[0]));    relay_conn far_6_7103_0_b(.in(layer_5[127]), .out(far_6_7103_0[1]));
    wire [1:0] far_6_7103_1;    relay_conn far_6_7103_1_a(.in(far_6_7103_0[0]), .out(far_6_7103_1[0]));    relay_conn far_6_7103_1_b(.in(far_6_7103_0[1]), .out(far_6_7103_1[1]));
    assign layer_6[983] = ~(far_6_7103_1[0] | far_6_7103_1[1]); 
    wire [1:0] far_6_7104_0;    relay_conn far_6_7104_0_a(.in(layer_5[651]), .out(far_6_7104_0[0]));    relay_conn far_6_7104_0_b(.in(layer_5[619]), .out(far_6_7104_0[1]));
    assign layer_6[984] = ~far_6_7104_0[0] | (far_6_7104_0[0] & far_6_7104_0[1]); 
    wire [1:0] far_6_7105_0;    relay_conn far_6_7105_0_a(.in(layer_5[426]), .out(far_6_7105_0[0]));    relay_conn far_6_7105_0_b(.in(layer_5[394]), .out(far_6_7105_0[1]));
    assign layer_6[985] = far_6_7105_0[0] & far_6_7105_0[1]; 
    wire [1:0] far_6_7106_0;    relay_conn far_6_7106_0_a(.in(layer_5[452]), .out(far_6_7106_0[0]));    relay_conn far_6_7106_0_b(.in(layer_5[381]), .out(far_6_7106_0[1]));
    wire [1:0] far_6_7106_1;    relay_conn far_6_7106_1_a(.in(far_6_7106_0[0]), .out(far_6_7106_1[0]));    relay_conn far_6_7106_1_b(.in(far_6_7106_0[1]), .out(far_6_7106_1[1]));
    assign layer_6[986] = ~far_6_7106_1[0]; 
    wire [1:0] far_6_7107_0;    relay_conn far_6_7107_0_a(.in(layer_5[795]), .out(far_6_7107_0[0]));    relay_conn far_6_7107_0_b(.in(layer_5[751]), .out(far_6_7107_0[1]));
    assign layer_6[987] = far_6_7107_0[0] | far_6_7107_0[1]; 
    wire [1:0] far_6_7108_0;    relay_conn far_6_7108_0_a(.in(layer_5[904]), .out(far_6_7108_0[0]));    relay_conn far_6_7108_0_b(.in(layer_5[974]), .out(far_6_7108_0[1]));
    wire [1:0] far_6_7108_1;    relay_conn far_6_7108_1_a(.in(far_6_7108_0[0]), .out(far_6_7108_1[0]));    relay_conn far_6_7108_1_b(.in(far_6_7108_0[1]), .out(far_6_7108_1[1]));
    assign layer_6[988] = far_6_7108_1[0] & far_6_7108_1[1]; 
    wire [1:0] far_6_7109_0;    relay_conn far_6_7109_0_a(.in(layer_5[430]), .out(far_6_7109_0[0]));    relay_conn far_6_7109_0_b(.in(layer_5[488]), .out(far_6_7109_0[1]));
    assign layer_6[989] = far_6_7109_0[0] & far_6_7109_0[1]; 
    wire [1:0] far_6_7110_0;    relay_conn far_6_7110_0_a(.in(layer_5[822]), .out(far_6_7110_0[0]));    relay_conn far_6_7110_0_b(.in(layer_5[948]), .out(far_6_7110_0[1]));
    wire [1:0] far_6_7110_1;    relay_conn far_6_7110_1_a(.in(far_6_7110_0[0]), .out(far_6_7110_1[0]));    relay_conn far_6_7110_1_b(.in(far_6_7110_0[1]), .out(far_6_7110_1[1]));
    wire [1:0] far_6_7110_2;    relay_conn far_6_7110_2_a(.in(far_6_7110_1[0]), .out(far_6_7110_2[0]));    relay_conn far_6_7110_2_b(.in(far_6_7110_1[1]), .out(far_6_7110_2[1]));
    assign layer_6[990] = ~far_6_7110_2[0]; 
    wire [1:0] far_6_7111_0;    relay_conn far_6_7111_0_a(.in(layer_5[471]), .out(far_6_7111_0[0]));    relay_conn far_6_7111_0_b(.in(layer_5[527]), .out(far_6_7111_0[1]));
    assign layer_6[991] = ~far_6_7111_0[0] | (far_6_7111_0[0] & far_6_7111_0[1]); 
    wire [1:0] far_6_7112_0;    relay_conn far_6_7112_0_a(.in(layer_5[396]), .out(far_6_7112_0[0]));    relay_conn far_6_7112_0_b(.in(layer_5[480]), .out(far_6_7112_0[1]));
    wire [1:0] far_6_7112_1;    relay_conn far_6_7112_1_a(.in(far_6_7112_0[0]), .out(far_6_7112_1[0]));    relay_conn far_6_7112_1_b(.in(far_6_7112_0[1]), .out(far_6_7112_1[1]));
    assign layer_6[992] = ~(far_6_7112_1[0] & far_6_7112_1[1]); 
    wire [1:0] far_6_7113_0;    relay_conn far_6_7113_0_a(.in(layer_5[720]), .out(far_6_7113_0[0]));    relay_conn far_6_7113_0_b(.in(layer_5[662]), .out(far_6_7113_0[1]));
    assign layer_6[993] = ~(far_6_7113_0[0] & far_6_7113_0[1]); 
    assign layer_6[994] = layer_5[656] ^ layer_5[673]; 
    wire [1:0] far_6_7115_0;    relay_conn far_6_7115_0_a(.in(layer_5[736]), .out(far_6_7115_0[0]));    relay_conn far_6_7115_0_b(.in(layer_5[849]), .out(far_6_7115_0[1]));
    wire [1:0] far_6_7115_1;    relay_conn far_6_7115_1_a(.in(far_6_7115_0[0]), .out(far_6_7115_1[0]));    relay_conn far_6_7115_1_b(.in(far_6_7115_0[1]), .out(far_6_7115_1[1]));
    wire [1:0] far_6_7115_2;    relay_conn far_6_7115_2_a(.in(far_6_7115_1[0]), .out(far_6_7115_2[0]));    relay_conn far_6_7115_2_b(.in(far_6_7115_1[1]), .out(far_6_7115_2[1]));
    assign layer_6[995] = far_6_7115_2[0]; 
    wire [1:0] far_6_7116_0;    relay_conn far_6_7116_0_a(.in(layer_5[521]), .out(far_6_7116_0[0]));    relay_conn far_6_7116_0_b(.in(layer_5[487]), .out(far_6_7116_0[1]));
    assign layer_6[996] = ~(far_6_7116_0[0] | far_6_7116_0[1]); 
    wire [1:0] far_6_7117_0;    relay_conn far_6_7117_0_a(.in(layer_5[746]), .out(far_6_7117_0[0]));    relay_conn far_6_7117_0_b(.in(layer_5[779]), .out(far_6_7117_0[1]));
    assign layer_6[997] = ~(far_6_7117_0[0] ^ far_6_7117_0[1]); 
    wire [1:0] far_6_7118_0;    relay_conn far_6_7118_0_a(.in(layer_5[430]), .out(far_6_7118_0[0]));    relay_conn far_6_7118_0_b(.in(layer_5[514]), .out(far_6_7118_0[1]));
    wire [1:0] far_6_7118_1;    relay_conn far_6_7118_1_a(.in(far_6_7118_0[0]), .out(far_6_7118_1[0]));    relay_conn far_6_7118_1_b(.in(far_6_7118_0[1]), .out(far_6_7118_1[1]));
    assign layer_6[998] = far_6_7118_1[0] | far_6_7118_1[1]; 
    wire [1:0] far_6_7119_0;    relay_conn far_6_7119_0_a(.in(layer_5[844]), .out(far_6_7119_0[0]));    relay_conn far_6_7119_0_b(.in(layer_5[760]), .out(far_6_7119_0[1]));
    wire [1:0] far_6_7119_1;    relay_conn far_6_7119_1_a(.in(far_6_7119_0[0]), .out(far_6_7119_1[0]));    relay_conn far_6_7119_1_b(.in(far_6_7119_0[1]), .out(far_6_7119_1[1]));
    assign layer_6[999] = ~(far_6_7119_1[0] & far_6_7119_1[1]); 
    wire [1:0] far_6_7120_0;    relay_conn far_6_7120_0_a(.in(layer_5[297]), .out(far_6_7120_0[0]));    relay_conn far_6_7120_0_b(.in(layer_5[368]), .out(far_6_7120_0[1]));
    wire [1:0] far_6_7120_1;    relay_conn far_6_7120_1_a(.in(far_6_7120_0[0]), .out(far_6_7120_1[0]));    relay_conn far_6_7120_1_b(.in(far_6_7120_0[1]), .out(far_6_7120_1[1]));
    assign layer_6[1000] = ~far_6_7120_1[1] | (far_6_7120_1[0] & far_6_7120_1[1]); 
    wire [1:0] far_6_7121_0;    relay_conn far_6_7121_0_a(.in(layer_5[466]), .out(far_6_7121_0[0]));    relay_conn far_6_7121_0_b(.in(layer_5[402]), .out(far_6_7121_0[1]));
    wire [1:0] far_6_7121_1;    relay_conn far_6_7121_1_a(.in(far_6_7121_0[0]), .out(far_6_7121_1[0]));    relay_conn far_6_7121_1_b(.in(far_6_7121_0[1]), .out(far_6_7121_1[1]));
    assign layer_6[1001] = ~far_6_7121_1[0] | (far_6_7121_1[0] & far_6_7121_1[1]); 
    wire [1:0] far_6_7122_0;    relay_conn far_6_7122_0_a(.in(layer_5[96]), .out(far_6_7122_0[0]));    relay_conn far_6_7122_0_b(.in(layer_5[64]), .out(far_6_7122_0[1]));
    assign layer_6[1002] = far_6_7122_0[0] & ~far_6_7122_0[1]; 
    wire [1:0] far_6_7123_0;    relay_conn far_6_7123_0_a(.in(layer_5[588]), .out(far_6_7123_0[0]));    relay_conn far_6_7123_0_b(.in(layer_5[553]), .out(far_6_7123_0[1]));
    assign layer_6[1003] = far_6_7123_0[0] & ~far_6_7123_0[1]; 
    assign layer_6[1004] = ~layer_5[753]; 
    wire [1:0] far_6_7125_0;    relay_conn far_6_7125_0_a(.in(layer_5[552]), .out(far_6_7125_0[0]));    relay_conn far_6_7125_0_b(.in(layer_5[640]), .out(far_6_7125_0[1]));
    wire [1:0] far_6_7125_1;    relay_conn far_6_7125_1_a(.in(far_6_7125_0[0]), .out(far_6_7125_1[0]));    relay_conn far_6_7125_1_b(.in(far_6_7125_0[1]), .out(far_6_7125_1[1]));
    assign layer_6[1005] = ~(far_6_7125_1[0] & far_6_7125_1[1]); 
    wire [1:0] far_6_7126_0;    relay_conn far_6_7126_0_a(.in(layer_5[952]), .out(far_6_7126_0[0]));    relay_conn far_6_7126_0_b(.in(layer_5[860]), .out(far_6_7126_0[1]));
    wire [1:0] far_6_7126_1;    relay_conn far_6_7126_1_a(.in(far_6_7126_0[0]), .out(far_6_7126_1[0]));    relay_conn far_6_7126_1_b(.in(far_6_7126_0[1]), .out(far_6_7126_1[1]));
    assign layer_6[1006] = far_6_7126_1[0] | far_6_7126_1[1]; 
    wire [1:0] far_6_7127_0;    relay_conn far_6_7127_0_a(.in(layer_5[216]), .out(far_6_7127_0[0]));    relay_conn far_6_7127_0_b(.in(layer_5[159]), .out(far_6_7127_0[1]));
    assign layer_6[1007] = far_6_7127_0[0] | far_6_7127_0[1]; 
    wire [1:0] far_6_7128_0;    relay_conn far_6_7128_0_a(.in(layer_5[224]), .out(far_6_7128_0[0]));    relay_conn far_6_7128_0_b(.in(layer_5[173]), .out(far_6_7128_0[1]));
    assign layer_6[1008] = ~(far_6_7128_0[0] | far_6_7128_0[1]); 
    wire [1:0] far_6_7129_0;    relay_conn far_6_7129_0_a(.in(layer_5[720]), .out(far_6_7129_0[0]));    relay_conn far_6_7129_0_b(.in(layer_5[753]), .out(far_6_7129_0[1]));
    assign layer_6[1009] = ~far_6_7129_0[1]; 
    wire [1:0] far_6_7130_0;    relay_conn far_6_7130_0_a(.in(layer_5[440]), .out(far_6_7130_0[0]));    relay_conn far_6_7130_0_b(.in(layer_5[521]), .out(far_6_7130_0[1]));
    wire [1:0] far_6_7130_1;    relay_conn far_6_7130_1_a(.in(far_6_7130_0[0]), .out(far_6_7130_1[0]));    relay_conn far_6_7130_1_b(.in(far_6_7130_0[1]), .out(far_6_7130_1[1]));
    assign layer_6[1010] = far_6_7130_1[0] | far_6_7130_1[1]; 
    wire [1:0] far_6_7131_0;    relay_conn far_6_7131_0_a(.in(layer_5[548]), .out(far_6_7131_0[0]));    relay_conn far_6_7131_0_b(.in(layer_5[505]), .out(far_6_7131_0[1]));
    assign layer_6[1011] = far_6_7131_0[1]; 
    assign layer_6[1012] = ~layer_5[86] | (layer_5[116] & layer_5[86]); 
    wire [1:0] far_6_7133_0;    relay_conn far_6_7133_0_a(.in(layer_5[391]), .out(far_6_7133_0[0]));    relay_conn far_6_7133_0_b(.in(layer_5[467]), .out(far_6_7133_0[1]));
    wire [1:0] far_6_7133_1;    relay_conn far_6_7133_1_a(.in(far_6_7133_0[0]), .out(far_6_7133_1[0]));    relay_conn far_6_7133_1_b(.in(far_6_7133_0[1]), .out(far_6_7133_1[1]));
    assign layer_6[1013] = ~(far_6_7133_1[0] ^ far_6_7133_1[1]); 
    wire [1:0] far_6_7134_0;    relay_conn far_6_7134_0_a(.in(layer_5[934]), .out(far_6_7134_0[0]));    relay_conn far_6_7134_0_b(.in(layer_5[968]), .out(far_6_7134_0[1]));
    assign layer_6[1014] = far_6_7134_0[0] & far_6_7134_0[1]; 
    wire [1:0] far_6_7135_0;    relay_conn far_6_7135_0_a(.in(layer_5[993]), .out(far_6_7135_0[0]));    relay_conn far_6_7135_0_b(.in(layer_5[901]), .out(far_6_7135_0[1]));
    wire [1:0] far_6_7135_1;    relay_conn far_6_7135_1_a(.in(far_6_7135_0[0]), .out(far_6_7135_1[0]));    relay_conn far_6_7135_1_b(.in(far_6_7135_0[1]), .out(far_6_7135_1[1]));
    assign layer_6[1015] = far_6_7135_1[0]; 
    wire [1:0] far_6_7136_0;    relay_conn far_6_7136_0_a(.in(layer_5[110]), .out(far_6_7136_0[0]));    relay_conn far_6_7136_0_b(.in(layer_5[169]), .out(far_6_7136_0[1]));
    assign layer_6[1016] = ~far_6_7136_0[0]; 
    wire [1:0] far_6_7137_0;    relay_conn far_6_7137_0_a(.in(layer_5[1019]), .out(far_6_7137_0[0]));    relay_conn far_6_7137_0_b(.in(layer_5[891]), .out(far_6_7137_0[1]));
    wire [1:0] far_6_7137_1;    relay_conn far_6_7137_1_a(.in(far_6_7137_0[0]), .out(far_6_7137_1[0]));    relay_conn far_6_7137_1_b(.in(far_6_7137_0[1]), .out(far_6_7137_1[1]));
    wire [1:0] far_6_7137_2;    relay_conn far_6_7137_2_a(.in(far_6_7137_1[0]), .out(far_6_7137_2[0]));    relay_conn far_6_7137_2_b(.in(far_6_7137_1[1]), .out(far_6_7137_2[1]));
    wire [1:0] far_6_7137_3;    relay_conn far_6_7137_3_a(.in(far_6_7137_2[0]), .out(far_6_7137_3[0]));    relay_conn far_6_7137_3_b(.in(far_6_7137_2[1]), .out(far_6_7137_3[1]));
    assign layer_6[1017] = far_6_7137_3[1]; 
    assign layer_6[1018] = ~layer_5[359]; 
    wire [1:0] far_6_7139_0;    relay_conn far_6_7139_0_a(.in(layer_5[390]), .out(far_6_7139_0[0]));    relay_conn far_6_7139_0_b(.in(layer_5[282]), .out(far_6_7139_0[1]));
    wire [1:0] far_6_7139_1;    relay_conn far_6_7139_1_a(.in(far_6_7139_0[0]), .out(far_6_7139_1[0]));    relay_conn far_6_7139_1_b(.in(far_6_7139_0[1]), .out(far_6_7139_1[1]));
    wire [1:0] far_6_7139_2;    relay_conn far_6_7139_2_a(.in(far_6_7139_1[0]), .out(far_6_7139_2[0]));    relay_conn far_6_7139_2_b(.in(far_6_7139_1[1]), .out(far_6_7139_2[1]));
    assign layer_6[1019] = far_6_7139_2[0] & far_6_7139_2[1]; 
    // Layer 7 ============================================================
    wire [1:0] far_7_7140_0;    relay_conn far_7_7140_0_a(.in(layer_6[906]), .out(far_7_7140_0[0]));    relay_conn far_7_7140_0_b(.in(layer_6[963]), .out(far_7_7140_0[1]));
    assign out[0] = ~far_7_7140_0[0]; 
    wire [1:0] far_7_7141_0;    relay_conn far_7_7141_0_a(.in(layer_6[913]), .out(far_7_7141_0[0]));    relay_conn far_7_7141_0_b(.in(layer_6[970]), .out(far_7_7141_0[1]));
    assign out[1] = far_7_7141_0[1] & ~far_7_7141_0[0]; 
    wire [1:0] far_7_7142_0;    relay_conn far_7_7142_0_a(.in(layer_6[30]), .out(far_7_7142_0[0]));    relay_conn far_7_7142_0_b(.in(layer_6[157]), .out(far_7_7142_0[1]));
    wire [1:0] far_7_7142_1;    relay_conn far_7_7142_1_a(.in(far_7_7142_0[0]), .out(far_7_7142_1[0]));    relay_conn far_7_7142_1_b(.in(far_7_7142_0[1]), .out(far_7_7142_1[1]));
    wire [1:0] far_7_7142_2;    relay_conn far_7_7142_2_a(.in(far_7_7142_1[0]), .out(far_7_7142_2[0]));    relay_conn far_7_7142_2_b(.in(far_7_7142_1[1]), .out(far_7_7142_2[1]));
    assign out[2] = ~far_7_7142_2[1]; 
    assign out[3] = ~layer_6[74]; 
    wire [1:0] far_7_7144_0;    relay_conn far_7_7144_0_a(.in(layer_6[750]), .out(far_7_7144_0[0]));    relay_conn far_7_7144_0_b(.in(layer_6[718]), .out(far_7_7144_0[1]));
    assign out[4] = far_7_7144_0[0]; 
    wire [1:0] far_7_7145_0;    relay_conn far_7_7145_0_a(.in(layer_6[360]), .out(far_7_7145_0[0]));    relay_conn far_7_7145_0_b(.in(layer_6[412]), .out(far_7_7145_0[1]));
    assign out[5] = far_7_7145_0[0] & far_7_7145_0[1]; 
    assign out[6] = ~layer_6[109]; 
    wire [1:0] far_7_7147_0;    relay_conn far_7_7147_0_a(.in(layer_6[374]), .out(far_7_7147_0[0]));    relay_conn far_7_7147_0_b(.in(layer_6[497]), .out(far_7_7147_0[1]));
    wire [1:0] far_7_7147_1;    relay_conn far_7_7147_1_a(.in(far_7_7147_0[0]), .out(far_7_7147_1[0]));    relay_conn far_7_7147_1_b(.in(far_7_7147_0[1]), .out(far_7_7147_1[1]));
    wire [1:0] far_7_7147_2;    relay_conn far_7_7147_2_a(.in(far_7_7147_1[0]), .out(far_7_7147_2[0]));    relay_conn far_7_7147_2_b(.in(far_7_7147_1[1]), .out(far_7_7147_2[1]));
    assign out[7] = far_7_7147_2[0] & far_7_7147_2[1]; 
    wire [1:0] far_7_7148_0;    relay_conn far_7_7148_0_a(.in(layer_6[464]), .out(far_7_7148_0[0]));    relay_conn far_7_7148_0_b(.in(layer_6[412]), .out(far_7_7148_0[1]));
    assign out[8] = far_7_7148_0[1]; 
    wire [1:0] far_7_7149_0;    relay_conn far_7_7149_0_a(.in(layer_6[404]), .out(far_7_7149_0[0]));    relay_conn far_7_7149_0_b(.in(layer_6[360]), .out(far_7_7149_0[1]));
    assign out[9] = far_7_7149_0[1] & ~far_7_7149_0[0]; 
    assign out[10] = layer_6[180]; 
    wire [1:0] far_7_7151_0;    relay_conn far_7_7151_0_a(.in(layer_6[109]), .out(far_7_7151_0[0]));    relay_conn far_7_7151_0_b(.in(layer_6[157]), .out(far_7_7151_0[1]));
    assign out[11] = ~(far_7_7151_0[0] | far_7_7151_0[1]); 
    wire [1:0] far_7_7152_0;    relay_conn far_7_7152_0_a(.in(layer_6[254]), .out(far_7_7152_0[0]));    relay_conn far_7_7152_0_b(.in(layer_6[157]), .out(far_7_7152_0[1]));
    wire [1:0] far_7_7152_1;    relay_conn far_7_7152_1_a(.in(far_7_7152_0[0]), .out(far_7_7152_1[0]));    relay_conn far_7_7152_1_b(.in(far_7_7152_0[1]), .out(far_7_7152_1[1]));
    wire [1:0] far_7_7152_2;    relay_conn far_7_7152_2_a(.in(far_7_7152_1[0]), .out(far_7_7152_2[0]));    relay_conn far_7_7152_2_b(.in(far_7_7152_1[1]), .out(far_7_7152_2[1]));
    assign out[12] = ~(far_7_7152_2[0] | far_7_7152_2[1]); 
    wire [1:0] far_7_7153_0;    relay_conn far_7_7153_0_a(.in(layer_6[261]), .out(far_7_7153_0[0]));    relay_conn far_7_7153_0_b(.in(layer_6[222]), .out(far_7_7153_0[1]));
    assign out[13] = far_7_7153_0[0] ^ far_7_7153_0[1]; 
    wire [1:0] far_7_7154_0;    relay_conn far_7_7154_0_a(.in(layer_6[686]), .out(far_7_7154_0[0]));    relay_conn far_7_7154_0_b(.in(layer_6[606]), .out(far_7_7154_0[1]));
    wire [1:0] far_7_7154_1;    relay_conn far_7_7154_1_a(.in(far_7_7154_0[0]), .out(far_7_7154_1[0]));    relay_conn far_7_7154_1_b(.in(far_7_7154_0[1]), .out(far_7_7154_1[1]));
    assign out[14] = ~far_7_7154_1[1]; 
    wire [1:0] far_7_7155_0;    relay_conn far_7_7155_0_a(.in(layer_6[672]), .out(far_7_7155_0[0]));    relay_conn far_7_7155_0_b(.in(layer_6[706]), .out(far_7_7155_0[1]));
    assign out[15] = ~(far_7_7155_0[0] ^ far_7_7155_0[1]); 
    assign out[16] = ~(layer_6[591] | layer_6[583]); 
    wire [1:0] far_7_7157_0;    relay_conn far_7_7157_0_a(.in(layer_6[575]), .out(far_7_7157_0[0]));    relay_conn far_7_7157_0_b(.in(layer_6[478]), .out(far_7_7157_0[1]));
    wire [1:0] far_7_7157_1;    relay_conn far_7_7157_1_a(.in(far_7_7157_0[0]), .out(far_7_7157_1[0]));    relay_conn far_7_7157_1_b(.in(far_7_7157_0[1]), .out(far_7_7157_1[1]));
    wire [1:0] far_7_7157_2;    relay_conn far_7_7157_2_a(.in(far_7_7157_1[0]), .out(far_7_7157_2[0]));    relay_conn far_7_7157_2_b(.in(far_7_7157_1[1]), .out(far_7_7157_2[1]));
    assign out[17] = far_7_7157_2[1] & ~far_7_7157_2[0]; 
    assign out[18] = layer_6[688] & layer_6[676]; 
    wire [1:0] far_7_7159_0;    relay_conn far_7_7159_0_a(.in(layer_6[904]), .out(far_7_7159_0[0]));    relay_conn far_7_7159_0_b(.in(layer_6[971]), .out(far_7_7159_0[1]));
    wire [1:0] far_7_7159_1;    relay_conn far_7_7159_1_a(.in(far_7_7159_0[0]), .out(far_7_7159_1[0]));    relay_conn far_7_7159_1_b(.in(far_7_7159_0[1]), .out(far_7_7159_1[1]));
    assign out[19] = ~far_7_7159_1[1] | (far_7_7159_1[0] & far_7_7159_1[1]); 
    assign out[20] = layer_6[510] ^ layer_6[512]; 
    wire [1:0] far_7_7161_0;    relay_conn far_7_7161_0_a(.in(layer_6[290]), .out(far_7_7161_0[0]));    relay_conn far_7_7161_0_b(.in(layer_6[392]), .out(far_7_7161_0[1]));
    wire [1:0] far_7_7161_1;    relay_conn far_7_7161_1_a(.in(far_7_7161_0[0]), .out(far_7_7161_1[0]));    relay_conn far_7_7161_1_b(.in(far_7_7161_0[1]), .out(far_7_7161_1[1]));
    wire [1:0] far_7_7161_2;    relay_conn far_7_7161_2_a(.in(far_7_7161_1[0]), .out(far_7_7161_2[0]));    relay_conn far_7_7161_2_b(.in(far_7_7161_1[1]), .out(far_7_7161_2[1]));
    assign out[21] = far_7_7161_2[0] & far_7_7161_2[1]; 
    assign out[22] = layer_6[394] & ~layer_6[404]; 
    assign out[23] = layer_6[920]; 
    assign out[24] = layer_6[789] & layer_6[777]; 
    wire [1:0] far_7_7165_0;    relay_conn far_7_7165_0_a(.in(layer_6[329]), .out(far_7_7165_0[0]));    relay_conn far_7_7165_0_b(.in(layer_6[404]), .out(far_7_7165_0[1]));
    wire [1:0] far_7_7165_1;    relay_conn far_7_7165_1_a(.in(far_7_7165_0[0]), .out(far_7_7165_1[0]));    relay_conn far_7_7165_1_b(.in(far_7_7165_0[1]), .out(far_7_7165_1[1]));
    assign out[25] = far_7_7165_1[0] ^ far_7_7165_1[1]; 
    assign out[26] = layer_6[4]; 
    wire [1:0] far_7_7167_0;    relay_conn far_7_7167_0_a(.in(layer_6[186]), .out(far_7_7167_0[0]));    relay_conn far_7_7167_0_b(.in(layer_6[109]), .out(far_7_7167_0[1]));
    wire [1:0] far_7_7167_1;    relay_conn far_7_7167_1_a(.in(far_7_7167_0[0]), .out(far_7_7167_1[0]));    relay_conn far_7_7167_1_b(.in(far_7_7167_0[1]), .out(far_7_7167_1[1]));
    assign out[27] = ~far_7_7167_1[1] | (far_7_7167_1[0] & far_7_7167_1[1]); 
    assign out[28] = layer_6[737] ^ layer_6[757]; 
    wire [1:0] far_7_7169_0;    relay_conn far_7_7169_0_a(.in(layer_6[368]), .out(far_7_7169_0[0]));    relay_conn far_7_7169_0_b(.in(layer_6[478]), .out(far_7_7169_0[1]));
    wire [1:0] far_7_7169_1;    relay_conn far_7_7169_1_a(.in(far_7_7169_0[0]), .out(far_7_7169_1[0]));    relay_conn far_7_7169_1_b(.in(far_7_7169_0[1]), .out(far_7_7169_1[1]));
    wire [1:0] far_7_7169_2;    relay_conn far_7_7169_2_a(.in(far_7_7169_1[0]), .out(far_7_7169_2[0]));    relay_conn far_7_7169_2_b(.in(far_7_7169_1[1]), .out(far_7_7169_2[1]));
    assign out[29] = far_7_7169_2[0] & far_7_7169_2[1]; 
    assign out[30] = layer_6[118]; 
    wire [1:0] far_7_7171_0;    relay_conn far_7_7171_0_a(.in(layer_6[942]), .out(far_7_7171_0[0]));    relay_conn far_7_7171_0_b(.in(layer_6[982]), .out(far_7_7171_0[1]));
    assign out[31] = far_7_7171_0[0] & ~far_7_7171_0[1]; 
    wire [1:0] far_7_7172_0;    relay_conn far_7_7172_0_a(.in(layer_6[53]), .out(far_7_7172_0[0]));    relay_conn far_7_7172_0_b(.in(layer_6[19]), .out(far_7_7172_0[1]));
    assign out[32] = far_7_7172_0[1] & ~far_7_7172_0[0]; 
    wire [1:0] far_7_7173_0;    relay_conn far_7_7173_0_a(.in(layer_6[201]), .out(far_7_7173_0[0]));    relay_conn far_7_7173_0_b(.in(layer_6[321]), .out(far_7_7173_0[1]));
    wire [1:0] far_7_7173_1;    relay_conn far_7_7173_1_a(.in(far_7_7173_0[0]), .out(far_7_7173_1[0]));    relay_conn far_7_7173_1_b(.in(far_7_7173_0[1]), .out(far_7_7173_1[1]));
    wire [1:0] far_7_7173_2;    relay_conn far_7_7173_2_a(.in(far_7_7173_1[0]), .out(far_7_7173_2[0]));    relay_conn far_7_7173_2_b(.in(far_7_7173_1[1]), .out(far_7_7173_2[1]));
    assign out[33] = ~far_7_7173_2[0]; 
    wire [1:0] far_7_7174_0;    relay_conn far_7_7174_0_a(.in(layer_6[548]), .out(far_7_7174_0[0]));    relay_conn far_7_7174_0_b(.in(layer_6[672]), .out(far_7_7174_0[1]));
    wire [1:0] far_7_7174_1;    relay_conn far_7_7174_1_a(.in(far_7_7174_0[0]), .out(far_7_7174_1[0]));    relay_conn far_7_7174_1_b(.in(far_7_7174_0[1]), .out(far_7_7174_1[1]));
    wire [1:0] far_7_7174_2;    relay_conn far_7_7174_2_a(.in(far_7_7174_1[0]), .out(far_7_7174_2[0]));    relay_conn far_7_7174_2_b(.in(far_7_7174_1[1]), .out(far_7_7174_2[1]));
    assign out[34] = ~far_7_7174_2[0] | (far_7_7174_2[0] & far_7_7174_2[1]); 
    wire [1:0] far_7_7175_0;    relay_conn far_7_7175_0_a(.in(layer_6[1011]), .out(far_7_7175_0[0]));    relay_conn far_7_7175_0_b(.in(layer_6[972]), .out(far_7_7175_0[1]));
    assign out[35] = ~far_7_7175_0[0]; 
    wire [1:0] far_7_7176_0;    relay_conn far_7_7176_0_a(.in(layer_6[629]), .out(far_7_7176_0[0]));    relay_conn far_7_7176_0_b(.in(layer_6[566]), .out(far_7_7176_0[1]));
    assign out[36] = ~far_7_7176_0[0] | (far_7_7176_0[0] & far_7_7176_0[1]); 
    assign out[37] = ~(layer_6[279] | layer_6[262]); 
    wire [1:0] far_7_7178_0;    relay_conn far_7_7178_0_a(.in(layer_6[944]), .out(far_7_7178_0[0]));    relay_conn far_7_7178_0_b(.in(layer_6[845]), .out(far_7_7178_0[1]));
    wire [1:0] far_7_7178_1;    relay_conn far_7_7178_1_a(.in(far_7_7178_0[0]), .out(far_7_7178_1[0]));    relay_conn far_7_7178_1_b(.in(far_7_7178_0[1]), .out(far_7_7178_1[1]));
    wire [1:0] far_7_7178_2;    relay_conn far_7_7178_2_a(.in(far_7_7178_1[0]), .out(far_7_7178_2[0]));    relay_conn far_7_7178_2_b(.in(far_7_7178_1[1]), .out(far_7_7178_2[1]));
    assign out[38] = ~(far_7_7178_2[0] ^ far_7_7178_2[1]); 
    wire [1:0] far_7_7179_0;    relay_conn far_7_7179_0_a(.in(layer_6[173]), .out(far_7_7179_0[0]));    relay_conn far_7_7179_0_b(.in(layer_6[212]), .out(far_7_7179_0[1]));
    assign out[39] = far_7_7179_0[1] & ~far_7_7179_0[0]; 
    assign out[40] = ~(layer_6[299] | layer_6[272]); 
    wire [1:0] far_7_7181_0;    relay_conn far_7_7181_0_a(.in(layer_6[471]), .out(far_7_7181_0[0]));    relay_conn far_7_7181_0_b(.in(layer_6[568]), .out(far_7_7181_0[1]));
    wire [1:0] far_7_7181_1;    relay_conn far_7_7181_1_a(.in(far_7_7181_0[0]), .out(far_7_7181_1[0]));    relay_conn far_7_7181_1_b(.in(far_7_7181_0[1]), .out(far_7_7181_1[1]));
    wire [1:0] far_7_7181_2;    relay_conn far_7_7181_2_a(.in(far_7_7181_1[0]), .out(far_7_7181_2[0]));    relay_conn far_7_7181_2_b(.in(far_7_7181_1[1]), .out(far_7_7181_2[1]));
    assign out[41] = far_7_7181_2[1]; 
    assign out[42] = ~layer_6[128]; 
    wire [1:0] far_7_7183_0;    relay_conn far_7_7183_0_a(.in(layer_6[1008]), .out(far_7_7183_0[0]));    relay_conn far_7_7183_0_b(.in(layer_6[941]), .out(far_7_7183_0[1]));
    wire [1:0] far_7_7183_1;    relay_conn far_7_7183_1_a(.in(far_7_7183_0[0]), .out(far_7_7183_1[0]));    relay_conn far_7_7183_1_b(.in(far_7_7183_0[1]), .out(far_7_7183_1[1]));
    assign out[43] = far_7_7183_1[0] & ~far_7_7183_1[1]; 
    wire [1:0] far_7_7184_0;    relay_conn far_7_7184_0_a(.in(layer_6[821]), .out(far_7_7184_0[0]));    relay_conn far_7_7184_0_b(.in(layer_6[942]), .out(far_7_7184_0[1]));
    wire [1:0] far_7_7184_1;    relay_conn far_7_7184_1_a(.in(far_7_7184_0[0]), .out(far_7_7184_1[0]));    relay_conn far_7_7184_1_b(.in(far_7_7184_0[1]), .out(far_7_7184_1[1]));
    wire [1:0] far_7_7184_2;    relay_conn far_7_7184_2_a(.in(far_7_7184_1[0]), .out(far_7_7184_2[0]));    relay_conn far_7_7184_2_b(.in(far_7_7184_1[1]), .out(far_7_7184_2[1]));
    assign out[44] = far_7_7184_2[1]; 
    wire [1:0] far_7_7185_0;    relay_conn far_7_7185_0_a(.in(layer_6[435]), .out(far_7_7185_0[0]));    relay_conn far_7_7185_0_b(.in(layer_6[549]), .out(far_7_7185_0[1]));
    wire [1:0] far_7_7185_1;    relay_conn far_7_7185_1_a(.in(far_7_7185_0[0]), .out(far_7_7185_1[0]));    relay_conn far_7_7185_1_b(.in(far_7_7185_0[1]), .out(far_7_7185_1[1]));
    wire [1:0] far_7_7185_2;    relay_conn far_7_7185_2_a(.in(far_7_7185_1[0]), .out(far_7_7185_2[0]));    relay_conn far_7_7185_2_b(.in(far_7_7185_1[1]), .out(far_7_7185_2[1]));
    assign out[45] = far_7_7185_2[1] & ~far_7_7185_2[0]; 
    wire [1:0] far_7_7186_0;    relay_conn far_7_7186_0_a(.in(layer_6[819]), .out(far_7_7186_0[0]));    relay_conn far_7_7186_0_b(.in(layer_6[718]), .out(far_7_7186_0[1]));
    wire [1:0] far_7_7186_1;    relay_conn far_7_7186_1_a(.in(far_7_7186_0[0]), .out(far_7_7186_1[0]));    relay_conn far_7_7186_1_b(.in(far_7_7186_0[1]), .out(far_7_7186_1[1]));
    wire [1:0] far_7_7186_2;    relay_conn far_7_7186_2_a(.in(far_7_7186_1[0]), .out(far_7_7186_2[0]));    relay_conn far_7_7186_2_b(.in(far_7_7186_1[1]), .out(far_7_7186_2[1]));
    assign out[46] = far_7_7186_2[0] | far_7_7186_2[1]; 
    wire [1:0] far_7_7187_0;    relay_conn far_7_7187_0_a(.in(layer_6[393]), .out(far_7_7187_0[0]));    relay_conn far_7_7187_0_b(.in(layer_6[478]), .out(far_7_7187_0[1]));
    wire [1:0] far_7_7187_1;    relay_conn far_7_7187_1_a(.in(far_7_7187_0[0]), .out(far_7_7187_1[0]));    relay_conn far_7_7187_1_b(.in(far_7_7187_0[1]), .out(far_7_7187_1[1]));
    assign out[47] = far_7_7187_1[1]; 
    wire [1:0] far_7_7188_0;    relay_conn far_7_7188_0_a(.in(layer_6[800]), .out(far_7_7188_0[0]));    relay_conn far_7_7188_0_b(.in(layer_6[765]), .out(far_7_7188_0[1]));
    assign out[48] = ~(far_7_7188_0[0] ^ far_7_7188_0[1]); 
    wire [1:0] far_7_7189_0;    relay_conn far_7_7189_0_a(.in(layer_6[194]), .out(far_7_7189_0[0]));    relay_conn far_7_7189_0_b(.in(layer_6[242]), .out(far_7_7189_0[1]));
    assign out[49] = far_7_7189_0[0] ^ far_7_7189_0[1]; 
    wire [1:0] far_7_7190_0;    relay_conn far_7_7190_0_a(.in(layer_6[659]), .out(far_7_7190_0[0]));    relay_conn far_7_7190_0_b(.in(layer_6[773]), .out(far_7_7190_0[1]));
    wire [1:0] far_7_7190_1;    relay_conn far_7_7190_1_a(.in(far_7_7190_0[0]), .out(far_7_7190_1[0]));    relay_conn far_7_7190_1_b(.in(far_7_7190_0[1]), .out(far_7_7190_1[1]));
    wire [1:0] far_7_7190_2;    relay_conn far_7_7190_2_a(.in(far_7_7190_1[0]), .out(far_7_7190_2[0]));    relay_conn far_7_7190_2_b(.in(far_7_7190_1[1]), .out(far_7_7190_2[1]));
    assign out[50] = ~(far_7_7190_2[0] | far_7_7190_2[1]); 
    wire [1:0] far_7_7191_0;    relay_conn far_7_7191_0_a(.in(layer_6[317]), .out(far_7_7191_0[0]));    relay_conn far_7_7191_0_b(.in(layer_6[387]), .out(far_7_7191_0[1]));
    wire [1:0] far_7_7191_1;    relay_conn far_7_7191_1_a(.in(far_7_7191_0[0]), .out(far_7_7191_1[0]));    relay_conn far_7_7191_1_b(.in(far_7_7191_0[1]), .out(far_7_7191_1[1]));
    assign out[51] = ~(far_7_7191_1[0] | far_7_7191_1[1]); 
    assign out[52] = ~layer_6[721]; 
    wire [1:0] far_7_7193_0;    relay_conn far_7_7193_0_a(.in(layer_6[272]), .out(far_7_7193_0[0]));    relay_conn far_7_7193_0_b(.in(layer_6[230]), .out(far_7_7193_0[1]));
    assign out[53] = far_7_7193_0[1] & ~far_7_7193_0[0]; 
    wire [1:0] far_7_7194_0;    relay_conn far_7_7194_0_a(.in(layer_6[614]), .out(far_7_7194_0[0]));    relay_conn far_7_7194_0_b(.in(layer_6[675]), .out(far_7_7194_0[1]));
    assign out[54] = ~(far_7_7194_0[0] ^ far_7_7194_0[1]); 
    wire [1:0] far_7_7195_0;    relay_conn far_7_7195_0_a(.in(layer_6[239]), .out(far_7_7195_0[0]));    relay_conn far_7_7195_0_b(.in(layer_6[197]), .out(far_7_7195_0[1]));
    assign out[55] = ~far_7_7195_0[1]; 
    wire [1:0] far_7_7196_0;    relay_conn far_7_7196_0_a(.in(layer_6[670]), .out(far_7_7196_0[0]));    relay_conn far_7_7196_0_b(.in(layer_6[542]), .out(far_7_7196_0[1]));
    wire [1:0] far_7_7196_1;    relay_conn far_7_7196_1_a(.in(far_7_7196_0[0]), .out(far_7_7196_1[0]));    relay_conn far_7_7196_1_b(.in(far_7_7196_0[1]), .out(far_7_7196_1[1]));
    wire [1:0] far_7_7196_2;    relay_conn far_7_7196_2_a(.in(far_7_7196_1[0]), .out(far_7_7196_2[0]));    relay_conn far_7_7196_2_b(.in(far_7_7196_1[1]), .out(far_7_7196_2[1]));
    wire [1:0] far_7_7196_3;    relay_conn far_7_7196_3_a(.in(far_7_7196_2[0]), .out(far_7_7196_3[0]));    relay_conn far_7_7196_3_b(.in(far_7_7196_2[1]), .out(far_7_7196_3[1]));
    assign out[56] = far_7_7196_3[0]; 
    wire [1:0] far_7_7197_0;    relay_conn far_7_7197_0_a(.in(layer_6[941]), .out(far_7_7197_0[0]));    relay_conn far_7_7197_0_b(.in(layer_6[828]), .out(far_7_7197_0[1]));
    wire [1:0] far_7_7197_1;    relay_conn far_7_7197_1_a(.in(far_7_7197_0[0]), .out(far_7_7197_1[0]));    relay_conn far_7_7197_1_b(.in(far_7_7197_0[1]), .out(far_7_7197_1[1]));
    wire [1:0] far_7_7197_2;    relay_conn far_7_7197_2_a(.in(far_7_7197_1[0]), .out(far_7_7197_2[0]));    relay_conn far_7_7197_2_b(.in(far_7_7197_1[1]), .out(far_7_7197_2[1]));
    assign out[57] = far_7_7197_2[1] & ~far_7_7197_2[0]; 
    wire [1:0] far_7_7198_0;    relay_conn far_7_7198_0_a(.in(layer_6[727]), .out(far_7_7198_0[0]));    relay_conn far_7_7198_0_b(.in(layer_6[599]), .out(far_7_7198_0[1]));
    wire [1:0] far_7_7198_1;    relay_conn far_7_7198_1_a(.in(far_7_7198_0[0]), .out(far_7_7198_1[0]));    relay_conn far_7_7198_1_b(.in(far_7_7198_0[1]), .out(far_7_7198_1[1]));
    wire [1:0] far_7_7198_2;    relay_conn far_7_7198_2_a(.in(far_7_7198_1[0]), .out(far_7_7198_2[0]));    relay_conn far_7_7198_2_b(.in(far_7_7198_1[1]), .out(far_7_7198_2[1]));
    wire [1:0] far_7_7198_3;    relay_conn far_7_7198_3_a(.in(far_7_7198_2[0]), .out(far_7_7198_3[0]));    relay_conn far_7_7198_3_b(.in(far_7_7198_2[1]), .out(far_7_7198_3[1]));
    assign out[58] = far_7_7198_3[0]; 
    wire [1:0] far_7_7199_0;    relay_conn far_7_7199_0_a(.in(layer_6[30]), .out(far_7_7199_0[0]));    relay_conn far_7_7199_0_b(.in(layer_6[103]), .out(far_7_7199_0[1]));
    wire [1:0] far_7_7199_1;    relay_conn far_7_7199_1_a(.in(far_7_7199_0[0]), .out(far_7_7199_1[0]));    relay_conn far_7_7199_1_b(.in(far_7_7199_0[1]), .out(far_7_7199_1[1]));
    assign out[59] = ~far_7_7199_1[1]; 
    wire [1:0] far_7_7200_0;    relay_conn far_7_7200_0_a(.in(layer_6[869]), .out(far_7_7200_0[0]));    relay_conn far_7_7200_0_b(.in(layer_6[831]), .out(far_7_7200_0[1]));
    assign out[60] = far_7_7200_0[1]; 
    wire [1:0] far_7_7201_0;    relay_conn far_7_7201_0_a(.in(layer_6[736]), .out(far_7_7201_0[0]));    relay_conn far_7_7201_0_b(.in(layer_6[670]), .out(far_7_7201_0[1]));
    wire [1:0] far_7_7201_1;    relay_conn far_7_7201_1_a(.in(far_7_7201_0[0]), .out(far_7_7201_1[0]));    relay_conn far_7_7201_1_b(.in(far_7_7201_0[1]), .out(far_7_7201_1[1]));
    assign out[61] = far_7_7201_1[0]; 
    wire [1:0] far_7_7202_0;    relay_conn far_7_7202_0_a(.in(layer_6[679]), .out(far_7_7202_0[0]));    relay_conn far_7_7202_0_b(.in(layer_6[631]), .out(far_7_7202_0[1]));
    assign out[62] = ~far_7_7202_0[1]; 
    assign out[63] = layer_6[153] & ~layer_6[139]; 
    wire [1:0] far_7_7204_0;    relay_conn far_7_7204_0_a(.in(layer_6[896]), .out(far_7_7204_0[0]));    relay_conn far_7_7204_0_b(.in(layer_6[825]), .out(far_7_7204_0[1]));
    wire [1:0] far_7_7204_1;    relay_conn far_7_7204_1_a(.in(far_7_7204_0[0]), .out(far_7_7204_1[0]));    relay_conn far_7_7204_1_b(.in(far_7_7204_0[1]), .out(far_7_7204_1[1]));
    assign out[64] = far_7_7204_1[0] | far_7_7204_1[1]; 
    wire [1:0] far_7_7205_0;    relay_conn far_7_7205_0_a(.in(layer_6[472]), .out(far_7_7205_0[0]));    relay_conn far_7_7205_0_b(.in(layer_6[556]), .out(far_7_7205_0[1]));
    wire [1:0] far_7_7205_1;    relay_conn far_7_7205_1_a(.in(far_7_7205_0[0]), .out(far_7_7205_1[0]));    relay_conn far_7_7205_1_b(.in(far_7_7205_0[1]), .out(far_7_7205_1[1]));
    assign out[65] = far_7_7205_1[0] & ~far_7_7205_1[1]; 
    wire [1:0] far_7_7206_0;    relay_conn far_7_7206_0_a(.in(layer_6[548]), .out(far_7_7206_0[0]));    relay_conn far_7_7206_0_b(.in(layer_6[437]), .out(far_7_7206_0[1]));
    wire [1:0] far_7_7206_1;    relay_conn far_7_7206_1_a(.in(far_7_7206_0[0]), .out(far_7_7206_1[0]));    relay_conn far_7_7206_1_b(.in(far_7_7206_0[1]), .out(far_7_7206_1[1]));
    wire [1:0] far_7_7206_2;    relay_conn far_7_7206_2_a(.in(far_7_7206_1[0]), .out(far_7_7206_2[0]));    relay_conn far_7_7206_2_b(.in(far_7_7206_1[1]), .out(far_7_7206_2[1]));
    assign out[66] = ~far_7_7206_2[0] | (far_7_7206_2[0] & far_7_7206_2[1]); 
    assign out[67] = layer_6[56] & ~layer_6[79]; 
    wire [1:0] far_7_7208_0;    relay_conn far_7_7208_0_a(.in(layer_6[129]), .out(far_7_7208_0[0]));    relay_conn far_7_7208_0_b(.in(layer_6[222]), .out(far_7_7208_0[1]));
    wire [1:0] far_7_7208_1;    relay_conn far_7_7208_1_a(.in(far_7_7208_0[0]), .out(far_7_7208_1[0]));    relay_conn far_7_7208_1_b(.in(far_7_7208_0[1]), .out(far_7_7208_1[1]));
    assign out[68] = far_7_7208_1[0]; 
    assign out[69] = layer_6[150] & ~layer_6[128]; 
    wire [1:0] far_7_7210_0;    relay_conn far_7_7210_0_a(.in(layer_6[660]), .out(far_7_7210_0[0]));    relay_conn far_7_7210_0_b(.in(layer_6[760]), .out(far_7_7210_0[1]));
    wire [1:0] far_7_7210_1;    relay_conn far_7_7210_1_a(.in(far_7_7210_0[0]), .out(far_7_7210_1[0]));    relay_conn far_7_7210_1_b(.in(far_7_7210_0[1]), .out(far_7_7210_1[1]));
    wire [1:0] far_7_7210_2;    relay_conn far_7_7210_2_a(.in(far_7_7210_1[0]), .out(far_7_7210_2[0]));    relay_conn far_7_7210_2_b(.in(far_7_7210_1[1]), .out(far_7_7210_2[1]));
    assign out[70] = far_7_7210_2[1] & ~far_7_7210_2[0]; 
    assign out[71] = layer_6[775]; 
    wire [1:0] far_7_7212_0;    relay_conn far_7_7212_0_a(.in(layer_6[888]), .out(far_7_7212_0[0]));    relay_conn far_7_7212_0_b(.in(layer_6[987]), .out(far_7_7212_0[1]));
    wire [1:0] far_7_7212_1;    relay_conn far_7_7212_1_a(.in(far_7_7212_0[0]), .out(far_7_7212_1[0]));    relay_conn far_7_7212_1_b(.in(far_7_7212_0[1]), .out(far_7_7212_1[1]));
    wire [1:0] far_7_7212_2;    relay_conn far_7_7212_2_a(.in(far_7_7212_1[0]), .out(far_7_7212_2[0]));    relay_conn far_7_7212_2_b(.in(far_7_7212_1[1]), .out(far_7_7212_2[1]));
    assign out[72] = far_7_7212_2[0] & far_7_7212_2[1]; 
    assign out[73] = ~(layer_6[116] | layer_6[103]); 
    wire [1:0] far_7_7214_0;    relay_conn far_7_7214_0_a(.in(layer_6[421]), .out(far_7_7214_0[0]));    relay_conn far_7_7214_0_b(.in(layer_6[497]), .out(far_7_7214_0[1]));
    wire [1:0] far_7_7214_1;    relay_conn far_7_7214_1_a(.in(far_7_7214_0[0]), .out(far_7_7214_1[0]));    relay_conn far_7_7214_1_b(.in(far_7_7214_0[1]), .out(far_7_7214_1[1]));
    assign out[74] = far_7_7214_1[1] & ~far_7_7214_1[0]; 
    wire [1:0] far_7_7215_0;    relay_conn far_7_7215_0_a(.in(layer_6[972]), .out(far_7_7215_0[0]));    relay_conn far_7_7215_0_b(.in(layer_6[1016]), .out(far_7_7215_0[1]));
    assign out[75] = far_7_7215_0[0] & far_7_7215_0[1]; 
    assign out[76] = layer_6[944] ^ layer_6[941]; 
    wire [1:0] far_7_7217_0;    relay_conn far_7_7217_0_a(.in(layer_6[249]), .out(far_7_7217_0[0]));    relay_conn far_7_7217_0_b(.in(layer_6[316]), .out(far_7_7217_0[1]));
    wire [1:0] far_7_7217_1;    relay_conn far_7_7217_1_a(.in(far_7_7217_0[0]), .out(far_7_7217_1[0]));    relay_conn far_7_7217_1_b(.in(far_7_7217_0[1]), .out(far_7_7217_1[1]));
    assign out[77] = far_7_7217_1[0] ^ far_7_7217_1[1]; 
    wire [1:0] far_7_7218_0;    relay_conn far_7_7218_0_a(.in(layer_6[576]), .out(far_7_7218_0[0]));    relay_conn far_7_7218_0_b(.in(layer_6[537]), .out(far_7_7218_0[1]));
    assign out[78] = ~far_7_7218_0[0]; 
    wire [1:0] far_7_7219_0;    relay_conn far_7_7219_0_a(.in(layer_6[434]), .out(far_7_7219_0[0]));    relay_conn far_7_7219_0_b(.in(layer_6[511]), .out(far_7_7219_0[1]));
    wire [1:0] far_7_7219_1;    relay_conn far_7_7219_1_a(.in(far_7_7219_0[0]), .out(far_7_7219_1[0]));    relay_conn far_7_7219_1_b(.in(far_7_7219_0[1]), .out(far_7_7219_1[1]));
    assign out[79] = far_7_7219_1[0] & ~far_7_7219_1[1]; 
    wire [1:0] far_7_7220_0;    relay_conn far_7_7220_0_a(.in(layer_6[575]), .out(far_7_7220_0[0]));    relay_conn far_7_7220_0_b(.in(layer_6[615]), .out(far_7_7220_0[1]));
    assign out[80] = ~far_7_7220_0[0]; 
    assign out[81] = ~layer_6[198]; 
    wire [1:0] far_7_7222_0;    relay_conn far_7_7222_0_a(.in(layer_6[456]), .out(far_7_7222_0[0]));    relay_conn far_7_7222_0_b(.in(layer_6[558]), .out(far_7_7222_0[1]));
    wire [1:0] far_7_7222_1;    relay_conn far_7_7222_1_a(.in(far_7_7222_0[0]), .out(far_7_7222_1[0]));    relay_conn far_7_7222_1_b(.in(far_7_7222_0[1]), .out(far_7_7222_1[1]));
    wire [1:0] far_7_7222_2;    relay_conn far_7_7222_2_a(.in(far_7_7222_1[0]), .out(far_7_7222_2[0]));    relay_conn far_7_7222_2_b(.in(far_7_7222_1[1]), .out(far_7_7222_2[1]));
    assign out[82] = far_7_7222_2[1]; 
    wire [1:0] far_7_7223_0;    relay_conn far_7_7223_0_a(.in(layer_6[752]), .out(far_7_7223_0[0]));    relay_conn far_7_7223_0_b(.in(layer_6[792]), .out(far_7_7223_0[1]));
    assign out[83] = far_7_7223_0[0]; 
    wire [1:0] far_7_7224_0;    relay_conn far_7_7224_0_a(.in(layer_6[644]), .out(far_7_7224_0[0]));    relay_conn far_7_7224_0_b(.in(layer_6[599]), .out(far_7_7224_0[1]));
    assign out[84] = far_7_7224_0[0] & ~far_7_7224_0[1]; 
    wire [1:0] far_7_7225_0;    relay_conn far_7_7225_0_a(.in(layer_6[280]), .out(far_7_7225_0[0]));    relay_conn far_7_7225_0_b(.in(layer_6[338]), .out(far_7_7225_0[1]));
    assign out[85] = ~(far_7_7225_0[0] | far_7_7225_0[1]); 
    wire [1:0] far_7_7226_0;    relay_conn far_7_7226_0_a(.in(layer_6[363]), .out(far_7_7226_0[0]));    relay_conn far_7_7226_0_b(.in(layer_6[469]), .out(far_7_7226_0[1]));
    wire [1:0] far_7_7226_1;    relay_conn far_7_7226_1_a(.in(far_7_7226_0[0]), .out(far_7_7226_1[0]));    relay_conn far_7_7226_1_b(.in(far_7_7226_0[1]), .out(far_7_7226_1[1]));
    wire [1:0] far_7_7226_2;    relay_conn far_7_7226_2_a(.in(far_7_7226_1[0]), .out(far_7_7226_2[0]));    relay_conn far_7_7226_2_b(.in(far_7_7226_1[1]), .out(far_7_7226_2[1]));
    assign out[86] = ~far_7_7226_2[1]; 
    wire [1:0] far_7_7227_0;    relay_conn far_7_7227_0_a(.in(layer_6[404]), .out(far_7_7227_0[0]));    relay_conn far_7_7227_0_b(.in(layer_6[310]), .out(far_7_7227_0[1]));
    wire [1:0] far_7_7227_1;    relay_conn far_7_7227_1_a(.in(far_7_7227_0[0]), .out(far_7_7227_1[0]));    relay_conn far_7_7227_1_b(.in(far_7_7227_0[1]), .out(far_7_7227_1[1]));
    assign out[87] = ~(far_7_7227_1[0] | far_7_7227_1[1]); 
    wire [1:0] far_7_7228_0;    relay_conn far_7_7228_0_a(.in(layer_6[632]), .out(far_7_7228_0[0]));    relay_conn far_7_7228_0_b(.in(layer_6[730]), .out(far_7_7228_0[1]));
    wire [1:0] far_7_7228_1;    relay_conn far_7_7228_1_a(.in(far_7_7228_0[0]), .out(far_7_7228_1[0]));    relay_conn far_7_7228_1_b(.in(far_7_7228_0[1]), .out(far_7_7228_1[1]));
    wire [1:0] far_7_7228_2;    relay_conn far_7_7228_2_a(.in(far_7_7228_1[0]), .out(far_7_7228_2[0]));    relay_conn far_7_7228_2_b(.in(far_7_7228_1[1]), .out(far_7_7228_2[1]));
    assign out[88] = ~far_7_7228_2[1]; 
    wire [1:0] far_7_7229_0;    relay_conn far_7_7229_0_a(.in(layer_6[21]), .out(far_7_7229_0[0]));    relay_conn far_7_7229_0_b(.in(layer_6[105]), .out(far_7_7229_0[1]));
    wire [1:0] far_7_7229_1;    relay_conn far_7_7229_1_a(.in(far_7_7229_0[0]), .out(far_7_7229_1[0]));    relay_conn far_7_7229_1_b(.in(far_7_7229_0[1]), .out(far_7_7229_1[1]));
    assign out[89] = ~(far_7_7229_1[0] | far_7_7229_1[1]); 
    assign out[90] = layer_6[118] ^ layer_6[141]; 
    wire [1:0] far_7_7231_0;    relay_conn far_7_7231_0_a(.in(layer_6[203]), .out(far_7_7231_0[0]));    relay_conn far_7_7231_0_b(.in(layer_6[312]), .out(far_7_7231_0[1]));
    wire [1:0] far_7_7231_1;    relay_conn far_7_7231_1_a(.in(far_7_7231_0[0]), .out(far_7_7231_1[0]));    relay_conn far_7_7231_1_b(.in(far_7_7231_0[1]), .out(far_7_7231_1[1]));
    wire [1:0] far_7_7231_2;    relay_conn far_7_7231_2_a(.in(far_7_7231_1[0]), .out(far_7_7231_2[0]));    relay_conn far_7_7231_2_b(.in(far_7_7231_1[1]), .out(far_7_7231_2[1]));
    assign out[91] = ~(far_7_7231_2[0] | far_7_7231_2[1]); 
    assign out[92] = ~layer_6[173]; 
    wire [1:0] far_7_7233_0;    relay_conn far_7_7233_0_a(.in(layer_6[253]), .out(far_7_7233_0[0]));    relay_conn far_7_7233_0_b(.in(layer_6[361]), .out(far_7_7233_0[1]));
    wire [1:0] far_7_7233_1;    relay_conn far_7_7233_1_a(.in(far_7_7233_0[0]), .out(far_7_7233_1[0]));    relay_conn far_7_7233_1_b(.in(far_7_7233_0[1]), .out(far_7_7233_1[1]));
    wire [1:0] far_7_7233_2;    relay_conn far_7_7233_2_a(.in(far_7_7233_1[0]), .out(far_7_7233_2[0]));    relay_conn far_7_7233_2_b(.in(far_7_7233_1[1]), .out(far_7_7233_2[1]));
    assign out[93] = far_7_7233_2[0] & far_7_7233_2[1]; 
    wire [1:0] far_7_7234_0;    relay_conn far_7_7234_0_a(.in(layer_6[511]), .out(far_7_7234_0[0]));    relay_conn far_7_7234_0_b(.in(layer_6[453]), .out(far_7_7234_0[1]));
    assign out[94] = far_7_7234_0[1] & ~far_7_7234_0[0]; 
    wire [1:0] far_7_7235_0;    relay_conn far_7_7235_0_a(.in(layer_6[270]), .out(far_7_7235_0[0]));    relay_conn far_7_7235_0_b(.in(layer_6[184]), .out(far_7_7235_0[1]));
    wire [1:0] far_7_7235_1;    relay_conn far_7_7235_1_a(.in(far_7_7235_0[0]), .out(far_7_7235_1[0]));    relay_conn far_7_7235_1_b(.in(far_7_7235_0[1]), .out(far_7_7235_1[1]));
    assign out[95] = far_7_7235_1[0]; 
    wire [1:0] far_7_7236_0;    relay_conn far_7_7236_0_a(.in(layer_6[785]), .out(far_7_7236_0[0]));    relay_conn far_7_7236_0_b(.in(layer_6[753]), .out(far_7_7236_0[1]));
    assign out[96] = far_7_7236_0[0] & far_7_7236_0[1]; 
    assign out[97] = layer_6[1008]; 
    wire [1:0] far_7_7238_0;    relay_conn far_7_7238_0_a(.in(layer_6[374]), .out(far_7_7238_0[0]));    relay_conn far_7_7238_0_b(.in(layer_6[491]), .out(far_7_7238_0[1]));
    wire [1:0] far_7_7238_1;    relay_conn far_7_7238_1_a(.in(far_7_7238_0[0]), .out(far_7_7238_1[0]));    relay_conn far_7_7238_1_b(.in(far_7_7238_0[1]), .out(far_7_7238_1[1]));
    wire [1:0] far_7_7238_2;    relay_conn far_7_7238_2_a(.in(far_7_7238_1[0]), .out(far_7_7238_2[0]));    relay_conn far_7_7238_2_b(.in(far_7_7238_1[1]), .out(far_7_7238_2[1]));
    assign out[98] = ~(far_7_7238_2[0] ^ far_7_7238_2[1]); 
    wire [1:0] far_7_7239_0;    relay_conn far_7_7239_0_a(.in(layer_6[157]), .out(far_7_7239_0[0]));    relay_conn far_7_7239_0_b(.in(layer_6[75]), .out(far_7_7239_0[1]));
    wire [1:0] far_7_7239_1;    relay_conn far_7_7239_1_a(.in(far_7_7239_0[0]), .out(far_7_7239_1[0]));    relay_conn far_7_7239_1_b(.in(far_7_7239_0[1]), .out(far_7_7239_1[1]));
    assign out[99] = far_7_7239_1[1]; 
    assign out[100] = ~(layer_6[981] | layer_6[1011]); 
    wire [1:0] far_7_7241_0;    relay_conn far_7_7241_0_a(.in(layer_6[117]), .out(far_7_7241_0[0]));    relay_conn far_7_7241_0_b(.in(layer_6[44]), .out(far_7_7241_0[1]));
    wire [1:0] far_7_7241_1;    relay_conn far_7_7241_1_a(.in(far_7_7241_0[0]), .out(far_7_7241_1[0]));    relay_conn far_7_7241_1_b(.in(far_7_7241_0[1]), .out(far_7_7241_1[1]));
    assign out[101] = far_7_7241_1[0] | far_7_7241_1[1]; 
    wire [1:0] far_7_7242_0;    relay_conn far_7_7242_0_a(.in(layer_6[881]), .out(far_7_7242_0[0]));    relay_conn far_7_7242_0_b(.in(layer_6[931]), .out(far_7_7242_0[1]));
    assign out[102] = ~far_7_7242_0[1]; 
    wire [1:0] far_7_7243_0;    relay_conn far_7_7243_0_a(.in(layer_6[17]), .out(far_7_7243_0[0]));    relay_conn far_7_7243_0_b(.in(layer_6[139]), .out(far_7_7243_0[1]));
    wire [1:0] far_7_7243_1;    relay_conn far_7_7243_1_a(.in(far_7_7243_0[0]), .out(far_7_7243_1[0]));    relay_conn far_7_7243_1_b(.in(far_7_7243_0[1]), .out(far_7_7243_1[1]));
    wire [1:0] far_7_7243_2;    relay_conn far_7_7243_2_a(.in(far_7_7243_1[0]), .out(far_7_7243_2[0]));    relay_conn far_7_7243_2_b(.in(far_7_7243_1[1]), .out(far_7_7243_2[1]));
    assign out[103] = ~far_7_7243_2[0] | (far_7_7243_2[0] & far_7_7243_2[1]); 
    assign out[104] = layer_6[681] | layer_6[668]; 
    wire [1:0] far_7_7245_0;    relay_conn far_7_7245_0_a(.in(layer_6[632]), .out(far_7_7245_0[0]));    relay_conn far_7_7245_0_b(.in(layer_6[681]), .out(far_7_7245_0[1]));
    assign out[105] = ~(far_7_7245_0[0] ^ far_7_7245_0[1]); 
    assign out[106] = ~(layer_6[513] | layer_6[503]); 
    wire [1:0] far_7_7247_0;    relay_conn far_7_7247_0_a(.in(layer_6[470]), .out(far_7_7247_0[0]));    relay_conn far_7_7247_0_b(.in(layer_6[350]), .out(far_7_7247_0[1]));
    wire [1:0] far_7_7247_1;    relay_conn far_7_7247_1_a(.in(far_7_7247_0[0]), .out(far_7_7247_1[0]));    relay_conn far_7_7247_1_b(.in(far_7_7247_0[1]), .out(far_7_7247_1[1]));
    wire [1:0] far_7_7247_2;    relay_conn far_7_7247_2_a(.in(far_7_7247_1[0]), .out(far_7_7247_2[0]));    relay_conn far_7_7247_2_b(.in(far_7_7247_1[1]), .out(far_7_7247_2[1]));
    assign out[107] = ~far_7_7247_2[1]; 
    wire [1:0] far_7_7248_0;    relay_conn far_7_7248_0_a(.in(layer_6[406]), .out(far_7_7248_0[0]));    relay_conn far_7_7248_0_b(.in(layer_6[478]), .out(far_7_7248_0[1]));
    wire [1:0] far_7_7248_1;    relay_conn far_7_7248_1_a(.in(far_7_7248_0[0]), .out(far_7_7248_1[0]));    relay_conn far_7_7248_1_b(.in(far_7_7248_0[1]), .out(far_7_7248_1[1]));
    assign out[108] = far_7_7248_1[0] & ~far_7_7248_1[1]; 
    wire [1:0] far_7_7249_0;    relay_conn far_7_7249_0_a(.in(layer_6[700]), .out(far_7_7249_0[0]));    relay_conn far_7_7249_0_b(.in(layer_6[581]), .out(far_7_7249_0[1]));
    wire [1:0] far_7_7249_1;    relay_conn far_7_7249_1_a(.in(far_7_7249_0[0]), .out(far_7_7249_1[0]));    relay_conn far_7_7249_1_b(.in(far_7_7249_0[1]), .out(far_7_7249_1[1]));
    wire [1:0] far_7_7249_2;    relay_conn far_7_7249_2_a(.in(far_7_7249_1[0]), .out(far_7_7249_2[0]));    relay_conn far_7_7249_2_b(.in(far_7_7249_1[1]), .out(far_7_7249_2[1]));
    assign out[109] = far_7_7249_2[0] & ~far_7_7249_2[1]; 
    wire [1:0] far_7_7250_0;    relay_conn far_7_7250_0_a(.in(layer_6[447]), .out(far_7_7250_0[0]));    relay_conn far_7_7250_0_b(.in(layer_6[558]), .out(far_7_7250_0[1]));
    wire [1:0] far_7_7250_1;    relay_conn far_7_7250_1_a(.in(far_7_7250_0[0]), .out(far_7_7250_1[0]));    relay_conn far_7_7250_1_b(.in(far_7_7250_0[1]), .out(far_7_7250_1[1]));
    wire [1:0] far_7_7250_2;    relay_conn far_7_7250_2_a(.in(far_7_7250_1[0]), .out(far_7_7250_2[0]));    relay_conn far_7_7250_2_b(.in(far_7_7250_1[1]), .out(far_7_7250_2[1]));
    assign out[110] = ~(far_7_7250_2[0] & far_7_7250_2[1]); 
    wire [1:0] far_7_7251_0;    relay_conn far_7_7251_0_a(.in(layer_6[835]), .out(far_7_7251_0[0]));    relay_conn far_7_7251_0_b(.in(layer_6[952]), .out(far_7_7251_0[1]));
    wire [1:0] far_7_7251_1;    relay_conn far_7_7251_1_a(.in(far_7_7251_0[0]), .out(far_7_7251_1[0]));    relay_conn far_7_7251_1_b(.in(far_7_7251_0[1]), .out(far_7_7251_1[1]));
    wire [1:0] far_7_7251_2;    relay_conn far_7_7251_2_a(.in(far_7_7251_1[0]), .out(far_7_7251_2[0]));    relay_conn far_7_7251_2_b(.in(far_7_7251_1[1]), .out(far_7_7251_2[1]));
    assign out[111] = far_7_7251_2[0] | far_7_7251_2[1]; 
    assign out[112] = layer_6[681] | layer_6[674]; 
    assign out[113] = ~layer_6[827]; 
    wire [1:0] far_7_7254_0;    relay_conn far_7_7254_0_a(.in(layer_6[1011]), .out(far_7_7254_0[0]));    relay_conn far_7_7254_0_b(.in(layer_6[902]), .out(far_7_7254_0[1]));
    wire [1:0] far_7_7254_1;    relay_conn far_7_7254_1_a(.in(far_7_7254_0[0]), .out(far_7_7254_1[0]));    relay_conn far_7_7254_1_b(.in(far_7_7254_0[1]), .out(far_7_7254_1[1]));
    wire [1:0] far_7_7254_2;    relay_conn far_7_7254_2_a(.in(far_7_7254_1[0]), .out(far_7_7254_2[0]));    relay_conn far_7_7254_2_b(.in(far_7_7254_1[1]), .out(far_7_7254_2[1]));
    assign out[114] = ~far_7_7254_2[1] | (far_7_7254_2[0] & far_7_7254_2[1]); 
    wire [1:0] far_7_7255_0;    relay_conn far_7_7255_0_a(.in(layer_6[210]), .out(far_7_7255_0[0]));    relay_conn far_7_7255_0_b(.in(layer_6[163]), .out(far_7_7255_0[1]));
    assign out[115] = ~(far_7_7255_0[0] | far_7_7255_0[1]); 
    assign out[116] = layer_6[659] & ~layer_6[663]; 
    wire [1:0] far_7_7257_0;    relay_conn far_7_7257_0_a(.in(layer_6[172]), .out(far_7_7257_0[0]));    relay_conn far_7_7257_0_b(.in(layer_6[100]), .out(far_7_7257_0[1]));
    wire [1:0] far_7_7257_1;    relay_conn far_7_7257_1_a(.in(far_7_7257_0[0]), .out(far_7_7257_1[0]));    relay_conn far_7_7257_1_b(.in(far_7_7257_0[1]), .out(far_7_7257_1[1]));
    assign out[117] = ~(far_7_7257_1[0] | far_7_7257_1[1]); 
    assign out[118] = layer_6[747]; 
    wire [1:0] far_7_7259_0;    relay_conn far_7_7259_0_a(.in(layer_6[272]), .out(far_7_7259_0[0]));    relay_conn far_7_7259_0_b(.in(layer_6[334]), .out(far_7_7259_0[1]));
    assign out[119] = far_7_7259_0[0] | far_7_7259_0[1]; 
    wire [1:0] far_7_7260_0;    relay_conn far_7_7260_0_a(.in(layer_6[811]), .out(far_7_7260_0[0]));    relay_conn far_7_7260_0_b(.in(layer_6[768]), .out(far_7_7260_0[1]));
    assign out[120] = far_7_7260_0[1]; 
    wire [1:0] far_7_7261_0;    relay_conn far_7_7261_0_a(.in(layer_6[541]), .out(far_7_7261_0[0]));    relay_conn far_7_7261_0_b(.in(layer_6[470]), .out(far_7_7261_0[1]));
    wire [1:0] far_7_7261_1;    relay_conn far_7_7261_1_a(.in(far_7_7261_0[0]), .out(far_7_7261_1[0]));    relay_conn far_7_7261_1_b(.in(far_7_7261_0[1]), .out(far_7_7261_1[1]));
    assign out[121] = far_7_7261_1[0] & far_7_7261_1[1]; 
    wire [1:0] far_7_7262_0;    relay_conn far_7_7262_0_a(.in(layer_6[9]), .out(far_7_7262_0[0]));    relay_conn far_7_7262_0_b(.in(layer_6[97]), .out(far_7_7262_0[1]));
    wire [1:0] far_7_7262_1;    relay_conn far_7_7262_1_a(.in(far_7_7262_0[0]), .out(far_7_7262_1[0]));    relay_conn far_7_7262_1_b(.in(far_7_7262_0[1]), .out(far_7_7262_1[1]));
    assign out[122] = ~(far_7_7262_1[0] ^ far_7_7262_1[1]); 
    wire [1:0] far_7_7263_0;    relay_conn far_7_7263_0_a(.in(layer_6[109]), .out(far_7_7263_0[0]));    relay_conn far_7_7263_0_b(.in(layer_6[225]), .out(far_7_7263_0[1]));
    wire [1:0] far_7_7263_1;    relay_conn far_7_7263_1_a(.in(far_7_7263_0[0]), .out(far_7_7263_1[0]));    relay_conn far_7_7263_1_b(.in(far_7_7263_0[1]), .out(far_7_7263_1[1]));
    wire [1:0] far_7_7263_2;    relay_conn far_7_7263_2_a(.in(far_7_7263_1[0]), .out(far_7_7263_2[0]));    relay_conn far_7_7263_2_b(.in(far_7_7263_1[1]), .out(far_7_7263_2[1]));
    assign out[123] = ~(far_7_7263_2[0] ^ far_7_7263_2[1]); 
    wire [1:0] far_7_7264_0;    relay_conn far_7_7264_0_a(.in(layer_6[157]), .out(far_7_7264_0[0]));    relay_conn far_7_7264_0_b(.in(layer_6[57]), .out(far_7_7264_0[1]));
    wire [1:0] far_7_7264_1;    relay_conn far_7_7264_1_a(.in(far_7_7264_0[0]), .out(far_7_7264_1[0]));    relay_conn far_7_7264_1_b(.in(far_7_7264_0[1]), .out(far_7_7264_1[1]));
    wire [1:0] far_7_7264_2;    relay_conn far_7_7264_2_a(.in(far_7_7264_1[0]), .out(far_7_7264_2[0]));    relay_conn far_7_7264_2_b(.in(far_7_7264_1[1]), .out(far_7_7264_2[1]));
    assign out[124] = far_7_7264_2[0] | far_7_7264_2[1]; 
    wire [1:0] far_7_7265_0;    relay_conn far_7_7265_0_a(.in(layer_6[881]), .out(far_7_7265_0[0]));    relay_conn far_7_7265_0_b(.in(layer_6[923]), .out(far_7_7265_0[1]));
    assign out[125] = far_7_7265_0[1]; 
    wire [1:0] far_7_7266_0;    relay_conn far_7_7266_0_a(.in(layer_6[623]), .out(far_7_7266_0[0]));    relay_conn far_7_7266_0_b(.in(layer_6[574]), .out(far_7_7266_0[1]));
    assign out[126] = ~far_7_7266_0[0]; 
    wire [1:0] far_7_7267_0;    relay_conn far_7_7267_0_a(.in(layer_6[388]), .out(far_7_7267_0[0]));    relay_conn far_7_7267_0_b(.in(layer_6[339]), .out(far_7_7267_0[1]));
    assign out[127] = far_7_7267_0[1]; 
    wire [1:0] far_7_7268_0;    relay_conn far_7_7268_0_a(.in(layer_6[475]), .out(far_7_7268_0[0]));    relay_conn far_7_7268_0_b(.in(layer_6[568]), .out(far_7_7268_0[1]));
    wire [1:0] far_7_7268_1;    relay_conn far_7_7268_1_a(.in(far_7_7268_0[0]), .out(far_7_7268_1[0]));    relay_conn far_7_7268_1_b(.in(far_7_7268_0[1]), .out(far_7_7268_1[1]));
    assign out[128] = ~(far_7_7268_1[0] | far_7_7268_1[1]); 
    wire [1:0] far_7_7269_0;    relay_conn far_7_7269_0_a(.in(layer_6[524]), .out(far_7_7269_0[0]));    relay_conn far_7_7269_0_b(.in(layer_6[415]), .out(far_7_7269_0[1]));
    wire [1:0] far_7_7269_1;    relay_conn far_7_7269_1_a(.in(far_7_7269_0[0]), .out(far_7_7269_1[0]));    relay_conn far_7_7269_1_b(.in(far_7_7269_0[1]), .out(far_7_7269_1[1]));
    wire [1:0] far_7_7269_2;    relay_conn far_7_7269_2_a(.in(far_7_7269_1[0]), .out(far_7_7269_2[0]));    relay_conn far_7_7269_2_b(.in(far_7_7269_1[1]), .out(far_7_7269_2[1]));
    assign out[129] = far_7_7269_2[1] & ~far_7_7269_2[0]; 
    wire [1:0] far_7_7270_0;    relay_conn far_7_7270_0_a(.in(layer_6[370]), .out(far_7_7270_0[0]));    relay_conn far_7_7270_0_b(.in(layer_6[455]), .out(far_7_7270_0[1]));
    wire [1:0] far_7_7270_1;    relay_conn far_7_7270_1_a(.in(far_7_7270_0[0]), .out(far_7_7270_1[0]));    relay_conn far_7_7270_1_b(.in(far_7_7270_0[1]), .out(far_7_7270_1[1]));
    assign out[130] = ~(far_7_7270_1[0] | far_7_7270_1[1]); 
    wire [1:0] far_7_7271_0;    relay_conn far_7_7271_0_a(.in(layer_6[272]), .out(far_7_7271_0[0]));    relay_conn far_7_7271_0_b(.in(layer_6[187]), .out(far_7_7271_0[1]));
    wire [1:0] far_7_7271_1;    relay_conn far_7_7271_1_a(.in(far_7_7271_0[0]), .out(far_7_7271_1[0]));    relay_conn far_7_7271_1_b(.in(far_7_7271_0[1]), .out(far_7_7271_1[1]));
    assign out[131] = far_7_7271_1[0] & ~far_7_7271_1[1]; 
    wire [1:0] far_7_7272_0;    relay_conn far_7_7272_0_a(.in(layer_6[553]), .out(far_7_7272_0[0]));    relay_conn far_7_7272_0_b(.in(layer_6[615]), .out(far_7_7272_0[1]));
    assign out[132] = ~far_7_7272_0[0]; 
    assign out[133] = ~(layer_6[718] ^ layer_6[711]); 
    wire [1:0] far_7_7274_0;    relay_conn far_7_7274_0_a(.in(layer_6[718]), .out(far_7_7274_0[0]));    relay_conn far_7_7274_0_b(.in(layer_6[829]), .out(far_7_7274_0[1]));
    wire [1:0] far_7_7274_1;    relay_conn far_7_7274_1_a(.in(far_7_7274_0[0]), .out(far_7_7274_1[0]));    relay_conn far_7_7274_1_b(.in(far_7_7274_0[1]), .out(far_7_7274_1[1]));
    wire [1:0] far_7_7274_2;    relay_conn far_7_7274_2_a(.in(far_7_7274_1[0]), .out(far_7_7274_2[0]));    relay_conn far_7_7274_2_b(.in(far_7_7274_1[1]), .out(far_7_7274_2[1]));
    assign out[134] = far_7_7274_2[0] ^ far_7_7274_2[1]; 
    wire [1:0] far_7_7275_0;    relay_conn far_7_7275_0_a(.in(layer_6[142]), .out(far_7_7275_0[0]));    relay_conn far_7_7275_0_b(.in(layer_6[203]), .out(far_7_7275_0[1]));
    assign out[135] = far_7_7275_0[0] & far_7_7275_0[1]; 
    assign out[136] = ~layer_6[315]; 
    assign out[137] = layer_6[159]; 
    wire [1:0] far_7_7278_0;    relay_conn far_7_7278_0_a(.in(layer_6[923]), .out(far_7_7278_0[0]));    relay_conn far_7_7278_0_b(.in(layer_6[1009]), .out(far_7_7278_0[1]));
    wire [1:0] far_7_7278_1;    relay_conn far_7_7278_1_a(.in(far_7_7278_0[0]), .out(far_7_7278_1[0]));    relay_conn far_7_7278_1_b(.in(far_7_7278_0[1]), .out(far_7_7278_1[1]));
    assign out[138] = ~far_7_7278_1[1] | (far_7_7278_1[0] & far_7_7278_1[1]); 
    assign out[139] = ~layer_6[136]; 
    assign out[140] = ~layer_6[163]; 
    wire [1:0] far_7_7281_0;    relay_conn far_7_7281_0_a(.in(layer_6[175]), .out(far_7_7281_0[0]));    relay_conn far_7_7281_0_b(.in(layer_6[261]), .out(far_7_7281_0[1]));
    wire [1:0] far_7_7281_1;    relay_conn far_7_7281_1_a(.in(far_7_7281_0[0]), .out(far_7_7281_1[0]));    relay_conn far_7_7281_1_b(.in(far_7_7281_0[1]), .out(far_7_7281_1[1]));
    assign out[141] = ~far_7_7281_1[1]; 
    assign out[142] = layer_6[406]; 
    wire [1:0] far_7_7283_0;    relay_conn far_7_7283_0_a(.in(layer_6[941]), .out(far_7_7283_0[0]));    relay_conn far_7_7283_0_b(.in(layer_6[1019]), .out(far_7_7283_0[1]));
    wire [1:0] far_7_7283_1;    relay_conn far_7_7283_1_a(.in(far_7_7283_0[0]), .out(far_7_7283_1[0]));    relay_conn far_7_7283_1_b(.in(far_7_7283_0[1]), .out(far_7_7283_1[1]));
    assign out[143] = far_7_7283_1[0]; 
    assign out[144] = ~layer_6[786] | (layer_6[786] & layer_6[814]); 
    assign out[145] = layer_6[407]; 
    assign out[146] = layer_6[601]; 
    assign out[147] = layer_6[157]; 
    wire [1:0] far_7_7288_0;    relay_conn far_7_7288_0_a(.in(layer_6[74]), .out(far_7_7288_0[0]));    relay_conn far_7_7288_0_b(.in(layer_6[24]), .out(far_7_7288_0[1]));
    assign out[148] = ~far_7_7288_0[1]; 
    wire [1:0] far_7_7289_0;    relay_conn far_7_7289_0_a(.in(layer_6[850]), .out(far_7_7289_0[0]));    relay_conn far_7_7289_0_b(.in(layer_6[789]), .out(far_7_7289_0[1]));
    assign out[149] = far_7_7289_0[0]; 
    wire [1:0] far_7_7290_0;    relay_conn far_7_7290_0_a(.in(layer_6[470]), .out(far_7_7290_0[0]));    relay_conn far_7_7290_0_b(.in(layer_6[571]), .out(far_7_7290_0[1]));
    wire [1:0] far_7_7290_1;    relay_conn far_7_7290_1_a(.in(far_7_7290_0[0]), .out(far_7_7290_1[0]));    relay_conn far_7_7290_1_b(.in(far_7_7290_0[1]), .out(far_7_7290_1[1]));
    wire [1:0] far_7_7290_2;    relay_conn far_7_7290_2_a(.in(far_7_7290_1[0]), .out(far_7_7290_2[0]));    relay_conn far_7_7290_2_b(.in(far_7_7290_1[1]), .out(far_7_7290_2[1]));
    assign out[150] = far_7_7290_2[1]; 
    wire [1:0] far_7_7291_0;    relay_conn far_7_7291_0_a(.in(layer_6[163]), .out(far_7_7291_0[0]));    relay_conn far_7_7291_0_b(.in(layer_6[56]), .out(far_7_7291_0[1]));
    wire [1:0] far_7_7291_1;    relay_conn far_7_7291_1_a(.in(far_7_7291_0[0]), .out(far_7_7291_1[0]));    relay_conn far_7_7291_1_b(.in(far_7_7291_0[1]), .out(far_7_7291_1[1]));
    wire [1:0] far_7_7291_2;    relay_conn far_7_7291_2_a(.in(far_7_7291_1[0]), .out(far_7_7291_2[0]));    relay_conn far_7_7291_2_b(.in(far_7_7291_1[1]), .out(far_7_7291_2[1]));
    assign out[151] = ~(far_7_7291_2[0] | far_7_7291_2[1]); 
    wire [1:0] far_7_7292_0;    relay_conn far_7_7292_0_a(.in(layer_6[543]), .out(far_7_7292_0[0]));    relay_conn far_7_7292_0_b(.in(layer_6[591]), .out(far_7_7292_0[1]));
    assign out[152] = far_7_7292_0[1] & ~far_7_7292_0[0]; 
    wire [1:0] far_7_7293_0;    relay_conn far_7_7293_0_a(.in(layer_6[449]), .out(far_7_7293_0[0]));    relay_conn far_7_7293_0_b(.in(layer_6[513]), .out(far_7_7293_0[1]));
    wire [1:0] far_7_7293_1;    relay_conn far_7_7293_1_a(.in(far_7_7293_0[0]), .out(far_7_7293_1[0]));    relay_conn far_7_7293_1_b(.in(far_7_7293_0[1]), .out(far_7_7293_1[1]));
    assign out[153] = ~far_7_7293_1[1]; 
    assign out[154] = layer_6[244] ^ layer_6[255]; 
    assign out[155] = ~(layer_6[676] & layer_6[699]); 
    wire [1:0] far_7_7296_0;    relay_conn far_7_7296_0_a(.in(layer_6[372]), .out(far_7_7296_0[0]));    relay_conn far_7_7296_0_b(.in(layer_6[435]), .out(far_7_7296_0[1]));
    assign out[156] = ~far_7_7296_0[0] | (far_7_7296_0[0] & far_7_7296_0[1]); 
    wire [1:0] far_7_7297_0;    relay_conn far_7_7297_0_a(.in(layer_6[489]), .out(far_7_7297_0[0]));    relay_conn far_7_7297_0_b(.in(layer_6[442]), .out(far_7_7297_0[1]));
    assign out[157] = ~far_7_7297_0[0]; 
    assign out[158] = layer_6[924] & ~layer_6[917]; 
    wire [1:0] far_7_7299_0;    relay_conn far_7_7299_0_a(.in(layer_6[71]), .out(far_7_7299_0[0]));    relay_conn far_7_7299_0_b(.in(layer_6[11]), .out(far_7_7299_0[1]));
    assign out[159] = ~far_7_7299_0[1]; 
    wire [1:0] far_7_7300_0;    relay_conn far_7_7300_0_a(.in(layer_6[621]), .out(far_7_7300_0[0]));    relay_conn far_7_7300_0_b(.in(layer_6[544]), .out(far_7_7300_0[1]));
    wire [1:0] far_7_7300_1;    relay_conn far_7_7300_1_a(.in(far_7_7300_0[0]), .out(far_7_7300_1[0]));    relay_conn far_7_7300_1_b(.in(far_7_7300_0[1]), .out(far_7_7300_1[1]));
    assign out[160] = far_7_7300_1[1]; 
    wire [1:0] far_7_7301_0;    relay_conn far_7_7301_0_a(.in(layer_6[923]), .out(far_7_7301_0[0]));    relay_conn far_7_7301_0_b(.in(layer_6[845]), .out(far_7_7301_0[1]));
    wire [1:0] far_7_7301_1;    relay_conn far_7_7301_1_a(.in(far_7_7301_0[0]), .out(far_7_7301_1[0]));    relay_conn far_7_7301_1_b(.in(far_7_7301_0[1]), .out(far_7_7301_1[1]));
    assign out[161] = far_7_7301_1[0] & far_7_7301_1[1]; 
    wire [1:0] far_7_7302_0;    relay_conn far_7_7302_0_a(.in(layer_6[659]), .out(far_7_7302_0[0]));    relay_conn far_7_7302_0_b(.in(layer_6[737]), .out(far_7_7302_0[1]));
    wire [1:0] far_7_7302_1;    relay_conn far_7_7302_1_a(.in(far_7_7302_0[0]), .out(far_7_7302_1[0]));    relay_conn far_7_7302_1_b(.in(far_7_7302_0[1]), .out(far_7_7302_1[1]));
    assign out[162] = ~far_7_7302_1[1] | (far_7_7302_1[0] & far_7_7302_1[1]); 
    assign out[163] = ~(layer_6[374] | layer_6[370]); 
    wire [1:0] far_7_7304_0;    relay_conn far_7_7304_0_a(.in(layer_6[777]), .out(far_7_7304_0[0]));    relay_conn far_7_7304_0_b(.in(layer_6[896]), .out(far_7_7304_0[1]));
    wire [1:0] far_7_7304_1;    relay_conn far_7_7304_1_a(.in(far_7_7304_0[0]), .out(far_7_7304_1[0]));    relay_conn far_7_7304_1_b(.in(far_7_7304_0[1]), .out(far_7_7304_1[1]));
    wire [1:0] far_7_7304_2;    relay_conn far_7_7304_2_a(.in(far_7_7304_1[0]), .out(far_7_7304_2[0]));    relay_conn far_7_7304_2_b(.in(far_7_7304_1[1]), .out(far_7_7304_2[1]));
    assign out[164] = far_7_7304_2[0] | far_7_7304_2[1]; 
    wire [1:0] far_7_7305_0;    relay_conn far_7_7305_0_a(.in(layer_6[465]), .out(far_7_7305_0[0]));    relay_conn far_7_7305_0_b(.in(layer_6[345]), .out(far_7_7305_0[1]));
    wire [1:0] far_7_7305_1;    relay_conn far_7_7305_1_a(.in(far_7_7305_0[0]), .out(far_7_7305_1[0]));    relay_conn far_7_7305_1_b(.in(far_7_7305_0[1]), .out(far_7_7305_1[1]));
    wire [1:0] far_7_7305_2;    relay_conn far_7_7305_2_a(.in(far_7_7305_1[0]), .out(far_7_7305_2[0]));    relay_conn far_7_7305_2_b(.in(far_7_7305_1[1]), .out(far_7_7305_2[1]));
    assign out[165] = far_7_7305_2[0] & ~far_7_7305_2[1]; 
    wire [1:0] far_7_7306_0;    relay_conn far_7_7306_0_a(.in(layer_6[139]), .out(far_7_7306_0[0]));    relay_conn far_7_7306_0_b(.in(layer_6[267]), .out(far_7_7306_0[1]));
    wire [1:0] far_7_7306_1;    relay_conn far_7_7306_1_a(.in(far_7_7306_0[0]), .out(far_7_7306_1[0]));    relay_conn far_7_7306_1_b(.in(far_7_7306_0[1]), .out(far_7_7306_1[1]));
    wire [1:0] far_7_7306_2;    relay_conn far_7_7306_2_a(.in(far_7_7306_1[0]), .out(far_7_7306_2[0]));    relay_conn far_7_7306_2_b(.in(far_7_7306_1[1]), .out(far_7_7306_2[1]));
    wire [1:0] far_7_7306_3;    relay_conn far_7_7306_3_a(.in(far_7_7306_2[0]), .out(far_7_7306_3[0]));    relay_conn far_7_7306_3_b(.in(far_7_7306_2[1]), .out(far_7_7306_3[1]));
    assign out[166] = far_7_7306_3[0]; 
    wire [1:0] far_7_7307_0;    relay_conn far_7_7307_0_a(.in(layer_6[46]), .out(far_7_7307_0[0]));    relay_conn far_7_7307_0_b(.in(layer_6[110]), .out(far_7_7307_0[1]));
    wire [1:0] far_7_7307_1;    relay_conn far_7_7307_1_a(.in(far_7_7307_0[0]), .out(far_7_7307_1[0]));    relay_conn far_7_7307_1_b(.in(far_7_7307_0[1]), .out(far_7_7307_1[1]));
    assign out[167] = far_7_7307_1[1]; 
    assign out[168] = ~layer_6[158] | (layer_6[158] & layer_6[157]); 
    wire [1:0] far_7_7309_0;    relay_conn far_7_7309_0_a(.in(layer_6[103]), .out(far_7_7309_0[0]));    relay_conn far_7_7309_0_b(.in(layer_6[149]), .out(far_7_7309_0[1]));
    assign out[169] = ~far_7_7309_0[0]; 
    wire [1:0] far_7_7310_0;    relay_conn far_7_7310_0_a(.in(layer_6[732]), .out(far_7_7310_0[0]));    relay_conn far_7_7310_0_b(.in(layer_6[644]), .out(far_7_7310_0[1]));
    wire [1:0] far_7_7310_1;    relay_conn far_7_7310_1_a(.in(far_7_7310_0[0]), .out(far_7_7310_1[0]));    relay_conn far_7_7310_1_b(.in(far_7_7310_0[1]), .out(far_7_7310_1[1]));
    assign out[170] = ~(far_7_7310_1[0] | far_7_7310_1[1]); 
    wire [1:0] far_7_7311_0;    relay_conn far_7_7311_0_a(.in(layer_6[816]), .out(far_7_7311_0[0]));    relay_conn far_7_7311_0_b(.in(layer_6[765]), .out(far_7_7311_0[1]));
    assign out[171] = far_7_7311_0[0]; 
    wire [1:0] far_7_7312_0;    relay_conn far_7_7312_0_a(.in(layer_6[896]), .out(far_7_7312_0[0]));    relay_conn far_7_7312_0_b(.in(layer_6[932]), .out(far_7_7312_0[1]));
    assign out[172] = ~far_7_7312_0[1] | (far_7_7312_0[0] & far_7_7312_0[1]); 
    wire [1:0] far_7_7313_0;    relay_conn far_7_7313_0_a(.in(layer_6[930]), .out(far_7_7313_0[0]));    relay_conn far_7_7313_0_b(.in(layer_6[967]), .out(far_7_7313_0[1]));
    assign out[173] = ~far_7_7313_0[0]; 
    wire [1:0] far_7_7314_0;    relay_conn far_7_7314_0_a(.in(layer_6[671]), .out(far_7_7314_0[0]));    relay_conn far_7_7314_0_b(.in(layer_6[708]), .out(far_7_7314_0[1]));
    assign out[174] = ~far_7_7314_0[1]; 
    wire [1:0] far_7_7315_0;    relay_conn far_7_7315_0_a(.in(layer_6[209]), .out(far_7_7315_0[0]));    relay_conn far_7_7315_0_b(.in(layer_6[336]), .out(far_7_7315_0[1]));
    wire [1:0] far_7_7315_1;    relay_conn far_7_7315_1_a(.in(far_7_7315_0[0]), .out(far_7_7315_1[0]));    relay_conn far_7_7315_1_b(.in(far_7_7315_0[1]), .out(far_7_7315_1[1]));
    wire [1:0] far_7_7315_2;    relay_conn far_7_7315_2_a(.in(far_7_7315_1[0]), .out(far_7_7315_2[0]));    relay_conn far_7_7315_2_b(.in(far_7_7315_1[1]), .out(far_7_7315_2[1]));
    assign out[175] = ~(far_7_7315_2[0] | far_7_7315_2[1]); 
    wire [1:0] far_7_7316_0;    relay_conn far_7_7316_0_a(.in(layer_6[273]), .out(far_7_7316_0[0]));    relay_conn far_7_7316_0_b(.in(layer_6[328]), .out(far_7_7316_0[1]));
    assign out[176] = far_7_7316_0[1]; 
    wire [1:0] far_7_7317_0;    relay_conn far_7_7317_0_a(.in(layer_6[535]), .out(far_7_7317_0[0]));    relay_conn far_7_7317_0_b(.in(layer_6[569]), .out(far_7_7317_0[1]));
    assign out[177] = ~(far_7_7317_0[0] & far_7_7317_0[1]); 
    wire [1:0] far_7_7318_0;    relay_conn far_7_7318_0_a(.in(layer_6[706]), .out(far_7_7318_0[0]));    relay_conn far_7_7318_0_b(.in(layer_6[629]), .out(far_7_7318_0[1]));
    wire [1:0] far_7_7318_1;    relay_conn far_7_7318_1_a(.in(far_7_7318_0[0]), .out(far_7_7318_1[0]));    relay_conn far_7_7318_1_b(.in(far_7_7318_0[1]), .out(far_7_7318_1[1]));
    assign out[178] = far_7_7318_1[1]; 
    wire [1:0] far_7_7319_0;    relay_conn far_7_7319_0_a(.in(layer_6[780]), .out(far_7_7319_0[0]));    relay_conn far_7_7319_0_b(.in(layer_6[849]), .out(far_7_7319_0[1]));
    wire [1:0] far_7_7319_1;    relay_conn far_7_7319_1_a(.in(far_7_7319_0[0]), .out(far_7_7319_1[0]));    relay_conn far_7_7319_1_b(.in(far_7_7319_0[1]), .out(far_7_7319_1[1]));
    assign out[179] = far_7_7319_1[0]; 
    wire [1:0] far_7_7320_0;    relay_conn far_7_7320_0_a(.in(layer_6[597]), .out(far_7_7320_0[0]));    relay_conn far_7_7320_0_b(.in(layer_6[499]), .out(far_7_7320_0[1]));
    wire [1:0] far_7_7320_1;    relay_conn far_7_7320_1_a(.in(far_7_7320_0[0]), .out(far_7_7320_1[0]));    relay_conn far_7_7320_1_b(.in(far_7_7320_0[1]), .out(far_7_7320_1[1]));
    wire [1:0] far_7_7320_2;    relay_conn far_7_7320_2_a(.in(far_7_7320_1[0]), .out(far_7_7320_2[0]));    relay_conn far_7_7320_2_b(.in(far_7_7320_1[1]), .out(far_7_7320_2[1]));
    assign out[180] = far_7_7320_2[0] ^ far_7_7320_2[1]; 
    wire [1:0] far_7_7321_0;    relay_conn far_7_7321_0_a(.in(layer_6[1011]), .out(far_7_7321_0[0]));    relay_conn far_7_7321_0_b(.in(layer_6[884]), .out(far_7_7321_0[1]));
    wire [1:0] far_7_7321_1;    relay_conn far_7_7321_1_a(.in(far_7_7321_0[0]), .out(far_7_7321_1[0]));    relay_conn far_7_7321_1_b(.in(far_7_7321_0[1]), .out(far_7_7321_1[1]));
    wire [1:0] far_7_7321_2;    relay_conn far_7_7321_2_a(.in(far_7_7321_1[0]), .out(far_7_7321_2[0]));    relay_conn far_7_7321_2_b(.in(far_7_7321_1[1]), .out(far_7_7321_2[1]));
    assign out[181] = far_7_7321_2[0]; 
    assign out[182] = ~layer_6[966]; 
    wire [1:0] far_7_7323_0;    relay_conn far_7_7323_0_a(.in(layer_6[913]), .out(far_7_7323_0[0]));    relay_conn far_7_7323_0_b(.in(layer_6[839]), .out(far_7_7323_0[1]));
    wire [1:0] far_7_7323_1;    relay_conn far_7_7323_1_a(.in(far_7_7323_0[0]), .out(far_7_7323_1[0]));    relay_conn far_7_7323_1_b(.in(far_7_7323_0[1]), .out(far_7_7323_1[1]));
    assign out[183] = far_7_7323_1[0]; 
    assign out[184] = layer_6[174] & layer_6[194]; 
    wire [1:0] far_7_7325_0;    relay_conn far_7_7325_0_a(.in(layer_6[764]), .out(far_7_7325_0[0]));    relay_conn far_7_7325_0_b(.in(layer_6[672]), .out(far_7_7325_0[1]));
    wire [1:0] far_7_7325_1;    relay_conn far_7_7325_1_a(.in(far_7_7325_0[0]), .out(far_7_7325_1[0]));    relay_conn far_7_7325_1_b(.in(far_7_7325_0[1]), .out(far_7_7325_1[1]));
    assign out[185] = ~(far_7_7325_1[0] | far_7_7325_1[1]); 
    wire [1:0] far_7_7326_0;    relay_conn far_7_7326_0_a(.in(layer_6[604]), .out(far_7_7326_0[0]));    relay_conn far_7_7326_0_b(.in(layer_6[485]), .out(far_7_7326_0[1]));
    wire [1:0] far_7_7326_1;    relay_conn far_7_7326_1_a(.in(far_7_7326_0[0]), .out(far_7_7326_1[0]));    relay_conn far_7_7326_1_b(.in(far_7_7326_0[1]), .out(far_7_7326_1[1]));
    wire [1:0] far_7_7326_2;    relay_conn far_7_7326_2_a(.in(far_7_7326_1[0]), .out(far_7_7326_2[0]));    relay_conn far_7_7326_2_b(.in(far_7_7326_1[1]), .out(far_7_7326_2[1]));
    assign out[186] = ~(far_7_7326_2[0] ^ far_7_7326_2[1]); 
    assign out[187] = layer_6[249]; 
    wire [1:0] far_7_7328_0;    relay_conn far_7_7328_0_a(.in(layer_6[265]), .out(far_7_7328_0[0]));    relay_conn far_7_7328_0_b(.in(layer_6[199]), .out(far_7_7328_0[1]));
    wire [1:0] far_7_7328_1;    relay_conn far_7_7328_1_a(.in(far_7_7328_0[0]), .out(far_7_7328_1[0]));    relay_conn far_7_7328_1_b(.in(far_7_7328_0[1]), .out(far_7_7328_1[1]));
    assign out[188] = far_7_7328_1[0] | far_7_7328_1[1]; 
    wire [1:0] far_7_7329_0;    relay_conn far_7_7329_0_a(.in(layer_6[416]), .out(far_7_7329_0[0]));    relay_conn far_7_7329_0_b(.in(layer_6[456]), .out(far_7_7329_0[1]));
    assign out[189] = ~far_7_7329_0[1] | (far_7_7329_0[0] & far_7_7329_0[1]); 
    wire [1:0] far_7_7330_0;    relay_conn far_7_7330_0_a(.in(layer_6[911]), .out(far_7_7330_0[0]));    relay_conn far_7_7330_0_b(.in(layer_6[803]), .out(far_7_7330_0[1]));
    wire [1:0] far_7_7330_1;    relay_conn far_7_7330_1_a(.in(far_7_7330_0[0]), .out(far_7_7330_1[0]));    relay_conn far_7_7330_1_b(.in(far_7_7330_0[1]), .out(far_7_7330_1[1]));
    wire [1:0] far_7_7330_2;    relay_conn far_7_7330_2_a(.in(far_7_7330_1[0]), .out(far_7_7330_2[0]));    relay_conn far_7_7330_2_b(.in(far_7_7330_1[1]), .out(far_7_7330_2[1]));
    assign out[190] = ~far_7_7330_2[0]; 
    wire [1:0] far_7_7331_0;    relay_conn far_7_7331_0_a(.in(layer_6[924]), .out(far_7_7331_0[0]));    relay_conn far_7_7331_0_b(.in(layer_6[959]), .out(far_7_7331_0[1]));
    assign out[191] = far_7_7331_0[0] | far_7_7331_0[1]; 
    wire [1:0] far_7_7332_0;    relay_conn far_7_7332_0_a(.in(layer_6[515]), .out(far_7_7332_0[0]));    relay_conn far_7_7332_0_b(.in(layer_6[404]), .out(far_7_7332_0[1]));
    wire [1:0] far_7_7332_1;    relay_conn far_7_7332_1_a(.in(far_7_7332_0[0]), .out(far_7_7332_1[0]));    relay_conn far_7_7332_1_b(.in(far_7_7332_0[1]), .out(far_7_7332_1[1]));
    wire [1:0] far_7_7332_2;    relay_conn far_7_7332_2_a(.in(far_7_7332_1[0]), .out(far_7_7332_2[0]));    relay_conn far_7_7332_2_b(.in(far_7_7332_1[1]), .out(far_7_7332_2[1]));
    assign out[192] = far_7_7332_2[0] & far_7_7332_2[1]; 
    assign out[193] = layer_6[539] & ~layer_6[516]; 
    assign out[194] = layer_6[317]; 
    wire [1:0] far_7_7335_0;    relay_conn far_7_7335_0_a(.in(layer_6[944]), .out(far_7_7335_0[0]));    relay_conn far_7_7335_0_b(.in(layer_6[1008]), .out(far_7_7335_0[1]));
    wire [1:0] far_7_7335_1;    relay_conn far_7_7335_1_a(.in(far_7_7335_0[0]), .out(far_7_7335_1[0]));    relay_conn far_7_7335_1_b(.in(far_7_7335_0[1]), .out(far_7_7335_1[1]));
    assign out[195] = far_7_7335_1[0] ^ far_7_7335_1[1]; 
    wire [1:0] far_7_7336_0;    relay_conn far_7_7336_0_a(.in(layer_6[681]), .out(far_7_7336_0[0]));    relay_conn far_7_7336_0_b(.in(layer_6[729]), .out(far_7_7336_0[1]));
    assign out[196] = ~far_7_7336_0[1]; 
    wire [1:0] far_7_7337_0;    relay_conn far_7_7337_0_a(.in(layer_6[329]), .out(far_7_7337_0[0]));    relay_conn far_7_7337_0_b(.in(layer_6[256]), .out(far_7_7337_0[1]));
    wire [1:0] far_7_7337_1;    relay_conn far_7_7337_1_a(.in(far_7_7337_0[0]), .out(far_7_7337_1[0]));    relay_conn far_7_7337_1_b(.in(far_7_7337_0[1]), .out(far_7_7337_1[1]));
    assign out[197] = ~far_7_7337_1[1]; 
    wire [1:0] far_7_7338_0;    relay_conn far_7_7338_0_a(.in(layer_6[79]), .out(far_7_7338_0[0]));    relay_conn far_7_7338_0_b(.in(layer_6[25]), .out(far_7_7338_0[1]));
    assign out[198] = far_7_7338_0[0] & ~far_7_7338_0[1]; 
    wire [1:0] far_7_7339_0;    relay_conn far_7_7339_0_a(.in(layer_6[253]), .out(far_7_7339_0[0]));    relay_conn far_7_7339_0_b(.in(layer_6[331]), .out(far_7_7339_0[1]));
    wire [1:0] far_7_7339_1;    relay_conn far_7_7339_1_a(.in(far_7_7339_0[0]), .out(far_7_7339_1[0]));    relay_conn far_7_7339_1_b(.in(far_7_7339_0[1]), .out(far_7_7339_1[1]));
    assign out[199] = ~(far_7_7339_1[0] & far_7_7339_1[1]); 
    wire [1:0] far_7_7340_0;    relay_conn far_7_7340_0_a(.in(layer_6[45]), .out(far_7_7340_0[0]));    relay_conn far_7_7340_0_b(.in(layer_6[153]), .out(far_7_7340_0[1]));
    wire [1:0] far_7_7340_1;    relay_conn far_7_7340_1_a(.in(far_7_7340_0[0]), .out(far_7_7340_1[0]));    relay_conn far_7_7340_1_b(.in(far_7_7340_0[1]), .out(far_7_7340_1[1]));
    wire [1:0] far_7_7340_2;    relay_conn far_7_7340_2_a(.in(far_7_7340_1[0]), .out(far_7_7340_2[0]));    relay_conn far_7_7340_2_b(.in(far_7_7340_1[1]), .out(far_7_7340_2[1]));
    assign out[200] = ~far_7_7340_2[1]; 
    wire [1:0] far_7_7341_0;    relay_conn far_7_7341_0_a(.in(layer_6[737]), .out(far_7_7341_0[0]));    relay_conn far_7_7341_0_b(.in(layer_6[693]), .out(far_7_7341_0[1]));
    assign out[201] = ~(far_7_7341_0[0] ^ far_7_7341_0[1]); 
    wire [1:0] far_7_7342_0;    relay_conn far_7_7342_0_a(.in(layer_6[515]), .out(far_7_7342_0[0]));    relay_conn far_7_7342_0_b(.in(layer_6[476]), .out(far_7_7342_0[1]));
    assign out[202] = far_7_7342_0[0]; 
    wire [1:0] far_7_7343_0;    relay_conn far_7_7343_0_a(.in(layer_6[484]), .out(far_7_7343_0[0]));    relay_conn far_7_7343_0_b(.in(layer_6[526]), .out(far_7_7343_0[1]));
    assign out[203] = ~far_7_7343_0[1] | (far_7_7343_0[0] & far_7_7343_0[1]); 
    assign out[204] = layer_6[195] & ~layer_6[222]; 
    assign out[205] = layer_6[552] & ~layer_6[536]; 
    wire [1:0] far_7_7346_0;    relay_conn far_7_7346_0_a(.in(layer_6[194]), .out(far_7_7346_0[0]));    relay_conn far_7_7346_0_b(.in(layer_6[315]), .out(far_7_7346_0[1]));
    wire [1:0] far_7_7346_1;    relay_conn far_7_7346_1_a(.in(far_7_7346_0[0]), .out(far_7_7346_1[0]));    relay_conn far_7_7346_1_b(.in(far_7_7346_0[1]), .out(far_7_7346_1[1]));
    wire [1:0] far_7_7346_2;    relay_conn far_7_7346_2_a(.in(far_7_7346_1[0]), .out(far_7_7346_2[0]));    relay_conn far_7_7346_2_b(.in(far_7_7346_1[1]), .out(far_7_7346_2[1]));
    assign out[206] = ~(far_7_7346_2[0] ^ far_7_7346_2[1]); 
    assign out[207] = layer_6[703]; 
    wire [1:0] far_7_7348_0;    relay_conn far_7_7348_0_a(.in(layer_6[329]), .out(far_7_7348_0[0]));    relay_conn far_7_7348_0_b(.in(layer_6[249]), .out(far_7_7348_0[1]));
    wire [1:0] far_7_7348_1;    relay_conn far_7_7348_1_a(.in(far_7_7348_0[0]), .out(far_7_7348_1[0]));    relay_conn far_7_7348_1_b(.in(far_7_7348_0[1]), .out(far_7_7348_1[1]));
    assign out[208] = ~(far_7_7348_1[0] & far_7_7348_1[1]); 
    wire [1:0] far_7_7349_0;    relay_conn far_7_7349_0_a(.in(layer_6[504]), .out(far_7_7349_0[0]));    relay_conn far_7_7349_0_b(.in(layer_6[624]), .out(far_7_7349_0[1]));
    wire [1:0] far_7_7349_1;    relay_conn far_7_7349_1_a(.in(far_7_7349_0[0]), .out(far_7_7349_1[0]));    relay_conn far_7_7349_1_b(.in(far_7_7349_0[1]), .out(far_7_7349_1[1]));
    wire [1:0] far_7_7349_2;    relay_conn far_7_7349_2_a(.in(far_7_7349_1[0]), .out(far_7_7349_2[0]));    relay_conn far_7_7349_2_b(.in(far_7_7349_1[1]), .out(far_7_7349_2[1]));
    assign out[209] = ~(far_7_7349_2[0] | far_7_7349_2[1]); 
    wire [1:0] far_7_7350_0;    relay_conn far_7_7350_0_a(.in(layer_6[567]), .out(far_7_7350_0[0]));    relay_conn far_7_7350_0_b(.in(layer_6[682]), .out(far_7_7350_0[1]));
    wire [1:0] far_7_7350_1;    relay_conn far_7_7350_1_a(.in(far_7_7350_0[0]), .out(far_7_7350_1[0]));    relay_conn far_7_7350_1_b(.in(far_7_7350_0[1]), .out(far_7_7350_1[1]));
    wire [1:0] far_7_7350_2;    relay_conn far_7_7350_2_a(.in(far_7_7350_1[0]), .out(far_7_7350_2[0]));    relay_conn far_7_7350_2_b(.in(far_7_7350_1[1]), .out(far_7_7350_2[1]));
    assign out[210] = ~far_7_7350_2[0]; 
    wire [1:0] far_7_7351_0;    relay_conn far_7_7351_0_a(.in(layer_6[407]), .out(far_7_7351_0[0]));    relay_conn far_7_7351_0_b(.in(layer_6[289]), .out(far_7_7351_0[1]));
    wire [1:0] far_7_7351_1;    relay_conn far_7_7351_1_a(.in(far_7_7351_0[0]), .out(far_7_7351_1[0]));    relay_conn far_7_7351_1_b(.in(far_7_7351_0[1]), .out(far_7_7351_1[1]));
    wire [1:0] far_7_7351_2;    relay_conn far_7_7351_2_a(.in(far_7_7351_1[0]), .out(far_7_7351_2[0]));    relay_conn far_7_7351_2_b(.in(far_7_7351_1[1]), .out(far_7_7351_2[1]));
    assign out[211] = ~(far_7_7351_2[0] & far_7_7351_2[1]); 
    wire [1:0] far_7_7352_0;    relay_conn far_7_7352_0_a(.in(layer_6[515]), .out(far_7_7352_0[0]));    relay_conn far_7_7352_0_b(.in(layer_6[548]), .out(far_7_7352_0[1]));
    assign out[212] = ~far_7_7352_0[0]; 
    wire [1:0] far_7_7353_0;    relay_conn far_7_7353_0_a(.in(layer_6[122]), .out(far_7_7353_0[0]));    relay_conn far_7_7353_0_b(.in(layer_6[7]), .out(far_7_7353_0[1]));
    wire [1:0] far_7_7353_1;    relay_conn far_7_7353_1_a(.in(far_7_7353_0[0]), .out(far_7_7353_1[0]));    relay_conn far_7_7353_1_b(.in(far_7_7353_0[1]), .out(far_7_7353_1[1]));
    wire [1:0] far_7_7353_2;    relay_conn far_7_7353_2_a(.in(far_7_7353_1[0]), .out(far_7_7353_2[0]));    relay_conn far_7_7353_2_b(.in(far_7_7353_1[1]), .out(far_7_7353_2[1]));
    assign out[213] = ~far_7_7353_2[0] | (far_7_7353_2[0] & far_7_7353_2[1]); 
    wire [1:0] far_7_7354_0;    relay_conn far_7_7354_0_a(.in(layer_6[829]), .out(far_7_7354_0[0]));    relay_conn far_7_7354_0_b(.in(layer_6[923]), .out(far_7_7354_0[1]));
    wire [1:0] far_7_7354_1;    relay_conn far_7_7354_1_a(.in(far_7_7354_0[0]), .out(far_7_7354_1[0]));    relay_conn far_7_7354_1_b(.in(far_7_7354_0[1]), .out(far_7_7354_1[1]));
    assign out[214] = far_7_7354_1[1]; 
    assign out[215] = ~layer_6[971] | (layer_6[971] & layer_6[941]); 
    assign out[216] = ~(layer_6[387] & layer_6[369]); 
    wire [1:0] far_7_7357_0;    relay_conn far_7_7357_0_a(.in(layer_6[419]), .out(far_7_7357_0[0]));    relay_conn far_7_7357_0_b(.in(layer_6[337]), .out(far_7_7357_0[1]));
    wire [1:0] far_7_7357_1;    relay_conn far_7_7357_1_a(.in(far_7_7357_0[0]), .out(far_7_7357_1[0]));    relay_conn far_7_7357_1_b(.in(far_7_7357_0[1]), .out(far_7_7357_1[1]));
    assign out[217] = far_7_7357_1[0]; 
    wire [1:0] far_7_7358_0;    relay_conn far_7_7358_0_a(.in(layer_6[320]), .out(far_7_7358_0[0]));    relay_conn far_7_7358_0_b(.in(layer_6[198]), .out(far_7_7358_0[1]));
    wire [1:0] far_7_7358_1;    relay_conn far_7_7358_1_a(.in(far_7_7358_0[0]), .out(far_7_7358_1[0]));    relay_conn far_7_7358_1_b(.in(far_7_7358_0[1]), .out(far_7_7358_1[1]));
    wire [1:0] far_7_7358_2;    relay_conn far_7_7358_2_a(.in(far_7_7358_1[0]), .out(far_7_7358_2[0]));    relay_conn far_7_7358_2_b(.in(far_7_7358_1[1]), .out(far_7_7358_2[1]));
    assign out[218] = far_7_7358_2[1] & ~far_7_7358_2[0]; 
    assign out[219] = layer_6[485] & ~layer_6[466]; 
    wire [1:0] far_7_7360_0;    relay_conn far_7_7360_0_a(.in(layer_6[40]), .out(far_7_7360_0[0]));    relay_conn far_7_7360_0_b(.in(layer_6[136]), .out(far_7_7360_0[1]));
    wire [1:0] far_7_7360_1;    relay_conn far_7_7360_1_a(.in(far_7_7360_0[0]), .out(far_7_7360_1[0]));    relay_conn far_7_7360_1_b(.in(far_7_7360_0[1]), .out(far_7_7360_1[1]));
    wire [1:0] far_7_7360_2;    relay_conn far_7_7360_2_a(.in(far_7_7360_1[0]), .out(far_7_7360_2[0]));    relay_conn far_7_7360_2_b(.in(far_7_7360_1[1]), .out(far_7_7360_2[1]));
    assign out[220] = ~far_7_7360_2[1]; 
    wire [1:0] far_7_7361_0;    relay_conn far_7_7361_0_a(.in(layer_6[497]), .out(far_7_7361_0[0]));    relay_conn far_7_7361_0_b(.in(layer_6[417]), .out(far_7_7361_0[1]));
    wire [1:0] far_7_7361_1;    relay_conn far_7_7361_1_a(.in(far_7_7361_0[0]), .out(far_7_7361_1[0]));    relay_conn far_7_7361_1_b(.in(far_7_7361_0[1]), .out(far_7_7361_1[1]));
    assign out[221] = far_7_7361_1[0] & far_7_7361_1[1]; 
    wire [1:0] far_7_7362_0;    relay_conn far_7_7362_0_a(.in(layer_6[608]), .out(far_7_7362_0[0]));    relay_conn far_7_7362_0_b(.in(layer_6[698]), .out(far_7_7362_0[1]));
    wire [1:0] far_7_7362_1;    relay_conn far_7_7362_1_a(.in(far_7_7362_0[0]), .out(far_7_7362_1[0]));    relay_conn far_7_7362_1_b(.in(far_7_7362_0[1]), .out(far_7_7362_1[1]));
    assign out[222] = far_7_7362_1[1]; 
    wire [1:0] far_7_7363_0;    relay_conn far_7_7363_0_a(.in(layer_6[207]), .out(far_7_7363_0[0]));    relay_conn far_7_7363_0_b(.in(layer_6[141]), .out(far_7_7363_0[1]));
    wire [1:0] far_7_7363_1;    relay_conn far_7_7363_1_a(.in(far_7_7363_0[0]), .out(far_7_7363_1[0]));    relay_conn far_7_7363_1_b(.in(far_7_7363_0[1]), .out(far_7_7363_1[1]));
    assign out[223] = far_7_7363_1[0] ^ far_7_7363_1[1]; 
    wire [1:0] far_7_7364_0;    relay_conn far_7_7364_0_a(.in(layer_6[705]), .out(far_7_7364_0[0]));    relay_conn far_7_7364_0_b(.in(layer_6[758]), .out(far_7_7364_0[1]));
    assign out[224] = ~far_7_7364_0[0]; 
    assign out[225] = ~(layer_6[718] ^ layer_6[737]); 
    wire [1:0] far_7_7366_0;    relay_conn far_7_7366_0_a(.in(layer_6[157]), .out(far_7_7366_0[0]));    relay_conn far_7_7366_0_b(.in(layer_6[57]), .out(far_7_7366_0[1]));
    wire [1:0] far_7_7366_1;    relay_conn far_7_7366_1_a(.in(far_7_7366_0[0]), .out(far_7_7366_1[0]));    relay_conn far_7_7366_1_b(.in(far_7_7366_0[1]), .out(far_7_7366_1[1]));
    wire [1:0] far_7_7366_2;    relay_conn far_7_7366_2_a(.in(far_7_7366_1[0]), .out(far_7_7366_2[0]));    relay_conn far_7_7366_2_b(.in(far_7_7366_1[1]), .out(far_7_7366_2[1]));
    assign out[226] = far_7_7366_2[1]; 
    wire [1:0] far_7_7367_0;    relay_conn far_7_7367_0_a(.in(layer_6[394]), .out(far_7_7367_0[0]));    relay_conn far_7_7367_0_b(.in(layer_6[513]), .out(far_7_7367_0[1]));
    wire [1:0] far_7_7367_1;    relay_conn far_7_7367_1_a(.in(far_7_7367_0[0]), .out(far_7_7367_1[0]));    relay_conn far_7_7367_1_b(.in(far_7_7367_0[1]), .out(far_7_7367_1[1]));
    wire [1:0] far_7_7367_2;    relay_conn far_7_7367_2_a(.in(far_7_7367_1[0]), .out(far_7_7367_2[0]));    relay_conn far_7_7367_2_b(.in(far_7_7367_1[1]), .out(far_7_7367_2[1]));
    assign out[227] = far_7_7367_2[0]; 
    wire [1:0] far_7_7368_0;    relay_conn far_7_7368_0_a(.in(layer_6[557]), .out(far_7_7368_0[0]));    relay_conn far_7_7368_0_b(.in(layer_6[615]), .out(far_7_7368_0[1]));
    assign out[228] = far_7_7368_0[0] & far_7_7368_0[1]; 
    assign out[229] = layer_6[190]; 
    wire [1:0] far_7_7370_0;    relay_conn far_7_7370_0_a(.in(layer_6[333]), .out(far_7_7370_0[0]));    relay_conn far_7_7370_0_b(.in(layer_6[214]), .out(far_7_7370_0[1]));
    wire [1:0] far_7_7370_1;    relay_conn far_7_7370_1_a(.in(far_7_7370_0[0]), .out(far_7_7370_1[0]));    relay_conn far_7_7370_1_b(.in(far_7_7370_0[1]), .out(far_7_7370_1[1]));
    wire [1:0] far_7_7370_2;    relay_conn far_7_7370_2_a(.in(far_7_7370_1[0]), .out(far_7_7370_2[0]));    relay_conn far_7_7370_2_b(.in(far_7_7370_1[1]), .out(far_7_7370_2[1]));
    assign out[230] = ~far_7_7370_2[1]; 
    assign out[231] = ~(layer_6[129] | layer_6[116]); 
    wire [1:0] far_7_7372_0;    relay_conn far_7_7372_0_a(.in(layer_6[635]), .out(far_7_7372_0[0]));    relay_conn far_7_7372_0_b(.in(layer_6[601]), .out(far_7_7372_0[1]));
    assign out[232] = ~far_7_7372_0[1]; 
    wire [1:0] far_7_7373_0;    relay_conn far_7_7373_0_a(.in(layer_6[1]), .out(far_7_7373_0[0]));    relay_conn far_7_7373_0_b(.in(layer_6[63]), .out(far_7_7373_0[1]));
    assign out[233] = ~far_7_7373_0[0]; 
    assign out[234] = layer_6[616] & ~layer_6[599]; 
    wire [1:0] far_7_7375_0;    relay_conn far_7_7375_0_a(.in(layer_6[332]), .out(far_7_7375_0[0]));    relay_conn far_7_7375_0_b(.in(layer_6[369]), .out(far_7_7375_0[1]));
    assign out[235] = ~far_7_7375_0[0]; 
    wire [1:0] far_7_7376_0;    relay_conn far_7_7376_0_a(.in(layer_6[558]), .out(far_7_7376_0[0]));    relay_conn far_7_7376_0_b(.in(layer_6[615]), .out(far_7_7376_0[1]));
    assign out[236] = far_7_7376_0[1] & ~far_7_7376_0[0]; 
    wire [1:0] far_7_7377_0;    relay_conn far_7_7377_0_a(.in(layer_6[141]), .out(far_7_7377_0[0]));    relay_conn far_7_7377_0_b(.in(layer_6[40]), .out(far_7_7377_0[1]));
    wire [1:0] far_7_7377_1;    relay_conn far_7_7377_1_a(.in(far_7_7377_0[0]), .out(far_7_7377_1[0]));    relay_conn far_7_7377_1_b(.in(far_7_7377_0[1]), .out(far_7_7377_1[1]));
    wire [1:0] far_7_7377_2;    relay_conn far_7_7377_2_a(.in(far_7_7377_1[0]), .out(far_7_7377_2[0]));    relay_conn far_7_7377_2_b(.in(far_7_7377_1[1]), .out(far_7_7377_2[1]));
    assign out[237] = far_7_7377_2[0] ^ far_7_7377_2[1]; 
    wire [1:0] far_7_7378_0;    relay_conn far_7_7378_0_a(.in(layer_6[317]), .out(far_7_7378_0[0]));    relay_conn far_7_7378_0_b(.in(layer_6[228]), .out(far_7_7378_0[1]));
    wire [1:0] far_7_7378_1;    relay_conn far_7_7378_1_a(.in(far_7_7378_0[0]), .out(far_7_7378_1[0]));    relay_conn far_7_7378_1_b(.in(far_7_7378_0[1]), .out(far_7_7378_1[1]));
    assign out[238] = far_7_7378_1[0] | far_7_7378_1[1]; 
    assign out[239] = layer_6[274] & layer_6[293]; 
    wire [1:0] far_7_7380_0;    relay_conn far_7_7380_0_a(.in(layer_6[828]), .out(far_7_7380_0[0]));    relay_conn far_7_7380_0_b(.in(layer_6[716]), .out(far_7_7380_0[1]));
    wire [1:0] far_7_7380_1;    relay_conn far_7_7380_1_a(.in(far_7_7380_0[0]), .out(far_7_7380_1[0]));    relay_conn far_7_7380_1_b(.in(far_7_7380_0[1]), .out(far_7_7380_1[1]));
    wire [1:0] far_7_7380_2;    relay_conn far_7_7380_2_a(.in(far_7_7380_1[0]), .out(far_7_7380_2[0]));    relay_conn far_7_7380_2_b(.in(far_7_7380_1[1]), .out(far_7_7380_2[1]));
    assign out[240] = ~far_7_7380_2[1]; 
    wire [1:0] far_7_7381_0;    relay_conn far_7_7381_0_a(.in(layer_6[624]), .out(far_7_7381_0[0]));    relay_conn far_7_7381_0_b(.in(layer_6[547]), .out(far_7_7381_0[1]));
    wire [1:0] far_7_7381_1;    relay_conn far_7_7381_1_a(.in(far_7_7381_0[0]), .out(far_7_7381_1[0]));    relay_conn far_7_7381_1_b(.in(far_7_7381_0[1]), .out(far_7_7381_1[1]));
    assign out[241] = ~far_7_7381_1[0]; 
    wire [1:0] far_7_7382_0;    relay_conn far_7_7382_0_a(.in(layer_6[318]), .out(far_7_7382_0[0]));    relay_conn far_7_7382_0_b(.in(layer_6[370]), .out(far_7_7382_0[1]));
    assign out[242] = far_7_7382_0[1]; 
    wire [1:0] far_7_7383_0;    relay_conn far_7_7383_0_a(.in(layer_6[884]), .out(far_7_7383_0[0]));    relay_conn far_7_7383_0_b(.in(layer_6[789]), .out(far_7_7383_0[1]));
    wire [1:0] far_7_7383_1;    relay_conn far_7_7383_1_a(.in(far_7_7383_0[0]), .out(far_7_7383_1[0]));    relay_conn far_7_7383_1_b(.in(far_7_7383_0[1]), .out(far_7_7383_1[1]));
    assign out[243] = ~(far_7_7383_1[0] | far_7_7383_1[1]); 
    wire [1:0] far_7_7384_0;    relay_conn far_7_7384_0_a(.in(layer_6[404]), .out(far_7_7384_0[0]));    relay_conn far_7_7384_0_b(.in(layer_6[449]), .out(far_7_7384_0[1]));
    assign out[244] = far_7_7384_0[0] & ~far_7_7384_0[1]; 
    wire [1:0] far_7_7385_0;    relay_conn far_7_7385_0_a(.in(layer_6[333]), .out(far_7_7385_0[0]));    relay_conn far_7_7385_0_b(.in(layer_6[396]), .out(far_7_7385_0[1]));
    assign out[245] = far_7_7385_0[0] | far_7_7385_0[1]; 
    wire [1:0] far_7_7386_0;    relay_conn far_7_7386_0_a(.in(layer_6[924]), .out(far_7_7386_0[0]));    relay_conn far_7_7386_0_b(.in(layer_6[991]), .out(far_7_7386_0[1]));
    wire [1:0] far_7_7386_1;    relay_conn far_7_7386_1_a(.in(far_7_7386_0[0]), .out(far_7_7386_1[0]));    relay_conn far_7_7386_1_b(.in(far_7_7386_0[1]), .out(far_7_7386_1[1]));
    assign out[246] = far_7_7386_1[1] & ~far_7_7386_1[0]; 
    assign out[247] = layer_6[208] ^ layer_6[198]; 
    wire [1:0] far_7_7388_0;    relay_conn far_7_7388_0_a(.in(layer_6[7]), .out(far_7_7388_0[0]));    relay_conn far_7_7388_0_b(.in(layer_6[110]), .out(far_7_7388_0[1]));
    wire [1:0] far_7_7388_1;    relay_conn far_7_7388_1_a(.in(far_7_7388_0[0]), .out(far_7_7388_1[0]));    relay_conn far_7_7388_1_b(.in(far_7_7388_0[1]), .out(far_7_7388_1[1]));
    wire [1:0] far_7_7388_2;    relay_conn far_7_7388_2_a(.in(far_7_7388_1[0]), .out(far_7_7388_2[0]));    relay_conn far_7_7388_2_b(.in(far_7_7388_1[1]), .out(far_7_7388_2[1]));
    assign out[248] = far_7_7388_2[1]; 
    wire [1:0] far_7_7389_0;    relay_conn far_7_7389_0_a(.in(layer_6[88]), .out(far_7_7389_0[0]));    relay_conn far_7_7389_0_b(.in(layer_6[176]), .out(far_7_7389_0[1]));
    wire [1:0] far_7_7389_1;    relay_conn far_7_7389_1_a(.in(far_7_7389_0[0]), .out(far_7_7389_1[0]));    relay_conn far_7_7389_1_b(.in(far_7_7389_0[1]), .out(far_7_7389_1[1]));
    assign out[249] = ~far_7_7389_1[1]; 
    wire [1:0] far_7_7390_0;    relay_conn far_7_7390_0_a(.in(layer_6[76]), .out(far_7_7390_0[0]));    relay_conn far_7_7390_0_b(.in(layer_6[138]), .out(far_7_7390_0[1]));
    assign out[250] = ~(far_7_7390_0[0] ^ far_7_7390_0[1]); 
    assign out[251] = ~layer_6[403]; 
    wire [1:0] far_7_7392_0;    relay_conn far_7_7392_0_a(.in(layer_6[57]), .out(far_7_7392_0[0]));    relay_conn far_7_7392_0_b(.in(layer_6[98]), .out(far_7_7392_0[1]));
    assign out[252] = far_7_7392_0[0]; 
    wire [1:0] far_7_7393_0;    relay_conn far_7_7393_0_a(.in(layer_6[966]), .out(far_7_7393_0[0]));    relay_conn far_7_7393_0_b(.in(layer_6[920]), .out(far_7_7393_0[1]));
    assign out[253] = far_7_7393_0[0]; 
    wire [1:0] far_7_7394_0;    relay_conn far_7_7394_0_a(.in(layer_6[887]), .out(far_7_7394_0[0]));    relay_conn far_7_7394_0_b(.in(layer_6[972]), .out(far_7_7394_0[1]));
    wire [1:0] far_7_7394_1;    relay_conn far_7_7394_1_a(.in(far_7_7394_0[0]), .out(far_7_7394_1[0]));    relay_conn far_7_7394_1_b(.in(far_7_7394_0[1]), .out(far_7_7394_1[1]));
    assign out[254] = ~(far_7_7394_1[0] ^ far_7_7394_1[1]); 
    wire [1:0] far_7_7395_0;    relay_conn far_7_7395_0_a(.in(layer_6[318]), .out(far_7_7395_0[0]));    relay_conn far_7_7395_0_b(.in(layer_6[207]), .out(far_7_7395_0[1]));
    wire [1:0] far_7_7395_1;    relay_conn far_7_7395_1_a(.in(far_7_7395_0[0]), .out(far_7_7395_1[0]));    relay_conn far_7_7395_1_b(.in(far_7_7395_0[1]), .out(far_7_7395_1[1]));
    wire [1:0] far_7_7395_2;    relay_conn far_7_7395_2_a(.in(far_7_7395_1[0]), .out(far_7_7395_2[0]));    relay_conn far_7_7395_2_b(.in(far_7_7395_1[1]), .out(far_7_7395_2[1]));
    assign out[255] = ~(far_7_7395_2[0] ^ far_7_7395_2[1]); 
    assign out[256] = ~(layer_6[802] | layer_6[774]); 
    wire [1:0] far_7_7397_0;    relay_conn far_7_7397_0_a(.in(layer_6[792]), .out(far_7_7397_0[0]));    relay_conn far_7_7397_0_b(.in(layer_6[895]), .out(far_7_7397_0[1]));
    wire [1:0] far_7_7397_1;    relay_conn far_7_7397_1_a(.in(far_7_7397_0[0]), .out(far_7_7397_1[0]));    relay_conn far_7_7397_1_b(.in(far_7_7397_0[1]), .out(far_7_7397_1[1]));
    wire [1:0] far_7_7397_2;    relay_conn far_7_7397_2_a(.in(far_7_7397_1[0]), .out(far_7_7397_2[0]));    relay_conn far_7_7397_2_b(.in(far_7_7397_1[1]), .out(far_7_7397_2[1]));
    assign out[257] = far_7_7397_2[0]; 
    assign out[258] = ~layer_6[930]; 
    wire [1:0] far_7_7399_0;    relay_conn far_7_7399_0_a(.in(layer_6[109]), .out(far_7_7399_0[0]));    relay_conn far_7_7399_0_b(.in(layer_6[71]), .out(far_7_7399_0[1]));
    assign out[259] = far_7_7399_0[1] & ~far_7_7399_0[0]; 
    wire [1:0] far_7_7400_0;    relay_conn far_7_7400_0_a(.in(layer_6[712]), .out(far_7_7400_0[0]));    relay_conn far_7_7400_0_b(.in(layer_6[676]), .out(far_7_7400_0[1]));
    assign out[260] = ~(far_7_7400_0[0] ^ far_7_7400_0[1]); 
    assign out[261] = ~(layer_6[601] ^ layer_6[597]); 
    assign out[262] = ~layer_6[778]; 
    assign out[263] = layer_6[324]; 
    wire [1:0] far_7_7404_0;    relay_conn far_7_7404_0_a(.in(layer_6[732]), .out(far_7_7404_0[0]));    relay_conn far_7_7404_0_b(.in(layer_6[840]), .out(far_7_7404_0[1]));
    wire [1:0] far_7_7404_1;    relay_conn far_7_7404_1_a(.in(far_7_7404_0[0]), .out(far_7_7404_1[0]));    relay_conn far_7_7404_1_b(.in(far_7_7404_0[1]), .out(far_7_7404_1[1]));
    wire [1:0] far_7_7404_2;    relay_conn far_7_7404_2_a(.in(far_7_7404_1[0]), .out(far_7_7404_2[0]));    relay_conn far_7_7404_2_b(.in(far_7_7404_1[1]), .out(far_7_7404_2[1]));
    assign out[264] = ~far_7_7404_2[0]; 
    assign out[265] = ~layer_6[387]; 
    assign out[266] = ~layer_6[68]; 
    assign out[267] = ~layer_6[1011]; 
    assign out[268] = layer_6[613] ^ layer_6[597]; 
    assign out[269] = layer_6[744]; 
    wire [1:0] far_7_7410_0;    relay_conn far_7_7410_0_a(.in(layer_6[673]), .out(far_7_7410_0[0]));    relay_conn far_7_7410_0_b(.in(layer_6[569]), .out(far_7_7410_0[1]));
    wire [1:0] far_7_7410_1;    relay_conn far_7_7410_1_a(.in(far_7_7410_0[0]), .out(far_7_7410_1[0]));    relay_conn far_7_7410_1_b(.in(far_7_7410_0[1]), .out(far_7_7410_1[1]));
    wire [1:0] far_7_7410_2;    relay_conn far_7_7410_2_a(.in(far_7_7410_1[0]), .out(far_7_7410_2[0]));    relay_conn far_7_7410_2_b(.in(far_7_7410_1[1]), .out(far_7_7410_2[1]));
    assign out[270] = ~far_7_7410_2[0]; 
    assign out[271] = ~layer_6[251]; 
    wire [1:0] far_7_7412_0;    relay_conn far_7_7412_0_a(.in(layer_6[931]), .out(far_7_7412_0[0]));    relay_conn far_7_7412_0_b(.in(layer_6[981]), .out(far_7_7412_0[1]));
    assign out[272] = ~far_7_7412_0[0] | (far_7_7412_0[0] & far_7_7412_0[1]); 
    wire [1:0] far_7_7413_0;    relay_conn far_7_7413_0_a(.in(layer_6[522]), .out(far_7_7413_0[0]));    relay_conn far_7_7413_0_b(.in(layer_6[586]), .out(far_7_7413_0[1]));
    wire [1:0] far_7_7413_1;    relay_conn far_7_7413_1_a(.in(far_7_7413_0[0]), .out(far_7_7413_1[0]));    relay_conn far_7_7413_1_b(.in(far_7_7413_0[1]), .out(far_7_7413_1[1]));
    assign out[273] = ~(far_7_7413_1[0] ^ far_7_7413_1[1]); 
    wire [1:0] far_7_7414_0;    relay_conn far_7_7414_0_a(.in(layer_6[755]), .out(far_7_7414_0[0]));    relay_conn far_7_7414_0_b(.in(layer_6[821]), .out(far_7_7414_0[1]));
    wire [1:0] far_7_7414_1;    relay_conn far_7_7414_1_a(.in(far_7_7414_0[0]), .out(far_7_7414_1[0]));    relay_conn far_7_7414_1_b(.in(far_7_7414_0[1]), .out(far_7_7414_1[1]));
    assign out[274] = far_7_7414_1[0] & ~far_7_7414_1[1]; 
    assign out[275] = layer_6[852] & ~layer_6[836]; 
    wire [1:0] far_7_7416_0;    relay_conn far_7_7416_0_a(.in(layer_6[468]), .out(far_7_7416_0[0]));    relay_conn far_7_7416_0_b(.in(layer_6[435]), .out(far_7_7416_0[1]));
    assign out[276] = ~(far_7_7416_0[0] | far_7_7416_0[1]); 
    wire [1:0] far_7_7417_0;    relay_conn far_7_7417_0_a(.in(layer_6[553]), .out(far_7_7417_0[0]));    relay_conn far_7_7417_0_b(.in(layer_6[449]), .out(far_7_7417_0[1]));
    wire [1:0] far_7_7417_1;    relay_conn far_7_7417_1_a(.in(far_7_7417_0[0]), .out(far_7_7417_1[0]));    relay_conn far_7_7417_1_b(.in(far_7_7417_0[1]), .out(far_7_7417_1[1]));
    wire [1:0] far_7_7417_2;    relay_conn far_7_7417_2_a(.in(far_7_7417_1[0]), .out(far_7_7417_2[0]));    relay_conn far_7_7417_2_b(.in(far_7_7417_1[1]), .out(far_7_7417_2[1]));
    assign out[277] = far_7_7417_2[0] & ~far_7_7417_2[1]; 
    wire [1:0] far_7_7418_0;    relay_conn far_7_7418_0_a(.in(layer_6[628]), .out(far_7_7418_0[0]));    relay_conn far_7_7418_0_b(.in(layer_6[557]), .out(far_7_7418_0[1]));
    wire [1:0] far_7_7418_1;    relay_conn far_7_7418_1_a(.in(far_7_7418_0[0]), .out(far_7_7418_1[0]));    relay_conn far_7_7418_1_b(.in(far_7_7418_0[1]), .out(far_7_7418_1[1]));
    assign out[278] = far_7_7418_1[0] & far_7_7418_1[1]; 
    wire [1:0] far_7_7419_0;    relay_conn far_7_7419_0_a(.in(layer_6[923]), .out(far_7_7419_0[0]));    relay_conn far_7_7419_0_b(.in(layer_6[884]), .out(far_7_7419_0[1]));
    assign out[279] = far_7_7419_0[0] & ~far_7_7419_0[1]; 
    wire [1:0] far_7_7420_0;    relay_conn far_7_7420_0_a(.in(layer_6[449]), .out(far_7_7420_0[0]));    relay_conn far_7_7420_0_b(.in(layer_6[534]), .out(far_7_7420_0[1]));
    wire [1:0] far_7_7420_1;    relay_conn far_7_7420_1_a(.in(far_7_7420_0[0]), .out(far_7_7420_1[0]));    relay_conn far_7_7420_1_b(.in(far_7_7420_0[1]), .out(far_7_7420_1[1]));
    assign out[280] = ~(far_7_7420_1[0] | far_7_7420_1[1]); 
    wire [1:0] far_7_7421_0;    relay_conn far_7_7421_0_a(.in(layer_6[597]), .out(far_7_7421_0[0]));    relay_conn far_7_7421_0_b(.in(layer_6[692]), .out(far_7_7421_0[1]));
    wire [1:0] far_7_7421_1;    relay_conn far_7_7421_1_a(.in(far_7_7421_0[0]), .out(far_7_7421_1[0]));    relay_conn far_7_7421_1_b(.in(far_7_7421_0[1]), .out(far_7_7421_1[1]));
    assign out[281] = ~far_7_7421_1[1]; 
    wire [1:0] far_7_7422_0;    relay_conn far_7_7422_0_a(.in(layer_6[222]), .out(far_7_7422_0[0]));    relay_conn far_7_7422_0_b(.in(layer_6[345]), .out(far_7_7422_0[1]));
    wire [1:0] far_7_7422_1;    relay_conn far_7_7422_1_a(.in(far_7_7422_0[0]), .out(far_7_7422_1[0]));    relay_conn far_7_7422_1_b(.in(far_7_7422_0[1]), .out(far_7_7422_1[1]));
    wire [1:0] far_7_7422_2;    relay_conn far_7_7422_2_a(.in(far_7_7422_1[0]), .out(far_7_7422_2[0]));    relay_conn far_7_7422_2_b(.in(far_7_7422_1[1]), .out(far_7_7422_2[1]));
    assign out[282] = ~(far_7_7422_2[0] | far_7_7422_2[1]); 
    wire [1:0] far_7_7423_0;    relay_conn far_7_7423_0_a(.in(layer_6[967]), .out(far_7_7423_0[0]));    relay_conn far_7_7423_0_b(.in(layer_6[1011]), .out(far_7_7423_0[1]));
    assign out[283] = far_7_7423_0[0] & ~far_7_7423_0[1]; 
    wire [1:0] far_7_7424_0;    relay_conn far_7_7424_0_a(.in(layer_6[496]), .out(far_7_7424_0[0]));    relay_conn far_7_7424_0_b(.in(layer_6[449]), .out(far_7_7424_0[1]));
    assign out[284] = ~(far_7_7424_0[0] | far_7_7424_0[1]); 
    assign out[285] = ~layer_6[84]; 
    assign out[286] = layer_6[773] & ~layer_6[777]; 
    wire [1:0] far_7_7427_0;    relay_conn far_7_7427_0_a(.in(layer_6[920]), .out(far_7_7427_0[0]));    relay_conn far_7_7427_0_b(.in(layer_6[845]), .out(far_7_7427_0[1]));
    wire [1:0] far_7_7427_1;    relay_conn far_7_7427_1_a(.in(far_7_7427_0[0]), .out(far_7_7427_1[0]));    relay_conn far_7_7427_1_b(.in(far_7_7427_0[1]), .out(far_7_7427_1[1]));
    assign out[287] = far_7_7427_1[0] & far_7_7427_1[1]; 
    wire [1:0] far_7_7428_0;    relay_conn far_7_7428_0_a(.in(layer_6[746]), .out(far_7_7428_0[0]));    relay_conn far_7_7428_0_b(.in(layer_6[672]), .out(far_7_7428_0[1]));
    wire [1:0] far_7_7428_1;    relay_conn far_7_7428_1_a(.in(far_7_7428_0[0]), .out(far_7_7428_1[0]));    relay_conn far_7_7428_1_b(.in(far_7_7428_0[1]), .out(far_7_7428_1[1]));
    assign out[288] = far_7_7428_1[1]; 
    wire [1:0] far_7_7429_0;    relay_conn far_7_7429_0_a(.in(layer_6[703]), .out(far_7_7429_0[0]));    relay_conn far_7_7429_0_b(.in(layer_6[633]), .out(far_7_7429_0[1]));
    wire [1:0] far_7_7429_1;    relay_conn far_7_7429_1_a(.in(far_7_7429_0[0]), .out(far_7_7429_1[0]));    relay_conn far_7_7429_1_b(.in(far_7_7429_0[1]), .out(far_7_7429_1[1]));
    assign out[289] = far_7_7429_1[0]; 
    wire [1:0] far_7_7430_0;    relay_conn far_7_7430_0_a(.in(layer_6[829]), .out(far_7_7430_0[0]));    relay_conn far_7_7430_0_b(.in(layer_6[789]), .out(far_7_7430_0[1]));
    assign out[290] = ~far_7_7430_0[1]; 
    wire [1:0] far_7_7431_0;    relay_conn far_7_7431_0_a(.in(layer_6[742]), .out(far_7_7431_0[0]));    relay_conn far_7_7431_0_b(.in(layer_6[683]), .out(far_7_7431_0[1]));
    assign out[291] = far_7_7431_0[0] & ~far_7_7431_0[1]; 
    assign out[292] = layer_6[773]; 
    wire [1:0] far_7_7433_0;    relay_conn far_7_7433_0_a(.in(layer_6[985]), .out(far_7_7433_0[0]));    relay_conn far_7_7433_0_b(.in(layer_6[908]), .out(far_7_7433_0[1]));
    wire [1:0] far_7_7433_1;    relay_conn far_7_7433_1_a(.in(far_7_7433_0[0]), .out(far_7_7433_1[0]));    relay_conn far_7_7433_1_b(.in(far_7_7433_0[1]), .out(far_7_7433_1[1]));
    assign out[293] = far_7_7433_1[0]; 
    wire [1:0] far_7_7434_0;    relay_conn far_7_7434_0_a(.in(layer_6[706]), .out(far_7_7434_0[0]));    relay_conn far_7_7434_0_b(.in(layer_6[600]), .out(far_7_7434_0[1]));
    wire [1:0] far_7_7434_1;    relay_conn far_7_7434_1_a(.in(far_7_7434_0[0]), .out(far_7_7434_1[0]));    relay_conn far_7_7434_1_b(.in(far_7_7434_0[1]), .out(far_7_7434_1[1]));
    wire [1:0] far_7_7434_2;    relay_conn far_7_7434_2_a(.in(far_7_7434_1[0]), .out(far_7_7434_2[0]));    relay_conn far_7_7434_2_b(.in(far_7_7434_1[1]), .out(far_7_7434_2[1]));
    assign out[294] = ~(far_7_7434_2[0] ^ far_7_7434_2[1]); 
    wire [1:0] far_7_7435_0;    relay_conn far_7_7435_0_a(.in(layer_6[416]), .out(far_7_7435_0[0]));    relay_conn far_7_7435_0_b(.in(layer_6[450]), .out(far_7_7435_0[1]));
    assign out[295] = far_7_7435_0[1]; 
    wire [1:0] far_7_7436_0;    relay_conn far_7_7436_0_a(.in(layer_6[282]), .out(far_7_7436_0[0]));    relay_conn far_7_7436_0_b(.in(layer_6[330]), .out(far_7_7436_0[1]));
    assign out[296] = far_7_7436_0[0] & far_7_7436_0[1]; 
    wire [1:0] far_7_7437_0;    relay_conn far_7_7437_0_a(.in(layer_6[720]), .out(far_7_7437_0[0]));    relay_conn far_7_7437_0_b(.in(layer_6[799]), .out(far_7_7437_0[1]));
    wire [1:0] far_7_7437_1;    relay_conn far_7_7437_1_a(.in(far_7_7437_0[0]), .out(far_7_7437_1[0]));    relay_conn far_7_7437_1_b(.in(far_7_7437_0[1]), .out(far_7_7437_1[1]));
    assign out[297] = far_7_7437_1[0] & ~far_7_7437_1[1]; 
    wire [1:0] far_7_7438_0;    relay_conn far_7_7438_0_a(.in(layer_6[623]), .out(far_7_7438_0[0]));    relay_conn far_7_7438_0_b(.in(layer_6[575]), .out(far_7_7438_0[1]));
    assign out[298] = far_7_7438_0[1]; 
    wire [1:0] far_7_7439_0;    relay_conn far_7_7439_0_a(.in(layer_6[774]), .out(far_7_7439_0[0]));    relay_conn far_7_7439_0_b(.in(layer_6[861]), .out(far_7_7439_0[1]));
    wire [1:0] far_7_7439_1;    relay_conn far_7_7439_1_a(.in(far_7_7439_0[0]), .out(far_7_7439_1[0]));    relay_conn far_7_7439_1_b(.in(far_7_7439_0[1]), .out(far_7_7439_1[1]));
    assign out[299] = far_7_7439_1[1]; 
    wire [1:0] far_7_7440_0;    relay_conn far_7_7440_0_a(.in(layer_6[451]), .out(far_7_7440_0[0]));    relay_conn far_7_7440_0_b(.in(layer_6[552]), .out(far_7_7440_0[1]));
    wire [1:0] far_7_7440_1;    relay_conn far_7_7440_1_a(.in(far_7_7440_0[0]), .out(far_7_7440_1[0]));    relay_conn far_7_7440_1_b(.in(far_7_7440_0[1]), .out(far_7_7440_1[1]));
    wire [1:0] far_7_7440_2;    relay_conn far_7_7440_2_a(.in(far_7_7440_1[0]), .out(far_7_7440_2[0]));    relay_conn far_7_7440_2_b(.in(far_7_7440_1[1]), .out(far_7_7440_2[1]));
    assign out[300] = far_7_7440_2[1] & ~far_7_7440_2[0]; 
    wire [1:0] far_7_7441_0;    relay_conn far_7_7441_0_a(.in(layer_6[393]), .out(far_7_7441_0[0]));    relay_conn far_7_7441_0_b(.in(layer_6[271]), .out(far_7_7441_0[1]));
    wire [1:0] far_7_7441_1;    relay_conn far_7_7441_1_a(.in(far_7_7441_0[0]), .out(far_7_7441_1[0]));    relay_conn far_7_7441_1_b(.in(far_7_7441_0[1]), .out(far_7_7441_1[1]));
    wire [1:0] far_7_7441_2;    relay_conn far_7_7441_2_a(.in(far_7_7441_1[0]), .out(far_7_7441_2[0]));    relay_conn far_7_7441_2_b(.in(far_7_7441_1[1]), .out(far_7_7441_2[1]));
    assign out[301] = far_7_7441_2[0] ^ far_7_7441_2[1]; 
    wire [1:0] far_7_7442_0;    relay_conn far_7_7442_0_a(.in(layer_6[136]), .out(far_7_7442_0[0]));    relay_conn far_7_7442_0_b(.in(layer_6[26]), .out(far_7_7442_0[1]));
    wire [1:0] far_7_7442_1;    relay_conn far_7_7442_1_a(.in(far_7_7442_0[0]), .out(far_7_7442_1[0]));    relay_conn far_7_7442_1_b(.in(far_7_7442_0[1]), .out(far_7_7442_1[1]));
    wire [1:0] far_7_7442_2;    relay_conn far_7_7442_2_a(.in(far_7_7442_1[0]), .out(far_7_7442_2[0]));    relay_conn far_7_7442_2_b(.in(far_7_7442_1[1]), .out(far_7_7442_2[1]));
    assign out[302] = ~(far_7_7442_2[0] | far_7_7442_2[1]); 
    wire [1:0] far_7_7443_0;    relay_conn far_7_7443_0_a(.in(layer_6[336]), .out(far_7_7443_0[0]));    relay_conn far_7_7443_0_b(.in(layer_6[279]), .out(far_7_7443_0[1]));
    assign out[303] = far_7_7443_0[1]; 
    assign out[304] = ~(layer_6[413] | layer_6[440]); 
    wire [1:0] far_7_7445_0;    relay_conn far_7_7445_0_a(.in(layer_6[659]), .out(far_7_7445_0[0]));    relay_conn far_7_7445_0_b(.in(layer_6[763]), .out(far_7_7445_0[1]));
    wire [1:0] far_7_7445_1;    relay_conn far_7_7445_1_a(.in(far_7_7445_0[0]), .out(far_7_7445_1[0]));    relay_conn far_7_7445_1_b(.in(far_7_7445_0[1]), .out(far_7_7445_1[1]));
    wire [1:0] far_7_7445_2;    relay_conn far_7_7445_2_a(.in(far_7_7445_1[0]), .out(far_7_7445_2[0]));    relay_conn far_7_7445_2_b(.in(far_7_7445_1[1]), .out(far_7_7445_2[1]));
    assign out[305] = ~far_7_7445_2[1]; 
    assign out[306] = layer_6[312]; 
    wire [1:0] far_7_7447_0;    relay_conn far_7_7447_0_a(.in(layer_6[237]), .out(far_7_7447_0[0]));    relay_conn far_7_7447_0_b(.in(layer_6[145]), .out(far_7_7447_0[1]));
    wire [1:0] far_7_7447_1;    relay_conn far_7_7447_1_a(.in(far_7_7447_0[0]), .out(far_7_7447_1[0]));    relay_conn far_7_7447_1_b(.in(far_7_7447_0[1]), .out(far_7_7447_1[1]));
    assign out[307] = far_7_7447_1[0] ^ far_7_7447_1[1]; 
    assign out[308] = ~layer_6[947]; 
    wire [1:0] far_7_7449_0;    relay_conn far_7_7449_0_a(.in(layer_6[51]), .out(far_7_7449_0[0]));    relay_conn far_7_7449_0_b(.in(layer_6[19]), .out(far_7_7449_0[1]));
    assign out[309] = ~(far_7_7449_0[0] ^ far_7_7449_0[1]); 
    assign out[310] = ~layer_6[750]; 
    assign out[311] = layer_6[771] & layer_6[755]; 
    assign out[312] = ~layer_6[187] | (layer_6[187] & layer_6[208]); 
    wire [1:0] far_7_7453_0;    relay_conn far_7_7453_0_a(.in(layer_6[146]), .out(far_7_7453_0[0]));    relay_conn far_7_7453_0_b(.in(layer_6[210]), .out(far_7_7453_0[1]));
    wire [1:0] far_7_7453_1;    relay_conn far_7_7453_1_a(.in(far_7_7453_0[0]), .out(far_7_7453_1[0]));    relay_conn far_7_7453_1_b(.in(far_7_7453_0[1]), .out(far_7_7453_1[1]));
    assign out[313] = ~(far_7_7453_1[0] | far_7_7453_1[1]); 
    wire [1:0] far_7_7454_0;    relay_conn far_7_7454_0_a(.in(layer_6[214]), .out(far_7_7454_0[0]));    relay_conn far_7_7454_0_b(.in(layer_6[117]), .out(far_7_7454_0[1]));
    wire [1:0] far_7_7454_1;    relay_conn far_7_7454_1_a(.in(far_7_7454_0[0]), .out(far_7_7454_1[0]));    relay_conn far_7_7454_1_b(.in(far_7_7454_0[1]), .out(far_7_7454_1[1]));
    wire [1:0] far_7_7454_2;    relay_conn far_7_7454_2_a(.in(far_7_7454_1[0]), .out(far_7_7454_2[0]));    relay_conn far_7_7454_2_b(.in(far_7_7454_1[1]), .out(far_7_7454_2[1]));
    assign out[314] = ~(far_7_7454_2[0] | far_7_7454_2[1]); 
    wire [1:0] far_7_7455_0;    relay_conn far_7_7455_0_a(.in(layer_6[128]), .out(far_7_7455_0[0]));    relay_conn far_7_7455_0_b(.in(layer_6[84]), .out(far_7_7455_0[1]));
    assign out[315] = far_7_7455_0[0] & far_7_7455_0[1]; 
    wire [1:0] far_7_7456_0;    relay_conn far_7_7456_0_a(.in(layer_6[505]), .out(far_7_7456_0[0]));    relay_conn far_7_7456_0_b(.in(layer_6[432]), .out(far_7_7456_0[1]));
    wire [1:0] far_7_7456_1;    relay_conn far_7_7456_1_a(.in(far_7_7456_0[0]), .out(far_7_7456_1[0]));    relay_conn far_7_7456_1_b(.in(far_7_7456_0[1]), .out(far_7_7456_1[1]));
    assign out[316] = far_7_7456_1[1]; 
    wire [1:0] far_7_7457_0;    relay_conn far_7_7457_0_a(.in(layer_6[214]), .out(far_7_7457_0[0]));    relay_conn far_7_7457_0_b(.in(layer_6[162]), .out(far_7_7457_0[1]));
    assign out[317] = far_7_7457_0[1] & ~far_7_7457_0[0]; 
    assign out[318] = ~layer_6[386]; 
    wire [1:0] far_7_7459_0;    relay_conn far_7_7459_0_a(.in(layer_6[931]), .out(far_7_7459_0[0]));    relay_conn far_7_7459_0_b(.in(layer_6[815]), .out(far_7_7459_0[1]));
    wire [1:0] far_7_7459_1;    relay_conn far_7_7459_1_a(.in(far_7_7459_0[0]), .out(far_7_7459_1[0]));    relay_conn far_7_7459_1_b(.in(far_7_7459_0[1]), .out(far_7_7459_1[1]));
    wire [1:0] far_7_7459_2;    relay_conn far_7_7459_2_a(.in(far_7_7459_1[0]), .out(far_7_7459_2[0]));    relay_conn far_7_7459_2_b(.in(far_7_7459_1[1]), .out(far_7_7459_2[1]));
    assign out[319] = ~far_7_7459_2[0] | (far_7_7459_2[0] & far_7_7459_2[1]); 
    assign out[320] = layer_6[198] & layer_6[211]; 
    wire [1:0] far_7_7461_0;    relay_conn far_7_7461_0_a(.in(layer_6[329]), .out(far_7_7461_0[0]));    relay_conn far_7_7461_0_b(.in(layer_6[394]), .out(far_7_7461_0[1]));
    wire [1:0] far_7_7461_1;    relay_conn far_7_7461_1_a(.in(far_7_7461_0[0]), .out(far_7_7461_1[0]));    relay_conn far_7_7461_1_b(.in(far_7_7461_0[1]), .out(far_7_7461_1[1]));
    assign out[321] = ~(far_7_7461_1[0] ^ far_7_7461_1[1]); 
    assign out[322] = ~layer_6[777]; 
    assign out[323] = ~(layer_6[622] | layer_6[648]); 
    wire [1:0] far_7_7464_0;    relay_conn far_7_7464_0_a(.in(layer_6[646]), .out(far_7_7464_0[0]));    relay_conn far_7_7464_0_b(.in(layer_6[524]), .out(far_7_7464_0[1]));
    wire [1:0] far_7_7464_1;    relay_conn far_7_7464_1_a(.in(far_7_7464_0[0]), .out(far_7_7464_1[0]));    relay_conn far_7_7464_1_b(.in(far_7_7464_0[1]), .out(far_7_7464_1[1]));
    wire [1:0] far_7_7464_2;    relay_conn far_7_7464_2_a(.in(far_7_7464_1[0]), .out(far_7_7464_2[0]));    relay_conn far_7_7464_2_b(.in(far_7_7464_1[1]), .out(far_7_7464_2[1]));
    assign out[324] = far_7_7464_2[0] & ~far_7_7464_2[1]; 
    wire [1:0] far_7_7465_0;    relay_conn far_7_7465_0_a(.in(layer_6[256]), .out(far_7_7465_0[0]));    relay_conn far_7_7465_0_b(.in(layer_6[321]), .out(far_7_7465_0[1]));
    wire [1:0] far_7_7465_1;    relay_conn far_7_7465_1_a(.in(far_7_7465_0[0]), .out(far_7_7465_1[0]));    relay_conn far_7_7465_1_b(.in(far_7_7465_0[1]), .out(far_7_7465_1[1]));
    assign out[325] = far_7_7465_1[0] | far_7_7465_1[1]; 
    wire [1:0] far_7_7466_0;    relay_conn far_7_7466_0_a(.in(layer_6[755]), .out(far_7_7466_0[0]));    relay_conn far_7_7466_0_b(.in(layer_6[642]), .out(far_7_7466_0[1]));
    wire [1:0] far_7_7466_1;    relay_conn far_7_7466_1_a(.in(far_7_7466_0[0]), .out(far_7_7466_1[0]));    relay_conn far_7_7466_1_b(.in(far_7_7466_0[1]), .out(far_7_7466_1[1]));
    wire [1:0] far_7_7466_2;    relay_conn far_7_7466_2_a(.in(far_7_7466_1[0]), .out(far_7_7466_2[0]));    relay_conn far_7_7466_2_b(.in(far_7_7466_1[1]), .out(far_7_7466_2[1]));
    assign out[326] = far_7_7466_2[0]; 
    wire [1:0] far_7_7467_0;    relay_conn far_7_7467_0_a(.in(layer_6[360]), .out(far_7_7467_0[0]));    relay_conn far_7_7467_0_b(.in(layer_6[271]), .out(far_7_7467_0[1]));
    wire [1:0] far_7_7467_1;    relay_conn far_7_7467_1_a(.in(far_7_7467_0[0]), .out(far_7_7467_1[0]));    relay_conn far_7_7467_1_b(.in(far_7_7467_0[1]), .out(far_7_7467_1[1]));
    assign out[327] = ~far_7_7467_1[1]; 
    wire [1:0] far_7_7468_0;    relay_conn far_7_7468_0_a(.in(layer_6[273]), .out(far_7_7468_0[0]));    relay_conn far_7_7468_0_b(.in(layer_6[320]), .out(far_7_7468_0[1]));
    assign out[328] = ~(far_7_7468_0[0] ^ far_7_7468_0[1]); 
    wire [1:0] far_7_7469_0;    relay_conn far_7_7469_0_a(.in(layer_6[93]), .out(far_7_7469_0[0]));    relay_conn far_7_7469_0_b(.in(layer_6[58]), .out(far_7_7469_0[1]));
    assign out[329] = ~far_7_7469_0[1]; 
    wire [1:0] far_7_7470_0;    relay_conn far_7_7470_0_a(.in(layer_6[750]), .out(far_7_7470_0[0]));    relay_conn far_7_7470_0_b(.in(layer_6[695]), .out(far_7_7470_0[1]));
    assign out[330] = ~far_7_7470_0[0]; 
    wire [1:0] far_7_7471_0;    relay_conn far_7_7471_0_a(.in(layer_6[497]), .out(far_7_7471_0[0]));    relay_conn far_7_7471_0_b(.in(layer_6[569]), .out(far_7_7471_0[1]));
    wire [1:0] far_7_7471_1;    relay_conn far_7_7471_1_a(.in(far_7_7471_0[0]), .out(far_7_7471_1[0]));    relay_conn far_7_7471_1_b(.in(far_7_7471_0[1]), .out(far_7_7471_1[1]));
    assign out[331] = far_7_7471_1[0] & ~far_7_7471_1[1]; 
    wire [1:0] far_7_7472_0;    relay_conn far_7_7472_0_a(.in(layer_6[329]), .out(far_7_7472_0[0]));    relay_conn far_7_7472_0_b(.in(layer_6[290]), .out(far_7_7472_0[1]));
    assign out[332] = far_7_7472_0[0] & far_7_7472_0[1]; 
    wire [1:0] far_7_7473_0;    relay_conn far_7_7473_0_a(.in(layer_6[558]), .out(far_7_7473_0[0]));    relay_conn far_7_7473_0_b(.in(layer_6[648]), .out(far_7_7473_0[1]));
    wire [1:0] far_7_7473_1;    relay_conn far_7_7473_1_a(.in(far_7_7473_0[0]), .out(far_7_7473_1[0]));    relay_conn far_7_7473_1_b(.in(far_7_7473_0[1]), .out(far_7_7473_1[1]));
    assign out[333] = far_7_7473_1[0]; 
    assign out[334] = ~layer_6[670]; 
    wire [1:0] far_7_7475_0;    relay_conn far_7_7475_0_a(.in(layer_6[632]), .out(far_7_7475_0[0]));    relay_conn far_7_7475_0_b(.in(layer_6[558]), .out(far_7_7475_0[1]));
    wire [1:0] far_7_7475_1;    relay_conn far_7_7475_1_a(.in(far_7_7475_0[0]), .out(far_7_7475_1[0]));    relay_conn far_7_7475_1_b(.in(far_7_7475_0[1]), .out(far_7_7475_1[1]));
    assign out[335] = ~(far_7_7475_1[0] ^ far_7_7475_1[1]); 
    wire [1:0] far_7_7476_0;    relay_conn far_7_7476_0_a(.in(layer_6[18]), .out(far_7_7476_0[0]));    relay_conn far_7_7476_0_b(.in(layer_6[74]), .out(far_7_7476_0[1]));
    assign out[336] = ~far_7_7476_0[0]; 
    wire [1:0] far_7_7477_0;    relay_conn far_7_7477_0_a(.in(layer_6[644]), .out(far_7_7477_0[0]));    relay_conn far_7_7477_0_b(.in(layer_6[594]), .out(far_7_7477_0[1]));
    assign out[337] = ~far_7_7477_0[0] | (far_7_7477_0[0] & far_7_7477_0[1]); 
    wire [1:0] far_7_7478_0;    relay_conn far_7_7478_0_a(.in(layer_6[361]), .out(far_7_7478_0[0]));    relay_conn far_7_7478_0_b(.in(layer_6[242]), .out(far_7_7478_0[1]));
    wire [1:0] far_7_7478_1;    relay_conn far_7_7478_1_a(.in(far_7_7478_0[0]), .out(far_7_7478_1[0]));    relay_conn far_7_7478_1_b(.in(far_7_7478_0[1]), .out(far_7_7478_1[1]));
    wire [1:0] far_7_7478_2;    relay_conn far_7_7478_2_a(.in(far_7_7478_1[0]), .out(far_7_7478_2[0]));    relay_conn far_7_7478_2_b(.in(far_7_7478_1[1]), .out(far_7_7478_2[1]));
    assign out[338] = far_7_7478_2[0]; 
    wire [1:0] far_7_7479_0;    relay_conn far_7_7479_0_a(.in(layer_6[394]), .out(far_7_7479_0[0]));    relay_conn far_7_7479_0_b(.in(layer_6[451]), .out(far_7_7479_0[1]));
    assign out[339] = ~far_7_7479_0[1]; 
    wire [1:0] far_7_7480_0;    relay_conn far_7_7480_0_a(.in(layer_6[229]), .out(far_7_7480_0[0]));    relay_conn far_7_7480_0_b(.in(layer_6[129]), .out(far_7_7480_0[1]));
    wire [1:0] far_7_7480_1;    relay_conn far_7_7480_1_a(.in(far_7_7480_0[0]), .out(far_7_7480_1[0]));    relay_conn far_7_7480_1_b(.in(far_7_7480_0[1]), .out(far_7_7480_1[1]));
    wire [1:0] far_7_7480_2;    relay_conn far_7_7480_2_a(.in(far_7_7480_1[0]), .out(far_7_7480_2[0]));    relay_conn far_7_7480_2_b(.in(far_7_7480_1[1]), .out(far_7_7480_2[1]));
    assign out[340] = ~far_7_7480_2[0] | (far_7_7480_2[0] & far_7_7480_2[1]); 
    assign out[341] = ~(layer_6[648] | layer_6[650]); 
    wire [1:0] far_7_7482_0;    relay_conn far_7_7482_0_a(.in(layer_6[781]), .out(far_7_7482_0[0]));    relay_conn far_7_7482_0_b(.in(layer_6[737]), .out(far_7_7482_0[1]));
    assign out[342] = ~far_7_7482_0[0]; 
    wire [1:0] far_7_7483_0;    relay_conn far_7_7483_0_a(.in(layer_6[574]), .out(far_7_7483_0[0]));    relay_conn far_7_7483_0_b(.in(layer_6[522]), .out(far_7_7483_0[1]));
    assign out[343] = ~far_7_7483_0[0]; 
    wire [1:0] far_7_7484_0;    relay_conn far_7_7484_0_a(.in(layer_6[497]), .out(far_7_7484_0[0]));    relay_conn far_7_7484_0_b(.in(layer_6[393]), .out(far_7_7484_0[1]));
    wire [1:0] far_7_7484_1;    relay_conn far_7_7484_1_a(.in(far_7_7484_0[0]), .out(far_7_7484_1[0]));    relay_conn far_7_7484_1_b(.in(far_7_7484_0[1]), .out(far_7_7484_1[1]));
    wire [1:0] far_7_7484_2;    relay_conn far_7_7484_2_a(.in(far_7_7484_1[0]), .out(far_7_7484_2[0]));    relay_conn far_7_7484_2_b(.in(far_7_7484_1[1]), .out(far_7_7484_2[1]));
    assign out[344] = ~(far_7_7484_2[0] ^ far_7_7484_2[1]); 
    wire [1:0] far_7_7485_0;    relay_conn far_7_7485_0_a(.in(layer_6[774]), .out(far_7_7485_0[0]));    relay_conn far_7_7485_0_b(.in(layer_6[676]), .out(far_7_7485_0[1]));
    wire [1:0] far_7_7485_1;    relay_conn far_7_7485_1_a(.in(far_7_7485_0[0]), .out(far_7_7485_1[0]));    relay_conn far_7_7485_1_b(.in(far_7_7485_0[1]), .out(far_7_7485_1[1]));
    wire [1:0] far_7_7485_2;    relay_conn far_7_7485_2_a(.in(far_7_7485_1[0]), .out(far_7_7485_2[0]));    relay_conn far_7_7485_2_b(.in(far_7_7485_1[1]), .out(far_7_7485_2[1]));
    assign out[345] = ~(far_7_7485_2[0] & far_7_7485_2[1]); 
    wire [1:0] far_7_7486_0;    relay_conn far_7_7486_0_a(.in(layer_6[840]), .out(far_7_7486_0[0]));    relay_conn far_7_7486_0_b(.in(layer_6[763]), .out(far_7_7486_0[1]));
    wire [1:0] far_7_7486_1;    relay_conn far_7_7486_1_a(.in(far_7_7486_0[0]), .out(far_7_7486_1[0]));    relay_conn far_7_7486_1_b(.in(far_7_7486_0[1]), .out(far_7_7486_1[1]));
    assign out[346] = far_7_7486_1[1]; 
    wire [1:0] far_7_7487_0;    relay_conn far_7_7487_0_a(.in(layer_6[742]), .out(far_7_7487_0[0]));    relay_conn far_7_7487_0_b(.in(layer_6[824]), .out(far_7_7487_0[1]));
    wire [1:0] far_7_7487_1;    relay_conn far_7_7487_1_a(.in(far_7_7487_0[0]), .out(far_7_7487_1[0]));    relay_conn far_7_7487_1_b(.in(far_7_7487_0[1]), .out(far_7_7487_1[1]));
    assign out[347] = far_7_7487_1[0] ^ far_7_7487_1[1]; 
    wire [1:0] far_7_7488_0;    relay_conn far_7_7488_0_a(.in(layer_6[939]), .out(far_7_7488_0[0]));    relay_conn far_7_7488_0_b(.in(layer_6[867]), .out(far_7_7488_0[1]));
    wire [1:0] far_7_7488_1;    relay_conn far_7_7488_1_a(.in(far_7_7488_0[0]), .out(far_7_7488_1[0]));    relay_conn far_7_7488_1_b(.in(far_7_7488_0[1]), .out(far_7_7488_1[1]));
    assign out[348] = far_7_7488_1[0] & ~far_7_7488_1[1]; 
    wire [1:0] far_7_7489_0;    relay_conn far_7_7489_0_a(.in(layer_6[181]), .out(far_7_7489_0[0]));    relay_conn far_7_7489_0_b(.in(layer_6[219]), .out(far_7_7489_0[1]));
    assign out[349] = far_7_7489_0[1]; 
    wire [1:0] far_7_7490_0;    relay_conn far_7_7490_0_a(.in(layer_6[229]), .out(far_7_7490_0[0]));    relay_conn far_7_7490_0_b(.in(layer_6[140]), .out(far_7_7490_0[1]));
    wire [1:0] far_7_7490_1;    relay_conn far_7_7490_1_a(.in(far_7_7490_0[0]), .out(far_7_7490_1[0]));    relay_conn far_7_7490_1_b(.in(far_7_7490_0[1]), .out(far_7_7490_1[1]));
    assign out[350] = ~far_7_7490_1[0]; 
    assign out[351] = ~(layer_6[297] & layer_6[267]); 
    wire [1:0] far_7_7492_0;    relay_conn far_7_7492_0_a(.in(layer_6[343]), .out(far_7_7492_0[0]));    relay_conn far_7_7492_0_b(.in(layer_6[456]), .out(far_7_7492_0[1]));
    wire [1:0] far_7_7492_1;    relay_conn far_7_7492_1_a(.in(far_7_7492_0[0]), .out(far_7_7492_1[0]));    relay_conn far_7_7492_1_b(.in(far_7_7492_0[1]), .out(far_7_7492_1[1]));
    wire [1:0] far_7_7492_2;    relay_conn far_7_7492_2_a(.in(far_7_7492_1[0]), .out(far_7_7492_2[0]));    relay_conn far_7_7492_2_b(.in(far_7_7492_1[1]), .out(far_7_7492_2[1]));
    assign out[352] = far_7_7492_2[1] & ~far_7_7492_2[0]; 
    wire [1:0] far_7_7493_0;    relay_conn far_7_7493_0_a(.in(layer_6[451]), .out(far_7_7493_0[0]));    relay_conn far_7_7493_0_b(.in(layer_6[326]), .out(far_7_7493_0[1]));
    wire [1:0] far_7_7493_1;    relay_conn far_7_7493_1_a(.in(far_7_7493_0[0]), .out(far_7_7493_1[0]));    relay_conn far_7_7493_1_b(.in(far_7_7493_0[1]), .out(far_7_7493_1[1]));
    wire [1:0] far_7_7493_2;    relay_conn far_7_7493_2_a(.in(far_7_7493_1[0]), .out(far_7_7493_2[0]));    relay_conn far_7_7493_2_b(.in(far_7_7493_1[1]), .out(far_7_7493_2[1]));
    assign out[353] = ~(far_7_7493_2[0] | far_7_7493_2[1]); 
    wire [1:0] far_7_7494_0;    relay_conn far_7_7494_0_a(.in(layer_6[845]), .out(far_7_7494_0[0]));    relay_conn far_7_7494_0_b(.in(layer_6[908]), .out(far_7_7494_0[1]));
    assign out[354] = far_7_7494_0[0] & far_7_7494_0[1]; 
    wire [1:0] far_7_7495_0;    relay_conn far_7_7495_0_a(.in(layer_6[39]), .out(far_7_7495_0[0]));    relay_conn far_7_7495_0_b(.in(layer_6[100]), .out(far_7_7495_0[1]));
    assign out[355] = ~far_7_7495_0[0]; 
    wire [1:0] far_7_7496_0;    relay_conn far_7_7496_0_a(.in(layer_6[550]), .out(far_7_7496_0[0]));    relay_conn far_7_7496_0_b(.in(layer_6[492]), .out(far_7_7496_0[1]));
    assign out[356] = ~(far_7_7496_0[0] | far_7_7496_0[1]); 
    wire [1:0] far_7_7497_0;    relay_conn far_7_7497_0_a(.in(layer_6[393]), .out(far_7_7497_0[0]));    relay_conn far_7_7497_0_b(.in(layer_6[453]), .out(far_7_7497_0[1]));
    assign out[357] = far_7_7497_0[1]; 
    assign out[358] = layer_6[48] & layer_6[51]; 
    wire [1:0] far_7_7499_0;    relay_conn far_7_7499_0_a(.in(layer_6[799]), .out(far_7_7499_0[0]));    relay_conn far_7_7499_0_b(.in(layer_6[721]), .out(far_7_7499_0[1]));
    wire [1:0] far_7_7499_1;    relay_conn far_7_7499_1_a(.in(far_7_7499_0[0]), .out(far_7_7499_1[0]));    relay_conn far_7_7499_1_b(.in(far_7_7499_0[1]), .out(far_7_7499_1[1]));
    assign out[359] = far_7_7499_1[1] & ~far_7_7499_1[0]; 
    wire [1:0] far_7_7500_0;    relay_conn far_7_7500_0_a(.in(layer_6[456]), .out(far_7_7500_0[0]));    relay_conn far_7_7500_0_b(.in(layer_6[339]), .out(far_7_7500_0[1]));
    wire [1:0] far_7_7500_1;    relay_conn far_7_7500_1_a(.in(far_7_7500_0[0]), .out(far_7_7500_1[0]));    relay_conn far_7_7500_1_b(.in(far_7_7500_0[1]), .out(far_7_7500_1[1]));
    wire [1:0] far_7_7500_2;    relay_conn far_7_7500_2_a(.in(far_7_7500_1[0]), .out(far_7_7500_2[0]));    relay_conn far_7_7500_2_b(.in(far_7_7500_1[1]), .out(far_7_7500_2[1]));
    assign out[360] = ~far_7_7500_2[1]; 
    assign out[361] = ~layer_6[874] | (layer_6[874] & layer_6[879]); 
    assign out[362] = layer_6[470] & ~layer_6[451]; 
    wire [1:0] far_7_7503_0;    relay_conn far_7_7503_0_a(.in(layer_6[387]), .out(far_7_7503_0[0]));    relay_conn far_7_7503_0_b(.in(layer_6[500]), .out(far_7_7503_0[1]));
    wire [1:0] far_7_7503_1;    relay_conn far_7_7503_1_a(.in(far_7_7503_0[0]), .out(far_7_7503_1[0]));    relay_conn far_7_7503_1_b(.in(far_7_7503_0[1]), .out(far_7_7503_1[1]));
    wire [1:0] far_7_7503_2;    relay_conn far_7_7503_2_a(.in(far_7_7503_1[0]), .out(far_7_7503_2[0]));    relay_conn far_7_7503_2_b(.in(far_7_7503_1[1]), .out(far_7_7503_2[1]));
    assign out[363] = far_7_7503_2[1]; 
    wire [1:0] far_7_7504_0;    relay_conn far_7_7504_0_a(.in(layer_6[456]), .out(far_7_7504_0[0]));    relay_conn far_7_7504_0_b(.in(layer_6[386]), .out(far_7_7504_0[1]));
    wire [1:0] far_7_7504_1;    relay_conn far_7_7504_1_a(.in(far_7_7504_0[0]), .out(far_7_7504_1[0]));    relay_conn far_7_7504_1_b(.in(far_7_7504_0[1]), .out(far_7_7504_1[1]));
    assign out[364] = ~far_7_7504_1[1]; 
    wire [1:0] far_7_7505_0;    relay_conn far_7_7505_0_a(.in(layer_6[387]), .out(far_7_7505_0[0]));    relay_conn far_7_7505_0_b(.in(layer_6[478]), .out(far_7_7505_0[1]));
    wire [1:0] far_7_7505_1;    relay_conn far_7_7505_1_a(.in(far_7_7505_0[0]), .out(far_7_7505_1[0]));    relay_conn far_7_7505_1_b(.in(far_7_7505_0[1]), .out(far_7_7505_1[1]));
    assign out[365] = ~far_7_7505_1[1]; 
    wire [1:0] far_7_7506_0;    relay_conn far_7_7506_0_a(.in(layer_6[194]), .out(far_7_7506_0[0]));    relay_conn far_7_7506_0_b(.in(layer_6[270]), .out(far_7_7506_0[1]));
    wire [1:0] far_7_7506_1;    relay_conn far_7_7506_1_a(.in(far_7_7506_0[0]), .out(far_7_7506_1[0]));    relay_conn far_7_7506_1_b(.in(far_7_7506_0[1]), .out(far_7_7506_1[1]));
    assign out[366] = far_7_7506_1[0]; 
    wire [1:0] far_7_7507_0;    relay_conn far_7_7507_0_a(.in(layer_6[473]), .out(far_7_7507_0[0]));    relay_conn far_7_7507_0_b(.in(layer_6[345]), .out(far_7_7507_0[1]));
    wire [1:0] far_7_7507_1;    relay_conn far_7_7507_1_a(.in(far_7_7507_0[0]), .out(far_7_7507_1[0]));    relay_conn far_7_7507_1_b(.in(far_7_7507_0[1]), .out(far_7_7507_1[1]));
    wire [1:0] far_7_7507_2;    relay_conn far_7_7507_2_a(.in(far_7_7507_1[0]), .out(far_7_7507_2[0]));    relay_conn far_7_7507_2_b(.in(far_7_7507_1[1]), .out(far_7_7507_2[1]));
    wire [1:0] far_7_7507_3;    relay_conn far_7_7507_3_a(.in(far_7_7507_2[0]), .out(far_7_7507_3[0]));    relay_conn far_7_7507_3_b(.in(far_7_7507_2[1]), .out(far_7_7507_3[1]));
    assign out[367] = ~far_7_7507_3[0]; 
    wire [1:0] far_7_7508_0;    relay_conn far_7_7508_0_a(.in(layer_6[802]), .out(far_7_7508_0[0]));    relay_conn far_7_7508_0_b(.in(layer_6[923]), .out(far_7_7508_0[1]));
    wire [1:0] far_7_7508_1;    relay_conn far_7_7508_1_a(.in(far_7_7508_0[0]), .out(far_7_7508_1[0]));    relay_conn far_7_7508_1_b(.in(far_7_7508_0[1]), .out(far_7_7508_1[1]));
    wire [1:0] far_7_7508_2;    relay_conn far_7_7508_2_a(.in(far_7_7508_1[0]), .out(far_7_7508_2[0]));    relay_conn far_7_7508_2_b(.in(far_7_7508_1[1]), .out(far_7_7508_2[1]));
    assign out[368] = far_7_7508_2[0] ^ far_7_7508_2[1]; 
    wire [1:0] far_7_7509_0;    relay_conn far_7_7509_0_a(.in(layer_6[24]), .out(far_7_7509_0[0]));    relay_conn far_7_7509_0_b(.in(layer_6[113]), .out(far_7_7509_0[1]));
    wire [1:0] far_7_7509_1;    relay_conn far_7_7509_1_a(.in(far_7_7509_0[0]), .out(far_7_7509_1[0]));    relay_conn far_7_7509_1_b(.in(far_7_7509_0[1]), .out(far_7_7509_1[1]));
    assign out[369] = far_7_7509_1[0] & ~far_7_7509_1[1]; 
    assign out[370] = layer_6[763] & ~layer_6[792]; 
    assign out[371] = ~layer_6[53]; 
    wire [1:0] far_7_7512_0;    relay_conn far_7_7512_0_a(.in(layer_6[976]), .out(far_7_7512_0[0]));    relay_conn far_7_7512_0_b(.in(layer_6[929]), .out(far_7_7512_0[1]));
    assign out[372] = ~far_7_7512_0[1]; 
    wire [1:0] far_7_7513_0;    relay_conn far_7_7513_0_a(.in(layer_6[821]), .out(far_7_7513_0[0]));    relay_conn far_7_7513_0_b(.in(layer_6[917]), .out(far_7_7513_0[1]));
    wire [1:0] far_7_7513_1;    relay_conn far_7_7513_1_a(.in(far_7_7513_0[0]), .out(far_7_7513_1[0]));    relay_conn far_7_7513_1_b(.in(far_7_7513_0[1]), .out(far_7_7513_1[1]));
    wire [1:0] far_7_7513_2;    relay_conn far_7_7513_2_a(.in(far_7_7513_1[0]), .out(far_7_7513_2[0]));    relay_conn far_7_7513_2_b(.in(far_7_7513_1[1]), .out(far_7_7513_2[1]));
    assign out[373] = far_7_7513_2[0]; 
    wire [1:0] far_7_7514_0;    relay_conn far_7_7514_0_a(.in(layer_6[1018]), .out(far_7_7514_0[0]));    relay_conn far_7_7514_0_b(.in(layer_6[951]), .out(far_7_7514_0[1]));
    wire [1:0] far_7_7514_1;    relay_conn far_7_7514_1_a(.in(far_7_7514_0[0]), .out(far_7_7514_1[0]));    relay_conn far_7_7514_1_b(.in(far_7_7514_0[1]), .out(far_7_7514_1[1]));
    assign out[374] = far_7_7514_1[1]; 
    assign out[375] = layer_6[591] & ~layer_6[601]; 
    wire [1:0] far_7_7516_0;    relay_conn far_7_7516_0_a(.in(layer_6[285]), .out(far_7_7516_0[0]));    relay_conn far_7_7516_0_b(.in(layer_6[404]), .out(far_7_7516_0[1]));
    wire [1:0] far_7_7516_1;    relay_conn far_7_7516_1_a(.in(far_7_7516_0[0]), .out(far_7_7516_1[0]));    relay_conn far_7_7516_1_b(.in(far_7_7516_0[1]), .out(far_7_7516_1[1]));
    wire [1:0] far_7_7516_2;    relay_conn far_7_7516_2_a(.in(far_7_7516_1[0]), .out(far_7_7516_2[0]));    relay_conn far_7_7516_2_b(.in(far_7_7516_1[1]), .out(far_7_7516_2[1]));
    assign out[376] = ~far_7_7516_2[1]; 
    wire [1:0] far_7_7517_0;    relay_conn far_7_7517_0_a(.in(layer_6[250]), .out(far_7_7517_0[0]));    relay_conn far_7_7517_0_b(.in(layer_6[333]), .out(far_7_7517_0[1]));
    wire [1:0] far_7_7517_1;    relay_conn far_7_7517_1_a(.in(far_7_7517_0[0]), .out(far_7_7517_1[0]));    relay_conn far_7_7517_1_b(.in(far_7_7517_0[1]), .out(far_7_7517_1[1]));
    assign out[377] = ~(far_7_7517_1[0] ^ far_7_7517_1[1]); 
    wire [1:0] far_7_7518_0;    relay_conn far_7_7518_0_a(.in(layer_6[230]), .out(far_7_7518_0[0]));    relay_conn far_7_7518_0_b(.in(layer_6[286]), .out(far_7_7518_0[1]));
    assign out[378] = ~far_7_7518_0[0]; 
    wire [1:0] far_7_7519_0;    relay_conn far_7_7519_0_a(.in(layer_6[834]), .out(far_7_7519_0[0]));    relay_conn far_7_7519_0_b(.in(layer_6[924]), .out(far_7_7519_0[1]));
    wire [1:0] far_7_7519_1;    relay_conn far_7_7519_1_a(.in(far_7_7519_0[0]), .out(far_7_7519_1[0]));    relay_conn far_7_7519_1_b(.in(far_7_7519_0[1]), .out(far_7_7519_1[1]));
    assign out[379] = ~far_7_7519_1[1]; 
    wire [1:0] far_7_7520_0;    relay_conn far_7_7520_0_a(.in(layer_6[323]), .out(far_7_7520_0[0]));    relay_conn far_7_7520_0_b(.in(layer_6[416]), .out(far_7_7520_0[1]));
    wire [1:0] far_7_7520_1;    relay_conn far_7_7520_1_a(.in(far_7_7520_0[0]), .out(far_7_7520_1[0]));    relay_conn far_7_7520_1_b(.in(far_7_7520_0[1]), .out(far_7_7520_1[1]));
    assign out[380] = far_7_7520_1[0] & ~far_7_7520_1[1]; 
    wire [1:0] far_7_7521_0;    relay_conn far_7_7521_0_a(.in(layer_6[550]), .out(far_7_7521_0[0]));    relay_conn far_7_7521_0_b(.in(layer_6[676]), .out(far_7_7521_0[1]));
    wire [1:0] far_7_7521_1;    relay_conn far_7_7521_1_a(.in(far_7_7521_0[0]), .out(far_7_7521_1[0]));    relay_conn far_7_7521_1_b(.in(far_7_7521_0[1]), .out(far_7_7521_1[1]));
    wire [1:0] far_7_7521_2;    relay_conn far_7_7521_2_a(.in(far_7_7521_1[0]), .out(far_7_7521_2[0]));    relay_conn far_7_7521_2_b(.in(far_7_7521_1[1]), .out(far_7_7521_2[1]));
    assign out[381] = ~(far_7_7521_2[0] | far_7_7521_2[1]); 
    wire [1:0] far_7_7522_0;    relay_conn far_7_7522_0_a(.in(layer_6[403]), .out(far_7_7522_0[0]));    relay_conn far_7_7522_0_b(.in(layer_6[342]), .out(far_7_7522_0[1]));
    assign out[382] = ~far_7_7522_0[0]; 
    wire [1:0] far_7_7523_0;    relay_conn far_7_7523_0_a(.in(layer_6[736]), .out(far_7_7523_0[0]));    relay_conn far_7_7523_0_b(.in(layer_6[642]), .out(far_7_7523_0[1]));
    wire [1:0] far_7_7523_1;    relay_conn far_7_7523_1_a(.in(far_7_7523_0[0]), .out(far_7_7523_1[0]));    relay_conn far_7_7523_1_b(.in(far_7_7523_0[1]), .out(far_7_7523_1[1]));
    assign out[383] = ~far_7_7523_1[0]; 
    wire [1:0] far_7_7524_0;    relay_conn far_7_7524_0_a(.in(layer_6[230]), .out(far_7_7524_0[0]));    relay_conn far_7_7524_0_b(.in(layer_6[190]), .out(far_7_7524_0[1]));
    assign out[384] = ~far_7_7524_0[0] | (far_7_7524_0[0] & far_7_7524_0[1]); 
    wire [1:0] far_7_7525_0;    relay_conn far_7_7525_0_a(.in(layer_6[262]), .out(far_7_7525_0[0]));    relay_conn far_7_7525_0_b(.in(layer_6[157]), .out(far_7_7525_0[1]));
    wire [1:0] far_7_7525_1;    relay_conn far_7_7525_1_a(.in(far_7_7525_0[0]), .out(far_7_7525_1[0]));    relay_conn far_7_7525_1_b(.in(far_7_7525_0[1]), .out(far_7_7525_1[1]));
    wire [1:0] far_7_7525_2;    relay_conn far_7_7525_2_a(.in(far_7_7525_1[0]), .out(far_7_7525_2[0]));    relay_conn far_7_7525_2_b(.in(far_7_7525_1[1]), .out(far_7_7525_2[1]));
    assign out[385] = ~far_7_7525_2[0]; 
    wire [1:0] far_7_7526_0;    relay_conn far_7_7526_0_a(.in(layer_6[315]), .out(far_7_7526_0[0]));    relay_conn far_7_7526_0_b(.in(layer_6[261]), .out(far_7_7526_0[1]));
    assign out[386] = far_7_7526_0[0] & ~far_7_7526_0[1]; 
    wire [1:0] far_7_7527_0;    relay_conn far_7_7527_0_a(.in(layer_6[886]), .out(far_7_7527_0[0]));    relay_conn far_7_7527_0_b(.in(layer_6[760]), .out(far_7_7527_0[1]));
    wire [1:0] far_7_7527_1;    relay_conn far_7_7527_1_a(.in(far_7_7527_0[0]), .out(far_7_7527_1[0]));    relay_conn far_7_7527_1_b(.in(far_7_7527_0[1]), .out(far_7_7527_1[1]));
    wire [1:0] far_7_7527_2;    relay_conn far_7_7527_2_a(.in(far_7_7527_1[0]), .out(far_7_7527_2[0]));    relay_conn far_7_7527_2_b(.in(far_7_7527_1[1]), .out(far_7_7527_2[1]));
    assign out[387] = far_7_7527_2[0] ^ far_7_7527_2[1]; 
    wire [1:0] far_7_7528_0;    relay_conn far_7_7528_0_a(.in(layer_6[315]), .out(far_7_7528_0[0]));    relay_conn far_7_7528_0_b(.in(layer_6[388]), .out(far_7_7528_0[1]));
    wire [1:0] far_7_7528_1;    relay_conn far_7_7528_1_a(.in(far_7_7528_0[0]), .out(far_7_7528_1[0]));    relay_conn far_7_7528_1_b(.in(far_7_7528_0[1]), .out(far_7_7528_1[1]));
    assign out[388] = ~(far_7_7528_1[0] ^ far_7_7528_1[1]); 
    wire [1:0] far_7_7529_0;    relay_conn far_7_7529_0_a(.in(layer_6[733]), .out(far_7_7529_0[0]));    relay_conn far_7_7529_0_b(.in(layer_6[847]), .out(far_7_7529_0[1]));
    wire [1:0] far_7_7529_1;    relay_conn far_7_7529_1_a(.in(far_7_7529_0[0]), .out(far_7_7529_1[0]));    relay_conn far_7_7529_1_b(.in(far_7_7529_0[1]), .out(far_7_7529_1[1]));
    wire [1:0] far_7_7529_2;    relay_conn far_7_7529_2_a(.in(far_7_7529_1[0]), .out(far_7_7529_2[0]));    relay_conn far_7_7529_2_b(.in(far_7_7529_1[1]), .out(far_7_7529_2[1]));
    assign out[389] = ~far_7_7529_2[1] | (far_7_7529_2[0] & far_7_7529_2[1]); 
    wire [1:0] far_7_7530_0;    relay_conn far_7_7530_0_a(.in(layer_6[681]), .out(far_7_7530_0[0]));    relay_conn far_7_7530_0_b(.in(layer_6[600]), .out(far_7_7530_0[1]));
    wire [1:0] far_7_7530_1;    relay_conn far_7_7530_1_a(.in(far_7_7530_0[0]), .out(far_7_7530_1[0]));    relay_conn far_7_7530_1_b(.in(far_7_7530_0[1]), .out(far_7_7530_1[1]));
    assign out[390] = ~far_7_7530_1[1]; 
    wire [1:0] far_7_7531_0;    relay_conn far_7_7531_0_a(.in(layer_6[711]), .out(far_7_7531_0[0]));    relay_conn far_7_7531_0_b(.in(layer_6[766]), .out(far_7_7531_0[1]));
    assign out[391] = far_7_7531_0[0] & far_7_7531_0[1]; 
    wire [1:0] far_7_7532_0;    relay_conn far_7_7532_0_a(.in(layer_6[825]), .out(far_7_7532_0[0]));    relay_conn far_7_7532_0_b(.in(layer_6[777]), .out(far_7_7532_0[1]));
    assign out[392] = ~far_7_7532_0[0]; 
    assign out[393] = layer_6[675] & ~layer_6[650]; 
    wire [1:0] far_7_7534_0;    relay_conn far_7_7534_0_a(.in(layer_6[766]), .out(far_7_7534_0[0]));    relay_conn far_7_7534_0_b(.in(layer_6[659]), .out(far_7_7534_0[1]));
    wire [1:0] far_7_7534_1;    relay_conn far_7_7534_1_a(.in(far_7_7534_0[0]), .out(far_7_7534_1[0]));    relay_conn far_7_7534_1_b(.in(far_7_7534_0[1]), .out(far_7_7534_1[1]));
    wire [1:0] far_7_7534_2;    relay_conn far_7_7534_2_a(.in(far_7_7534_1[0]), .out(far_7_7534_2[0]));    relay_conn far_7_7534_2_b(.in(far_7_7534_1[1]), .out(far_7_7534_2[1]));
    assign out[394] = far_7_7534_2[0] & ~far_7_7534_2[1]; 
    wire [1:0] far_7_7535_0;    relay_conn far_7_7535_0_a(.in(layer_6[159]), .out(far_7_7535_0[0]));    relay_conn far_7_7535_0_b(.in(layer_6[210]), .out(far_7_7535_0[1]));
    assign out[395] = ~(far_7_7535_0[0] | far_7_7535_0[1]); 
    wire [1:0] far_7_7536_0;    relay_conn far_7_7536_0_a(.in(layer_6[632]), .out(far_7_7536_0[0]));    relay_conn far_7_7536_0_b(.in(layer_6[587]), .out(far_7_7536_0[1]));
    assign out[396] = far_7_7536_0[1]; 
    assign out[397] = layer_6[194] & layer_6[215]; 
    assign out[398] = ~layer_6[416]; 
    wire [1:0] far_7_7539_0;    relay_conn far_7_7539_0_a(.in(layer_6[322]), .out(far_7_7539_0[0]));    relay_conn far_7_7539_0_b(.in(layer_6[424]), .out(far_7_7539_0[1]));
    wire [1:0] far_7_7539_1;    relay_conn far_7_7539_1_a(.in(far_7_7539_0[0]), .out(far_7_7539_1[0]));    relay_conn far_7_7539_1_b(.in(far_7_7539_0[1]), .out(far_7_7539_1[1]));
    wire [1:0] far_7_7539_2;    relay_conn far_7_7539_2_a(.in(far_7_7539_1[0]), .out(far_7_7539_2[0]));    relay_conn far_7_7539_2_b(.in(far_7_7539_1[1]), .out(far_7_7539_2[1]));
    assign out[399] = far_7_7539_2[0]; 
    wire [1:0] far_7_7540_0;    relay_conn far_7_7540_0_a(.in(layer_6[109]), .out(far_7_7540_0[0]));    relay_conn far_7_7540_0_b(.in(layer_6[198]), .out(far_7_7540_0[1]));
    wire [1:0] far_7_7540_1;    relay_conn far_7_7540_1_a(.in(far_7_7540_0[0]), .out(far_7_7540_1[0]));    relay_conn far_7_7540_1_b(.in(far_7_7540_0[1]), .out(far_7_7540_1[1]));
    assign out[400] = far_7_7540_1[1] & ~far_7_7540_1[0]; 
    assign out[401] = ~(layer_6[786] ^ layer_6[815]); 
    assign out[402] = layer_6[614]; 
    wire [1:0] far_7_7543_0;    relay_conn far_7_7543_0_a(.in(layer_6[632]), .out(far_7_7543_0[0]));    relay_conn far_7_7543_0_b(.in(layer_6[558]), .out(far_7_7543_0[1]));
    wire [1:0] far_7_7543_1;    relay_conn far_7_7543_1_a(.in(far_7_7543_0[0]), .out(far_7_7543_1[0]));    relay_conn far_7_7543_1_b(.in(far_7_7543_0[1]), .out(far_7_7543_1[1]));
    assign out[403] = far_7_7543_1[0] & far_7_7543_1[1]; 
    wire [1:0] far_7_7544_0;    relay_conn far_7_7544_0_a(.in(layer_6[995]), .out(far_7_7544_0[0]));    relay_conn far_7_7544_0_b(.in(layer_6[910]), .out(far_7_7544_0[1]));
    wire [1:0] far_7_7544_1;    relay_conn far_7_7544_1_a(.in(far_7_7544_0[0]), .out(far_7_7544_1[0]));    relay_conn far_7_7544_1_b(.in(far_7_7544_0[1]), .out(far_7_7544_1[1]));
    assign out[404] = ~(far_7_7544_1[0] | far_7_7544_1[1]); 
    wire [1:0] far_7_7545_0;    relay_conn far_7_7545_0_a(.in(layer_6[577]), .out(far_7_7545_0[0]));    relay_conn far_7_7545_0_b(.in(layer_6[646]), .out(far_7_7545_0[1]));
    wire [1:0] far_7_7545_1;    relay_conn far_7_7545_1_a(.in(far_7_7545_0[0]), .out(far_7_7545_1[0]));    relay_conn far_7_7545_1_b(.in(far_7_7545_0[1]), .out(far_7_7545_1[1]));
    assign out[405] = far_7_7545_1[0] & far_7_7545_1[1]; 
    wire [1:0] far_7_7546_0;    relay_conn far_7_7546_0_a(.in(layer_6[683]), .out(far_7_7546_0[0]));    relay_conn far_7_7546_0_b(.in(layer_6[577]), .out(far_7_7546_0[1]));
    wire [1:0] far_7_7546_1;    relay_conn far_7_7546_1_a(.in(far_7_7546_0[0]), .out(far_7_7546_1[0]));    relay_conn far_7_7546_1_b(.in(far_7_7546_0[1]), .out(far_7_7546_1[1]));
    wire [1:0] far_7_7546_2;    relay_conn far_7_7546_2_a(.in(far_7_7546_1[0]), .out(far_7_7546_2[0]));    relay_conn far_7_7546_2_b(.in(far_7_7546_1[1]), .out(far_7_7546_2[1]));
    assign out[406] = far_7_7546_2[1]; 
    wire [1:0] far_7_7547_0;    relay_conn far_7_7547_0_a(.in(layer_6[277]), .out(far_7_7547_0[0]));    relay_conn far_7_7547_0_b(.in(layer_6[176]), .out(far_7_7547_0[1]));
    wire [1:0] far_7_7547_1;    relay_conn far_7_7547_1_a(.in(far_7_7547_0[0]), .out(far_7_7547_1[0]));    relay_conn far_7_7547_1_b(.in(far_7_7547_0[1]), .out(far_7_7547_1[1]));
    wire [1:0] far_7_7547_2;    relay_conn far_7_7547_2_a(.in(far_7_7547_1[0]), .out(far_7_7547_2[0]));    relay_conn far_7_7547_2_b(.in(far_7_7547_1[1]), .out(far_7_7547_2[1]));
    assign out[407] = far_7_7547_2[0] & far_7_7547_2[1]; 
    wire [1:0] far_7_7548_0;    relay_conn far_7_7548_0_a(.in(layer_6[650]), .out(far_7_7548_0[0]));    relay_conn far_7_7548_0_b(.in(layer_6[607]), .out(far_7_7548_0[1]));
    assign out[408] = far_7_7548_0[0]; 
    wire [1:0] far_7_7549_0;    relay_conn far_7_7549_0_a(.in(layer_6[575]), .out(far_7_7549_0[0]));    relay_conn far_7_7549_0_b(.in(layer_6[469]), .out(far_7_7549_0[1]));
    wire [1:0] far_7_7549_1;    relay_conn far_7_7549_1_a(.in(far_7_7549_0[0]), .out(far_7_7549_1[0]));    relay_conn far_7_7549_1_b(.in(far_7_7549_0[1]), .out(far_7_7549_1[1]));
    wire [1:0] far_7_7549_2;    relay_conn far_7_7549_2_a(.in(far_7_7549_1[0]), .out(far_7_7549_2[0]));    relay_conn far_7_7549_2_b(.in(far_7_7549_1[1]), .out(far_7_7549_2[1]));
    assign out[409] = far_7_7549_2[0] & ~far_7_7549_2[1]; 
    wire [1:0] far_7_7550_0;    relay_conn far_7_7550_0_a(.in(layer_6[908]), .out(far_7_7550_0[0]));    relay_conn far_7_7550_0_b(.in(layer_6[873]), .out(far_7_7550_0[1]));
    assign out[410] = ~(far_7_7550_0[0] ^ far_7_7550_0[1]); 
    wire [1:0] far_7_7551_0;    relay_conn far_7_7551_0_a(.in(layer_6[57]), .out(far_7_7551_0[0]));    relay_conn far_7_7551_0_b(.in(layer_6[151]), .out(far_7_7551_0[1]));
    wire [1:0] far_7_7551_1;    relay_conn far_7_7551_1_a(.in(far_7_7551_0[0]), .out(far_7_7551_1[0]));    relay_conn far_7_7551_1_b(.in(far_7_7551_0[1]), .out(far_7_7551_1[1]));
    assign out[411] = ~(far_7_7551_1[0] | far_7_7551_1[1]); 
    wire [1:0] far_7_7552_0;    relay_conn far_7_7552_0_a(.in(layer_6[424]), .out(far_7_7552_0[0]));    relay_conn far_7_7552_0_b(.in(layer_6[531]), .out(far_7_7552_0[1]));
    wire [1:0] far_7_7552_1;    relay_conn far_7_7552_1_a(.in(far_7_7552_0[0]), .out(far_7_7552_1[0]));    relay_conn far_7_7552_1_b(.in(far_7_7552_0[1]), .out(far_7_7552_1[1]));
    wire [1:0] far_7_7552_2;    relay_conn far_7_7552_2_a(.in(far_7_7552_1[0]), .out(far_7_7552_2[0]));    relay_conn far_7_7552_2_b(.in(far_7_7552_1[1]), .out(far_7_7552_2[1]));
    assign out[412] = far_7_7552_2[1]; 
    wire [1:0] far_7_7553_0;    relay_conn far_7_7553_0_a(.in(layer_6[142]), .out(far_7_7553_0[0]));    relay_conn far_7_7553_0_b(.in(layer_6[100]), .out(far_7_7553_0[1]));
    assign out[413] = ~(far_7_7553_0[0] | far_7_7553_0[1]); 
    assign out[414] = ~(layer_6[777] | layer_6[762]); 
    wire [1:0] far_7_7555_0;    relay_conn far_7_7555_0_a(.in(layer_6[317]), .out(far_7_7555_0[0]));    relay_conn far_7_7555_0_b(.in(layer_6[425]), .out(far_7_7555_0[1]));
    wire [1:0] far_7_7555_1;    relay_conn far_7_7555_1_a(.in(far_7_7555_0[0]), .out(far_7_7555_1[0]));    relay_conn far_7_7555_1_b(.in(far_7_7555_0[1]), .out(far_7_7555_1[1]));
    wire [1:0] far_7_7555_2;    relay_conn far_7_7555_2_a(.in(far_7_7555_1[0]), .out(far_7_7555_2[0]));    relay_conn far_7_7555_2_b(.in(far_7_7555_1[1]), .out(far_7_7555_2[1]));
    assign out[415] = ~far_7_7555_2[0]; 
    wire [1:0] far_7_7556_0;    relay_conn far_7_7556_0_a(.in(layer_6[794]), .out(far_7_7556_0[0]));    relay_conn far_7_7556_0_b(.in(layer_6[687]), .out(far_7_7556_0[1]));
    wire [1:0] far_7_7556_1;    relay_conn far_7_7556_1_a(.in(far_7_7556_0[0]), .out(far_7_7556_1[0]));    relay_conn far_7_7556_1_b(.in(far_7_7556_0[1]), .out(far_7_7556_1[1]));
    wire [1:0] far_7_7556_2;    relay_conn far_7_7556_2_a(.in(far_7_7556_1[0]), .out(far_7_7556_2[0]));    relay_conn far_7_7556_2_b(.in(far_7_7556_1[1]), .out(far_7_7556_2[1]));
    assign out[416] = far_7_7556_2[0] & far_7_7556_2[1]; 
    wire [1:0] far_7_7557_0;    relay_conn far_7_7557_0_a(.in(layer_6[117]), .out(far_7_7557_0[0]));    relay_conn far_7_7557_0_b(.in(layer_6[226]), .out(far_7_7557_0[1]));
    wire [1:0] far_7_7557_1;    relay_conn far_7_7557_1_a(.in(far_7_7557_0[0]), .out(far_7_7557_1[0]));    relay_conn far_7_7557_1_b(.in(far_7_7557_0[1]), .out(far_7_7557_1[1]));
    wire [1:0] far_7_7557_2;    relay_conn far_7_7557_2_a(.in(far_7_7557_1[0]), .out(far_7_7557_2[0]));    relay_conn far_7_7557_2_b(.in(far_7_7557_1[1]), .out(far_7_7557_2[1]));
    assign out[417] = far_7_7557_2[1] & ~far_7_7557_2[0]; 
    wire [1:0] far_7_7558_0;    relay_conn far_7_7558_0_a(.in(layer_6[312]), .out(far_7_7558_0[0]));    relay_conn far_7_7558_0_b(.in(layer_6[210]), .out(far_7_7558_0[1]));
    wire [1:0] far_7_7558_1;    relay_conn far_7_7558_1_a(.in(far_7_7558_0[0]), .out(far_7_7558_1[0]));    relay_conn far_7_7558_1_b(.in(far_7_7558_0[1]), .out(far_7_7558_1[1]));
    wire [1:0] far_7_7558_2;    relay_conn far_7_7558_2_a(.in(far_7_7558_1[0]), .out(far_7_7558_2[0]));    relay_conn far_7_7558_2_b(.in(far_7_7558_1[1]), .out(far_7_7558_2[1]));
    assign out[418] = far_7_7558_2[1] & ~far_7_7558_2[0]; 
    wire [1:0] far_7_7559_0;    relay_conn far_7_7559_0_a(.in(layer_6[550]), .out(far_7_7559_0[0]));    relay_conn far_7_7559_0_b(.in(layer_6[483]), .out(far_7_7559_0[1]));
    wire [1:0] far_7_7559_1;    relay_conn far_7_7559_1_a(.in(far_7_7559_0[0]), .out(far_7_7559_1[0]));    relay_conn far_7_7559_1_b(.in(far_7_7559_0[1]), .out(far_7_7559_1[1]));
    assign out[419] = far_7_7559_1[1] & ~far_7_7559_1[0]; 
    wire [1:0] far_7_7560_0;    relay_conn far_7_7560_0_a(.in(layer_6[57]), .out(far_7_7560_0[0]));    relay_conn far_7_7560_0_b(.in(layer_6[140]), .out(far_7_7560_0[1]));
    wire [1:0] far_7_7560_1;    relay_conn far_7_7560_1_a(.in(far_7_7560_0[0]), .out(far_7_7560_1[0]));    relay_conn far_7_7560_1_b(.in(far_7_7560_0[1]), .out(far_7_7560_1[1]));
    assign out[420] = far_7_7560_1[1] & ~far_7_7560_1[0]; 
    wire [1:0] far_7_7561_0;    relay_conn far_7_7561_0_a(.in(layer_6[443]), .out(far_7_7561_0[0]));    relay_conn far_7_7561_0_b(.in(layer_6[384]), .out(far_7_7561_0[1]));
    assign out[421] = ~(far_7_7561_0[0] | far_7_7561_0[1]); 
    wire [1:0] far_7_7562_0;    relay_conn far_7_7562_0_a(.in(layer_6[203]), .out(far_7_7562_0[0]));    relay_conn far_7_7562_0_b(.in(layer_6[100]), .out(far_7_7562_0[1]));
    wire [1:0] far_7_7562_1;    relay_conn far_7_7562_1_a(.in(far_7_7562_0[0]), .out(far_7_7562_1[0]));    relay_conn far_7_7562_1_b(.in(far_7_7562_0[1]), .out(far_7_7562_1[1]));
    wire [1:0] far_7_7562_2;    relay_conn far_7_7562_2_a(.in(far_7_7562_1[0]), .out(far_7_7562_2[0]));    relay_conn far_7_7562_2_b(.in(far_7_7562_1[1]), .out(far_7_7562_2[1]));
    assign out[422] = ~(far_7_7562_2[0] | far_7_7562_2[1]); 
    wire [1:0] far_7_7563_0;    relay_conn far_7_7563_0_a(.in(layer_6[716]), .out(far_7_7563_0[0]));    relay_conn far_7_7563_0_b(.in(layer_6[629]), .out(far_7_7563_0[1]));
    wire [1:0] far_7_7563_1;    relay_conn far_7_7563_1_a(.in(far_7_7563_0[0]), .out(far_7_7563_1[0]));    relay_conn far_7_7563_1_b(.in(far_7_7563_0[1]), .out(far_7_7563_1[1]));
    assign out[423] = ~(far_7_7563_1[0] ^ far_7_7563_1[1]); 
    wire [1:0] far_7_7564_0;    relay_conn far_7_7564_0_a(.in(layer_6[117]), .out(far_7_7564_0[0]));    relay_conn far_7_7564_0_b(.in(layer_6[48]), .out(far_7_7564_0[1]));
    wire [1:0] far_7_7564_1;    relay_conn far_7_7564_1_a(.in(far_7_7564_0[0]), .out(far_7_7564_1[0]));    relay_conn far_7_7564_1_b(.in(far_7_7564_0[1]), .out(far_7_7564_1[1]));
    assign out[424] = ~(far_7_7564_1[0] | far_7_7564_1[1]); 
    assign out[425] = layer_6[569]; 
    wire [1:0] far_7_7566_0;    relay_conn far_7_7566_0_a(.in(layer_6[765]), .out(far_7_7566_0[0]));    relay_conn far_7_7566_0_b(.in(layer_6[663]), .out(far_7_7566_0[1]));
    wire [1:0] far_7_7566_1;    relay_conn far_7_7566_1_a(.in(far_7_7566_0[0]), .out(far_7_7566_1[0]));    relay_conn far_7_7566_1_b(.in(far_7_7566_0[1]), .out(far_7_7566_1[1]));
    wire [1:0] far_7_7566_2;    relay_conn far_7_7566_2_a(.in(far_7_7566_1[0]), .out(far_7_7566_2[0]));    relay_conn far_7_7566_2_b(.in(far_7_7566_1[1]), .out(far_7_7566_2[1]));
    assign out[426] = ~(far_7_7566_2[0] ^ far_7_7566_2[1]); 
    assign out[427] = layer_6[261]; 
    assign out[428] = ~(layer_6[583] | layer_6[611]); 
    wire [1:0] far_7_7569_0;    relay_conn far_7_7569_0_a(.in(layer_6[908]), .out(far_7_7569_0[0]));    relay_conn far_7_7569_0_b(.in(layer_6[821]), .out(far_7_7569_0[1]));
    wire [1:0] far_7_7569_1;    relay_conn far_7_7569_1_a(.in(far_7_7569_0[0]), .out(far_7_7569_1[0]));    relay_conn far_7_7569_1_b(.in(far_7_7569_0[1]), .out(far_7_7569_1[1]));
    assign out[429] = far_7_7569_1[0] ^ far_7_7569_1[1]; 
    wire [1:0] far_7_7570_0;    relay_conn far_7_7570_0_a(.in(layer_6[336]), .out(far_7_7570_0[0]));    relay_conn far_7_7570_0_b(.in(layer_6[268]), .out(far_7_7570_0[1]));
    wire [1:0] far_7_7570_1;    relay_conn far_7_7570_1_a(.in(far_7_7570_0[0]), .out(far_7_7570_1[0]));    relay_conn far_7_7570_1_b(.in(far_7_7570_0[1]), .out(far_7_7570_1[1]));
    assign out[430] = far_7_7570_1[0] & far_7_7570_1[1]; 
    wire [1:0] far_7_7571_0;    relay_conn far_7_7571_0_a(.in(layer_6[76]), .out(far_7_7571_0[0]));    relay_conn far_7_7571_0_b(.in(layer_6[175]), .out(far_7_7571_0[1]));
    wire [1:0] far_7_7571_1;    relay_conn far_7_7571_1_a(.in(far_7_7571_0[0]), .out(far_7_7571_1[0]));    relay_conn far_7_7571_1_b(.in(far_7_7571_0[1]), .out(far_7_7571_1[1]));
    wire [1:0] far_7_7571_2;    relay_conn far_7_7571_2_a(.in(far_7_7571_1[0]), .out(far_7_7571_2[0]));    relay_conn far_7_7571_2_b(.in(far_7_7571_1[1]), .out(far_7_7571_2[1]));
    assign out[431] = ~far_7_7571_2[0]; 
    wire [1:0] far_7_7572_0;    relay_conn far_7_7572_0_a(.in(layer_6[117]), .out(far_7_7572_0[0]));    relay_conn far_7_7572_0_b(.in(layer_6[208]), .out(far_7_7572_0[1]));
    wire [1:0] far_7_7572_1;    relay_conn far_7_7572_1_a(.in(far_7_7572_0[0]), .out(far_7_7572_1[0]));    relay_conn far_7_7572_1_b(.in(far_7_7572_0[1]), .out(far_7_7572_1[1]));
    assign out[432] = ~(far_7_7572_1[0] | far_7_7572_1[1]); 
    wire [1:0] far_7_7573_0;    relay_conn far_7_7573_0_a(.in(layer_6[336]), .out(far_7_7573_0[0]));    relay_conn far_7_7573_0_b(.in(layer_6[257]), .out(far_7_7573_0[1]));
    wire [1:0] far_7_7573_1;    relay_conn far_7_7573_1_a(.in(far_7_7573_0[0]), .out(far_7_7573_1[0]));    relay_conn far_7_7573_1_b(.in(far_7_7573_0[1]), .out(far_7_7573_1[1]));
    assign out[433] = far_7_7573_1[0] & far_7_7573_1[1]; 
    wire [1:0] far_7_7574_0;    relay_conn far_7_7574_0_a(.in(layer_6[434]), .out(far_7_7574_0[0]));    relay_conn far_7_7574_0_b(.in(layer_6[387]), .out(far_7_7574_0[1]));
    assign out[434] = ~far_7_7574_0[0]; 
    assign out[435] = ~(layer_6[923] | layer_6[910]); 
    wire [1:0] far_7_7576_0;    relay_conn far_7_7576_0_a(.in(layer_6[995]), .out(far_7_7576_0[0]));    relay_conn far_7_7576_0_b(.in(layer_6[892]), .out(far_7_7576_0[1]));
    wire [1:0] far_7_7576_1;    relay_conn far_7_7576_1_a(.in(far_7_7576_0[0]), .out(far_7_7576_1[0]));    relay_conn far_7_7576_1_b(.in(far_7_7576_0[1]), .out(far_7_7576_1[1]));
    wire [1:0] far_7_7576_2;    relay_conn far_7_7576_2_a(.in(far_7_7576_1[0]), .out(far_7_7576_2[0]));    relay_conn far_7_7576_2_b(.in(far_7_7576_1[1]), .out(far_7_7576_2[1]));
    assign out[436] = ~far_7_7576_2[1]; 
    wire [1:0] far_7_7577_0;    relay_conn far_7_7577_0_a(.in(layer_6[257]), .out(far_7_7577_0[0]));    relay_conn far_7_7577_0_b(.in(layer_6[177]), .out(far_7_7577_0[1]));
    wire [1:0] far_7_7577_1;    relay_conn far_7_7577_1_a(.in(far_7_7577_0[0]), .out(far_7_7577_1[0]));    relay_conn far_7_7577_1_b(.in(far_7_7577_0[1]), .out(far_7_7577_1[1]));
    assign out[437] = far_7_7577_1[0] & ~far_7_7577_1[1]; 
    assign out[438] = ~layer_6[898]; 
    wire [1:0] far_7_7579_0;    relay_conn far_7_7579_0_a(.in(layer_6[919]), .out(far_7_7579_0[0]));    relay_conn far_7_7579_0_b(.in(layer_6[952]), .out(far_7_7579_0[1]));
    assign out[439] = far_7_7579_0[0] & ~far_7_7579_0[1]; 
    wire [1:0] far_7_7580_0;    relay_conn far_7_7580_0_a(.in(layer_6[802]), .out(far_7_7580_0[0]));    relay_conn far_7_7580_0_b(.in(layer_6[895]), .out(far_7_7580_0[1]));
    wire [1:0] far_7_7580_1;    relay_conn far_7_7580_1_a(.in(far_7_7580_0[0]), .out(far_7_7580_1[0]));    relay_conn far_7_7580_1_b(.in(far_7_7580_0[1]), .out(far_7_7580_1[1]));
    assign out[440] = ~(far_7_7580_1[0] | far_7_7580_1[1]); 
    wire [1:0] far_7_7581_0;    relay_conn far_7_7581_0_a(.in(layer_6[260]), .out(far_7_7581_0[0]));    relay_conn far_7_7581_0_b(.in(layer_6[190]), .out(far_7_7581_0[1]));
    wire [1:0] far_7_7581_1;    relay_conn far_7_7581_1_a(.in(far_7_7581_0[0]), .out(far_7_7581_1[0]));    relay_conn far_7_7581_1_b(.in(far_7_7581_0[1]), .out(far_7_7581_1[1]));
    assign out[441] = ~(far_7_7581_1[0] | far_7_7581_1[1]); 
    wire [1:0] far_7_7582_0;    relay_conn far_7_7582_0_a(.in(layer_6[770]), .out(far_7_7582_0[0]));    relay_conn far_7_7582_0_b(.in(layer_6[718]), .out(far_7_7582_0[1]));
    assign out[442] = ~(far_7_7582_0[0] | far_7_7582_0[1]); 
    wire [1:0] far_7_7583_0;    relay_conn far_7_7583_0_a(.in(layer_6[181]), .out(far_7_7583_0[0]));    relay_conn far_7_7583_0_b(.in(layer_6[57]), .out(far_7_7583_0[1]));
    wire [1:0] far_7_7583_1;    relay_conn far_7_7583_1_a(.in(far_7_7583_0[0]), .out(far_7_7583_1[0]));    relay_conn far_7_7583_1_b(.in(far_7_7583_0[1]), .out(far_7_7583_1[1]));
    wire [1:0] far_7_7583_2;    relay_conn far_7_7583_2_a(.in(far_7_7583_1[0]), .out(far_7_7583_2[0]));    relay_conn far_7_7583_2_b(.in(far_7_7583_1[1]), .out(far_7_7583_2[1]));
    assign out[443] = ~(far_7_7583_2[0] | far_7_7583_2[1]); 
    assign out[444] = layer_6[109] & ~layer_6[100]; 
    wire [1:0] far_7_7585_0;    relay_conn far_7_7585_0_a(.in(layer_6[747]), .out(far_7_7585_0[0]));    relay_conn far_7_7585_0_b(.in(layer_6[663]), .out(far_7_7585_0[1]));
    wire [1:0] far_7_7585_1;    relay_conn far_7_7585_1_a(.in(far_7_7585_0[0]), .out(far_7_7585_1[0]));    relay_conn far_7_7585_1_b(.in(far_7_7585_0[1]), .out(far_7_7585_1[1]));
    assign out[445] = far_7_7585_1[0]; 
    assign out[446] = layer_6[122] & ~layer_6[117]; 
    wire [1:0] far_7_7587_0;    relay_conn far_7_7587_0_a(.in(layer_6[628]), .out(far_7_7587_0[0]));    relay_conn far_7_7587_0_b(.in(layer_6[532]), .out(far_7_7587_0[1]));
    wire [1:0] far_7_7587_1;    relay_conn far_7_7587_1_a(.in(far_7_7587_0[0]), .out(far_7_7587_1[0]));    relay_conn far_7_7587_1_b(.in(far_7_7587_0[1]), .out(far_7_7587_1[1]));
    wire [1:0] far_7_7587_2;    relay_conn far_7_7587_2_a(.in(far_7_7587_1[0]), .out(far_7_7587_2[0]));    relay_conn far_7_7587_2_b(.in(far_7_7587_1[1]), .out(far_7_7587_2[1]));
    assign out[447] = ~(far_7_7587_2[0] & far_7_7587_2[1]); 
    wire [1:0] far_7_7588_0;    relay_conn far_7_7588_0_a(.in(layer_6[472]), .out(far_7_7588_0[0]));    relay_conn far_7_7588_0_b(.in(layer_6[562]), .out(far_7_7588_0[1]));
    wire [1:0] far_7_7588_1;    relay_conn far_7_7588_1_a(.in(far_7_7588_0[0]), .out(far_7_7588_1[0]));    relay_conn far_7_7588_1_b(.in(far_7_7588_0[1]), .out(far_7_7588_1[1]));
    assign out[448] = ~(far_7_7588_1[0] | far_7_7588_1[1]); 
    wire [1:0] far_7_7589_0;    relay_conn far_7_7589_0_a(.in(layer_6[723]), .out(far_7_7589_0[0]));    relay_conn far_7_7589_0_b(.in(layer_6[788]), .out(far_7_7589_0[1]));
    wire [1:0] far_7_7589_1;    relay_conn far_7_7589_1_a(.in(far_7_7589_0[0]), .out(far_7_7589_1[0]));    relay_conn far_7_7589_1_b(.in(far_7_7589_0[1]), .out(far_7_7589_1[1]));
    assign out[449] = far_7_7589_1[0]; 
    wire [1:0] far_7_7590_0;    relay_conn far_7_7590_0_a(.in(layer_6[827]), .out(far_7_7590_0[0]));    relay_conn far_7_7590_0_b(.in(layer_6[887]), .out(far_7_7590_0[1]));
    assign out[450] = far_7_7590_0[0] ^ far_7_7590_0[1]; 
    wire [1:0] far_7_7591_0;    relay_conn far_7_7591_0_a(.in(layer_6[215]), .out(far_7_7591_0[0]));    relay_conn far_7_7591_0_b(.in(layer_6[136]), .out(far_7_7591_0[1]));
    wire [1:0] far_7_7591_1;    relay_conn far_7_7591_1_a(.in(far_7_7591_0[0]), .out(far_7_7591_1[0]));    relay_conn far_7_7591_1_b(.in(far_7_7591_0[1]), .out(far_7_7591_1[1]));
    assign out[451] = far_7_7591_1[1]; 
    wire [1:0] far_7_7592_0;    relay_conn far_7_7592_0_a(.in(layer_6[777]), .out(far_7_7592_0[0]));    relay_conn far_7_7592_0_b(.in(layer_6[721]), .out(far_7_7592_0[1]));
    assign out[452] = far_7_7592_0[1] & ~far_7_7592_0[0]; 
    assign out[453] = ~layer_6[821]; 
    wire [1:0] far_7_7594_0;    relay_conn far_7_7594_0_a(.in(layer_6[360]), .out(far_7_7594_0[0]));    relay_conn far_7_7594_0_b(.in(layer_6[461]), .out(far_7_7594_0[1]));
    wire [1:0] far_7_7594_1;    relay_conn far_7_7594_1_a(.in(far_7_7594_0[0]), .out(far_7_7594_1[0]));    relay_conn far_7_7594_1_b(.in(far_7_7594_0[1]), .out(far_7_7594_1[1]));
    wire [1:0] far_7_7594_2;    relay_conn far_7_7594_2_a(.in(far_7_7594_1[0]), .out(far_7_7594_2[0]));    relay_conn far_7_7594_2_b(.in(far_7_7594_1[1]), .out(far_7_7594_2[1]));
    assign out[454] = far_7_7594_2[1] & ~far_7_7594_2[0]; 
    assign out[455] = layer_6[717]; 
    wire [1:0] far_7_7596_0;    relay_conn far_7_7596_0_a(.in(layer_6[56]), .out(far_7_7596_0[0]));    relay_conn far_7_7596_0_b(.in(layer_6[128]), .out(far_7_7596_0[1]));
    wire [1:0] far_7_7596_1;    relay_conn far_7_7596_1_a(.in(far_7_7596_0[0]), .out(far_7_7596_1[0]));    relay_conn far_7_7596_1_b(.in(far_7_7596_0[1]), .out(far_7_7596_1[1]));
    assign out[456] = ~(far_7_7596_1[0] ^ far_7_7596_1[1]); 
    assign out[457] = layer_6[599] & ~layer_6[629]; 
    wire [1:0] far_7_7598_0;    relay_conn far_7_7598_0_a(.in(layer_6[779]), .out(far_7_7598_0[0]));    relay_conn far_7_7598_0_b(.in(layer_6[846]), .out(far_7_7598_0[1]));
    wire [1:0] far_7_7598_1;    relay_conn far_7_7598_1_a(.in(far_7_7598_0[0]), .out(far_7_7598_1[0]));    relay_conn far_7_7598_1_b(.in(far_7_7598_0[1]), .out(far_7_7598_1[1]));
    assign out[458] = far_7_7598_1[0] ^ far_7_7598_1[1]; 
    assign out[459] = layer_6[822]; 
    wire [1:0] far_7_7600_0;    relay_conn far_7_7600_0_a(.in(layer_6[315]), .out(far_7_7600_0[0]));    relay_conn far_7_7600_0_b(.in(layer_6[197]), .out(far_7_7600_0[1]));
    wire [1:0] far_7_7600_1;    relay_conn far_7_7600_1_a(.in(far_7_7600_0[0]), .out(far_7_7600_1[0]));    relay_conn far_7_7600_1_b(.in(far_7_7600_0[1]), .out(far_7_7600_1[1]));
    wire [1:0] far_7_7600_2;    relay_conn far_7_7600_2_a(.in(far_7_7600_1[0]), .out(far_7_7600_2[0]));    relay_conn far_7_7600_2_b(.in(far_7_7600_1[1]), .out(far_7_7600_2[1]));
    assign out[460] = far_7_7600_2[0]; 
    assign out[461] = layer_6[333] ^ layer_6[303]; 
    wire [1:0] far_7_7602_0;    relay_conn far_7_7602_0_a(.in(layer_6[448]), .out(far_7_7602_0[0]));    relay_conn far_7_7602_0_b(.in(layer_6[393]), .out(far_7_7602_0[1]));
    assign out[462] = far_7_7602_0[0] & ~far_7_7602_0[1]; 
    wire [1:0] far_7_7603_0;    relay_conn far_7_7603_0_a(.in(layer_6[318]), .out(far_7_7603_0[0]));    relay_conn far_7_7603_0_b(.in(layer_6[387]), .out(far_7_7603_0[1]));
    wire [1:0] far_7_7603_1;    relay_conn far_7_7603_1_a(.in(far_7_7603_0[0]), .out(far_7_7603_1[0]));    relay_conn far_7_7603_1_b(.in(far_7_7603_0[1]), .out(far_7_7603_1[1]));
    assign out[463] = ~(far_7_7603_1[0] ^ far_7_7603_1[1]); 
    assign out[464] = ~(layer_6[284] | layer_6[299]); 
    wire [1:0] far_7_7605_0;    relay_conn far_7_7605_0_a(.in(layer_6[416]), .out(far_7_7605_0[0]));    relay_conn far_7_7605_0_b(.in(layer_6[497]), .out(far_7_7605_0[1]));
    wire [1:0] far_7_7605_1;    relay_conn far_7_7605_1_a(.in(far_7_7605_0[0]), .out(far_7_7605_1[0]));    relay_conn far_7_7605_1_b(.in(far_7_7605_0[1]), .out(far_7_7605_1[1]));
    assign out[465] = ~far_7_7605_1[1]; 
    wire [1:0] far_7_7606_0;    relay_conn far_7_7606_0_a(.in(layer_6[468]), .out(far_7_7606_0[0]));    relay_conn far_7_7606_0_b(.in(layer_6[510]), .out(far_7_7606_0[1]));
    assign out[466] = far_7_7606_0[1]; 
    wire [1:0] far_7_7607_0;    relay_conn far_7_7607_0_a(.in(layer_6[534]), .out(far_7_7607_0[0]));    relay_conn far_7_7607_0_b(.in(layer_6[499]), .out(far_7_7607_0[1]));
    assign out[467] = far_7_7607_0[0]; 
    wire [1:0] far_7_7608_0;    relay_conn far_7_7608_0_a(.in(layer_6[764]), .out(far_7_7608_0[0]));    relay_conn far_7_7608_0_b(.in(layer_6[814]), .out(far_7_7608_0[1]));
    assign out[468] = far_7_7608_0[0]; 
    assign out[469] = ~layer_6[777]; 
    wire [1:0] far_7_7610_0;    relay_conn far_7_7610_0_a(.in(layer_6[811]), .out(far_7_7610_0[0]));    relay_conn far_7_7610_0_b(.in(layer_6[845]), .out(far_7_7610_0[1]));
    assign out[470] = far_7_7610_0[0] & far_7_7610_0[1]; 
    wire [1:0] far_7_7611_0;    relay_conn far_7_7611_0_a(.in(layer_6[398]), .out(far_7_7611_0[0]));    relay_conn far_7_7611_0_b(.in(layer_6[319]), .out(far_7_7611_0[1]));
    wire [1:0] far_7_7611_1;    relay_conn far_7_7611_1_a(.in(far_7_7611_0[0]), .out(far_7_7611_1[0]));    relay_conn far_7_7611_1_b(.in(far_7_7611_0[1]), .out(far_7_7611_1[1]));
    assign out[471] = ~far_7_7611_1[1]; 
    wire [1:0] far_7_7612_0;    relay_conn far_7_7612_0_a(.in(layer_6[691]), .out(far_7_7612_0[0]));    relay_conn far_7_7612_0_b(.in(layer_6[626]), .out(far_7_7612_0[1]));
    wire [1:0] far_7_7612_1;    relay_conn far_7_7612_1_a(.in(far_7_7612_0[0]), .out(far_7_7612_1[0]));    relay_conn far_7_7612_1_b(.in(far_7_7612_0[1]), .out(far_7_7612_1[1]));
    assign out[472] = far_7_7612_1[0] & far_7_7612_1[1]; 
    wire [1:0] far_7_7613_0;    relay_conn far_7_7613_0_a(.in(layer_6[682]), .out(far_7_7613_0[0]));    relay_conn far_7_7613_0_b(.in(layer_6[582]), .out(far_7_7613_0[1]));
    wire [1:0] far_7_7613_1;    relay_conn far_7_7613_1_a(.in(far_7_7613_0[0]), .out(far_7_7613_1[0]));    relay_conn far_7_7613_1_b(.in(far_7_7613_0[1]), .out(far_7_7613_1[1]));
    wire [1:0] far_7_7613_2;    relay_conn far_7_7613_2_a(.in(far_7_7613_1[0]), .out(far_7_7613_2[0]));    relay_conn far_7_7613_2_b(.in(far_7_7613_1[1]), .out(far_7_7613_2[1]));
    assign out[473] = far_7_7613_2[0] & ~far_7_7613_2[1]; 
    wire [1:0] far_7_7614_0;    relay_conn far_7_7614_0_a(.in(layer_6[358]), .out(far_7_7614_0[0]));    relay_conn far_7_7614_0_b(.in(layer_6[442]), .out(far_7_7614_0[1]));
    wire [1:0] far_7_7614_1;    relay_conn far_7_7614_1_a(.in(far_7_7614_0[0]), .out(far_7_7614_1[0]));    relay_conn far_7_7614_1_b(.in(far_7_7614_0[1]), .out(far_7_7614_1[1]));
    assign out[474] = ~(far_7_7614_1[0] ^ far_7_7614_1[1]); 
    assign out[475] = ~(layer_6[744] | layer_6[767]); 
    wire [1:0] far_7_7616_0;    relay_conn far_7_7616_0_a(.in(layer_6[76]), .out(far_7_7616_0[0]));    relay_conn far_7_7616_0_b(.in(layer_6[38]), .out(far_7_7616_0[1]));
    assign out[476] = far_7_7616_0[1] & ~far_7_7616_0[0]; 
    wire [1:0] far_7_7617_0;    relay_conn far_7_7617_0_a(.in(layer_6[450]), .out(far_7_7617_0[0]));    relay_conn far_7_7617_0_b(.in(layer_6[575]), .out(far_7_7617_0[1]));
    wire [1:0] far_7_7617_1;    relay_conn far_7_7617_1_a(.in(far_7_7617_0[0]), .out(far_7_7617_1[0]));    relay_conn far_7_7617_1_b(.in(far_7_7617_0[1]), .out(far_7_7617_1[1]));
    wire [1:0] far_7_7617_2;    relay_conn far_7_7617_2_a(.in(far_7_7617_1[0]), .out(far_7_7617_2[0]));    relay_conn far_7_7617_2_b(.in(far_7_7617_1[1]), .out(far_7_7617_2[1]));
    assign out[477] = far_7_7617_2[1]; 
    wire [1:0] far_7_7618_0;    relay_conn far_7_7618_0_a(.in(layer_6[896]), .out(far_7_7618_0[0]));    relay_conn far_7_7618_0_b(.in(layer_6[848]), .out(far_7_7618_0[1]));
    assign out[478] = far_7_7618_0[1]; 
    wire [1:0] far_7_7619_0;    relay_conn far_7_7619_0_a(.in(layer_6[913]), .out(far_7_7619_0[0]));    relay_conn far_7_7619_0_b(.in(layer_6[794]), .out(far_7_7619_0[1]));
    wire [1:0] far_7_7619_1;    relay_conn far_7_7619_1_a(.in(far_7_7619_0[0]), .out(far_7_7619_1[0]));    relay_conn far_7_7619_1_b(.in(far_7_7619_0[1]), .out(far_7_7619_1[1]));
    wire [1:0] far_7_7619_2;    relay_conn far_7_7619_2_a(.in(far_7_7619_1[0]), .out(far_7_7619_2[0]));    relay_conn far_7_7619_2_b(.in(far_7_7619_1[1]), .out(far_7_7619_2[1]));
    assign out[479] = far_7_7619_2[1] & ~far_7_7619_2[0]; 
    assign out[480] = layer_6[22]; 
    wire [1:0] far_7_7621_0;    relay_conn far_7_7621_0_a(.in(layer_6[613]), .out(far_7_7621_0[0]));    relay_conn far_7_7621_0_b(.in(layer_6[534]), .out(far_7_7621_0[1]));
    wire [1:0] far_7_7621_1;    relay_conn far_7_7621_1_a(.in(far_7_7621_0[0]), .out(far_7_7621_1[0]));    relay_conn far_7_7621_1_b(.in(far_7_7621_0[1]), .out(far_7_7621_1[1]));
    assign out[481] = ~far_7_7621_1[0]; 
    assign out[482] = ~(layer_6[802] | layer_6[812]); 
    wire [1:0] far_7_7623_0;    relay_conn far_7_7623_0_a(.in(layer_6[30]), .out(far_7_7623_0[0]));    relay_conn far_7_7623_0_b(.in(layer_6[143]), .out(far_7_7623_0[1]));
    wire [1:0] far_7_7623_1;    relay_conn far_7_7623_1_a(.in(far_7_7623_0[0]), .out(far_7_7623_1[0]));    relay_conn far_7_7623_1_b(.in(far_7_7623_0[1]), .out(far_7_7623_1[1]));
    wire [1:0] far_7_7623_2;    relay_conn far_7_7623_2_a(.in(far_7_7623_1[0]), .out(far_7_7623_2[0]));    relay_conn far_7_7623_2_b(.in(far_7_7623_1[1]), .out(far_7_7623_2[1]));
    assign out[483] = far_7_7623_2[0] & far_7_7623_2[1]; 
    wire [1:0] far_7_7624_0;    relay_conn far_7_7624_0_a(.in(layer_6[773]), .out(far_7_7624_0[0]));    relay_conn far_7_7624_0_b(.in(layer_6[673]), .out(far_7_7624_0[1]));
    wire [1:0] far_7_7624_1;    relay_conn far_7_7624_1_a(.in(far_7_7624_0[0]), .out(far_7_7624_1[0]));    relay_conn far_7_7624_1_b(.in(far_7_7624_0[1]), .out(far_7_7624_1[1]));
    wire [1:0] far_7_7624_2;    relay_conn far_7_7624_2_a(.in(far_7_7624_1[0]), .out(far_7_7624_2[0]));    relay_conn far_7_7624_2_b(.in(far_7_7624_1[1]), .out(far_7_7624_2[1]));
    assign out[484] = far_7_7624_2[1]; 
    wire [1:0] far_7_7625_0;    relay_conn far_7_7625_0_a(.in(layer_6[416]), .out(far_7_7625_0[0]));    relay_conn far_7_7625_0_b(.in(layer_6[478]), .out(far_7_7625_0[1]));
    assign out[485] = ~far_7_7625_0[1]; 
    wire [1:0] far_7_7626_0;    relay_conn far_7_7626_0_a(.in(layer_6[205]), .out(far_7_7626_0[0]));    relay_conn far_7_7626_0_b(.in(layer_6[304]), .out(far_7_7626_0[1]));
    wire [1:0] far_7_7626_1;    relay_conn far_7_7626_1_a(.in(far_7_7626_0[0]), .out(far_7_7626_1[0]));    relay_conn far_7_7626_1_b(.in(far_7_7626_0[1]), .out(far_7_7626_1[1]));
    wire [1:0] far_7_7626_2;    relay_conn far_7_7626_2_a(.in(far_7_7626_1[0]), .out(far_7_7626_2[0]));    relay_conn far_7_7626_2_b(.in(far_7_7626_1[1]), .out(far_7_7626_2[1]));
    assign out[486] = far_7_7626_2[0] & ~far_7_7626_2[1]; 
    wire [1:0] far_7_7627_0;    relay_conn far_7_7627_0_a(.in(layer_6[45]), .out(far_7_7627_0[0]));    relay_conn far_7_7627_0_b(.in(layer_6[6]), .out(far_7_7627_0[1]));
    assign out[487] = far_7_7627_0[0] & far_7_7627_0[1]; 
    wire [1:0] far_7_7628_0;    relay_conn far_7_7628_0_a(.in(layer_6[308]), .out(far_7_7628_0[0]));    relay_conn far_7_7628_0_b(.in(layer_6[230]), .out(far_7_7628_0[1]));
    wire [1:0] far_7_7628_1;    relay_conn far_7_7628_1_a(.in(far_7_7628_0[0]), .out(far_7_7628_1[0]));    relay_conn far_7_7628_1_b(.in(far_7_7628_0[1]), .out(far_7_7628_1[1]));
    assign out[488] = far_7_7628_1[1] & ~far_7_7628_1[0]; 
    assign out[489] = ~(layer_6[981] | layer_6[954]); 
    wire [1:0] far_7_7630_0;    relay_conn far_7_7630_0_a(.in(layer_6[21]), .out(far_7_7630_0[0]));    relay_conn far_7_7630_0_b(.in(layer_6[146]), .out(far_7_7630_0[1]));
    wire [1:0] far_7_7630_1;    relay_conn far_7_7630_1_a(.in(far_7_7630_0[0]), .out(far_7_7630_1[0]));    relay_conn far_7_7630_1_b(.in(far_7_7630_0[1]), .out(far_7_7630_1[1]));
    wire [1:0] far_7_7630_2;    relay_conn far_7_7630_2_a(.in(far_7_7630_1[0]), .out(far_7_7630_2[0]));    relay_conn far_7_7630_2_b(.in(far_7_7630_1[1]), .out(far_7_7630_2[1]));
    assign out[490] = ~far_7_7630_2[0]; 
    wire [1:0] far_7_7631_0;    relay_conn far_7_7631_0_a(.in(layer_6[476]), .out(far_7_7631_0[0]));    relay_conn far_7_7631_0_b(.in(layer_6[425]), .out(far_7_7631_0[1]));
    assign out[491] = far_7_7631_0[1] & ~far_7_7631_0[0]; 
    assign out[492] = layer_6[526] & layer_6[516]; 
    assign out[493] = ~(layer_6[675] & layer_6[703]); 
    wire [1:0] far_7_7634_0;    relay_conn far_7_7634_0_a(.in(layer_6[908]), .out(far_7_7634_0[0]));    relay_conn far_7_7634_0_b(.in(layer_6[1016]), .out(far_7_7634_0[1]));
    wire [1:0] far_7_7634_1;    relay_conn far_7_7634_1_a(.in(far_7_7634_0[0]), .out(far_7_7634_1[0]));    relay_conn far_7_7634_1_b(.in(far_7_7634_0[1]), .out(far_7_7634_1[1]));
    wire [1:0] far_7_7634_2;    relay_conn far_7_7634_2_a(.in(far_7_7634_1[0]), .out(far_7_7634_2[0]));    relay_conn far_7_7634_2_b(.in(far_7_7634_1[1]), .out(far_7_7634_2[1]));
    assign out[494] = far_7_7634_2[1]; 
    wire [1:0] far_7_7635_0;    relay_conn far_7_7635_0_a(.in(layer_6[903]), .out(far_7_7635_0[0]));    relay_conn far_7_7635_0_b(.in(layer_6[802]), .out(far_7_7635_0[1]));
    wire [1:0] far_7_7635_1;    relay_conn far_7_7635_1_a(.in(far_7_7635_0[0]), .out(far_7_7635_1[0]));    relay_conn far_7_7635_1_b(.in(far_7_7635_0[1]), .out(far_7_7635_1[1]));
    wire [1:0] far_7_7635_2;    relay_conn far_7_7635_2_a(.in(far_7_7635_1[0]), .out(far_7_7635_2[0]));    relay_conn far_7_7635_2_b(.in(far_7_7635_1[1]), .out(far_7_7635_2[1]));
    assign out[495] = ~(far_7_7635_2[0] | far_7_7635_2[1]); 
    wire [1:0] far_7_7636_0;    relay_conn far_7_7636_0_a(.in(layer_6[778]), .out(far_7_7636_0[0]));    relay_conn far_7_7636_0_b(.in(layer_6[660]), .out(far_7_7636_0[1]));
    wire [1:0] far_7_7636_1;    relay_conn far_7_7636_1_a(.in(far_7_7636_0[0]), .out(far_7_7636_1[0]));    relay_conn far_7_7636_1_b(.in(far_7_7636_0[1]), .out(far_7_7636_1[1]));
    wire [1:0] far_7_7636_2;    relay_conn far_7_7636_2_a(.in(far_7_7636_1[0]), .out(far_7_7636_2[0]));    relay_conn far_7_7636_2_b(.in(far_7_7636_1[1]), .out(far_7_7636_2[1]));
    assign out[496] = far_7_7636_2[1]; 
    assign out[497] = layer_6[678] & ~layer_6[648]; 
    wire [1:0] far_7_7638_0;    relay_conn far_7_7638_0_a(.in(layer_6[822]), .out(far_7_7638_0[0]));    relay_conn far_7_7638_0_b(.in(layer_6[778]), .out(far_7_7638_0[1]));
    assign out[498] = far_7_7638_0[0]; 
    assign out[499] = layer_6[510]; 
    wire [1:0] far_7_7640_0;    relay_conn far_7_7640_0_a(.in(layer_6[742]), .out(far_7_7640_0[0]));    relay_conn far_7_7640_0_b(.in(layer_6[793]), .out(far_7_7640_0[1]));
    assign out[500] = ~far_7_7640_0[0]; 
    wire [1:0] far_7_7641_0;    relay_conn far_7_7641_0_a(.in(layer_6[605]), .out(far_7_7641_0[0]));    relay_conn far_7_7641_0_b(.in(layer_6[643]), .out(far_7_7641_0[1]));
    assign out[501] = far_7_7641_0[1]; 
    wire [1:0] far_7_7642_0;    relay_conn far_7_7642_0_a(.in(layer_6[539]), .out(far_7_7642_0[0]));    relay_conn far_7_7642_0_b(.in(layer_6[460]), .out(far_7_7642_0[1]));
    wire [1:0] far_7_7642_1;    relay_conn far_7_7642_1_a(.in(far_7_7642_0[0]), .out(far_7_7642_1[0]));    relay_conn far_7_7642_1_b(.in(far_7_7642_0[1]), .out(far_7_7642_1[1]));
    assign out[502] = ~(far_7_7642_1[0] | far_7_7642_1[1]); 
    wire [1:0] far_7_7643_0;    relay_conn far_7_7643_0_a(.in(layer_6[866]), .out(far_7_7643_0[0]));    relay_conn far_7_7643_0_b(.in(layer_6[942]), .out(far_7_7643_0[1]));
    wire [1:0] far_7_7643_1;    relay_conn far_7_7643_1_a(.in(far_7_7643_0[0]), .out(far_7_7643_1[0]));    relay_conn far_7_7643_1_b(.in(far_7_7643_0[1]), .out(far_7_7643_1[1]));
    assign out[503] = ~(far_7_7643_1[0] | far_7_7643_1[1]); 
    wire [1:0] far_7_7644_0;    relay_conn far_7_7644_0_a(.in(layer_6[422]), .out(far_7_7644_0[0]));    relay_conn far_7_7644_0_b(.in(layer_6[456]), .out(far_7_7644_0[1]));
    assign out[504] = far_7_7644_0[0]; 
    wire [1:0] far_7_7645_0;    relay_conn far_7_7645_0_a(.in(layer_6[456]), .out(far_7_7645_0[0]));    relay_conn far_7_7645_0_b(.in(layer_6[388]), .out(far_7_7645_0[1]));
    wire [1:0] far_7_7645_1;    relay_conn far_7_7645_1_a(.in(far_7_7645_0[0]), .out(far_7_7645_1[0]));    relay_conn far_7_7645_1_b(.in(far_7_7645_0[1]), .out(far_7_7645_1[1]));
    assign out[505] = ~far_7_7645_1[1]; 
    wire [1:0] far_7_7646_0;    relay_conn far_7_7646_0_a(.in(layer_6[419]), .out(far_7_7646_0[0]));    relay_conn far_7_7646_0_b(.in(layer_6[321]), .out(far_7_7646_0[1]));
    wire [1:0] far_7_7646_1;    relay_conn far_7_7646_1_a(.in(far_7_7646_0[0]), .out(far_7_7646_1[0]));    relay_conn far_7_7646_1_b(.in(far_7_7646_0[1]), .out(far_7_7646_1[1]));
    wire [1:0] far_7_7646_2;    relay_conn far_7_7646_2_a(.in(far_7_7646_1[0]), .out(far_7_7646_2[0]));    relay_conn far_7_7646_2_b(.in(far_7_7646_1[1]), .out(far_7_7646_2[1]));
    assign out[506] = far_7_7646_2[0] & ~far_7_7646_2[1]; 
    assign out[507] = ~(layer_6[220] | layer_6[222]); 
    wire [1:0] far_7_7648_0;    relay_conn far_7_7648_0_a(.in(layer_6[852]), .out(far_7_7648_0[0]));    relay_conn far_7_7648_0_b(.in(layer_6[799]), .out(far_7_7648_0[1]));
    assign out[508] = ~far_7_7648_0[0]; 
    wire [1:0] far_7_7649_0;    relay_conn far_7_7649_0_a(.in(layer_6[62]), .out(far_7_7649_0[0]));    relay_conn far_7_7649_0_b(.in(layer_6[187]), .out(far_7_7649_0[1]));
    wire [1:0] far_7_7649_1;    relay_conn far_7_7649_1_a(.in(far_7_7649_0[0]), .out(far_7_7649_1[0]));    relay_conn far_7_7649_1_b(.in(far_7_7649_0[1]), .out(far_7_7649_1[1]));
    wire [1:0] far_7_7649_2;    relay_conn far_7_7649_2_a(.in(far_7_7649_1[0]), .out(far_7_7649_2[0]));    relay_conn far_7_7649_2_b(.in(far_7_7649_1[1]), .out(far_7_7649_2[1]));
    assign out[509] = far_7_7649_2[0]; 
    wire [1:0] far_7_7650_0;    relay_conn far_7_7650_0_a(.in(layer_6[826]), .out(far_7_7650_0[0]));    relay_conn far_7_7650_0_b(.in(layer_6[886]), .out(far_7_7650_0[1]));
    assign out[510] = far_7_7650_0[1]; 
    assign out[511] = layer_6[591] & ~layer_6[601]; 
    wire [1:0] far_7_7652_0;    relay_conn far_7_7652_0_a(.in(layer_6[226]), .out(far_7_7652_0[0]));    relay_conn far_7_7652_0_b(.in(layer_6[183]), .out(far_7_7652_0[1]));
    assign out[512] = far_7_7652_0[1] & ~far_7_7652_0[0]; 
    assign out[513] = ~(layer_6[57] | layer_6[88]); 
    wire [1:0] far_7_7654_0;    relay_conn far_7_7654_0_a(.in(layer_6[496]), .out(far_7_7654_0[0]));    relay_conn far_7_7654_0_b(.in(layer_6[597]), .out(far_7_7654_0[1]));
    wire [1:0] far_7_7654_1;    relay_conn far_7_7654_1_a(.in(far_7_7654_0[0]), .out(far_7_7654_1[0]));    relay_conn far_7_7654_1_b(.in(far_7_7654_0[1]), .out(far_7_7654_1[1]));
    wire [1:0] far_7_7654_2;    relay_conn far_7_7654_2_a(.in(far_7_7654_1[0]), .out(far_7_7654_2[0]));    relay_conn far_7_7654_2_b(.in(far_7_7654_1[1]), .out(far_7_7654_2[1]));
    assign out[514] = far_7_7654_2[0] & ~far_7_7654_2[1]; 
    wire [1:0] far_7_7655_0;    relay_conn far_7_7655_0_a(.in(layer_6[919]), .out(far_7_7655_0[0]));    relay_conn far_7_7655_0_b(.in(layer_6[834]), .out(far_7_7655_0[1]));
    wire [1:0] far_7_7655_1;    relay_conn far_7_7655_1_a(.in(far_7_7655_0[0]), .out(far_7_7655_1[0]));    relay_conn far_7_7655_1_b(.in(far_7_7655_0[1]), .out(far_7_7655_1[1]));
    assign out[515] = far_7_7655_1[0] & far_7_7655_1[1]; 
    assign out[516] = layer_6[808] & ~layer_6[814]; 
    wire [1:0] far_7_7657_0;    relay_conn far_7_7657_0_a(.in(layer_6[574]), .out(far_7_7657_0[0]));    relay_conn far_7_7657_0_b(.in(layer_6[645]), .out(far_7_7657_0[1]));
    wire [1:0] far_7_7657_1;    relay_conn far_7_7657_1_a(.in(far_7_7657_0[0]), .out(far_7_7657_1[0]));    relay_conn far_7_7657_1_b(.in(far_7_7657_0[1]), .out(far_7_7657_1[1]));
    assign out[517] = ~far_7_7657_1[1]; 
    wire [1:0] far_7_7658_0;    relay_conn far_7_7658_0_a(.in(layer_6[410]), .out(far_7_7658_0[0]));    relay_conn far_7_7658_0_b(.in(layer_6[511]), .out(far_7_7658_0[1]));
    wire [1:0] far_7_7658_1;    relay_conn far_7_7658_1_a(.in(far_7_7658_0[0]), .out(far_7_7658_1[0]));    relay_conn far_7_7658_1_b(.in(far_7_7658_0[1]), .out(far_7_7658_1[1]));
    wire [1:0] far_7_7658_2;    relay_conn far_7_7658_2_a(.in(far_7_7658_1[0]), .out(far_7_7658_2[0]));    relay_conn far_7_7658_2_b(.in(far_7_7658_1[1]), .out(far_7_7658_2[1]));
    assign out[518] = far_7_7658_2[1] & ~far_7_7658_2[0]; 
    wire [1:0] far_7_7659_0;    relay_conn far_7_7659_0_a(.in(layer_6[80]), .out(far_7_7659_0[0]));    relay_conn far_7_7659_0_b(.in(layer_6[12]), .out(far_7_7659_0[1]));
    wire [1:0] far_7_7659_1;    relay_conn far_7_7659_1_a(.in(far_7_7659_0[0]), .out(far_7_7659_1[0]));    relay_conn far_7_7659_1_b(.in(far_7_7659_0[1]), .out(far_7_7659_1[1]));
    assign out[519] = ~(far_7_7659_1[0] ^ far_7_7659_1[1]); 
    wire [1:0] far_7_7660_0;    relay_conn far_7_7660_0_a(.in(layer_6[982]), .out(far_7_7660_0[0]));    relay_conn far_7_7660_0_b(.in(layer_6[892]), .out(far_7_7660_0[1]));
    wire [1:0] far_7_7660_1;    relay_conn far_7_7660_1_a(.in(far_7_7660_0[0]), .out(far_7_7660_1[0]));    relay_conn far_7_7660_1_b(.in(far_7_7660_0[1]), .out(far_7_7660_1[1]));
    assign out[520] = ~(far_7_7660_1[0] | far_7_7660_1[1]); 
    wire [1:0] far_7_7661_0;    relay_conn far_7_7661_0_a(.in(layer_6[273]), .out(far_7_7661_0[0]));    relay_conn far_7_7661_0_b(.in(layer_6[370]), .out(far_7_7661_0[1]));
    wire [1:0] far_7_7661_1;    relay_conn far_7_7661_1_a(.in(far_7_7661_0[0]), .out(far_7_7661_1[0]));    relay_conn far_7_7661_1_b(.in(far_7_7661_0[1]), .out(far_7_7661_1[1]));
    wire [1:0] far_7_7661_2;    relay_conn far_7_7661_2_a(.in(far_7_7661_1[0]), .out(far_7_7661_2[0]));    relay_conn far_7_7661_2_b(.in(far_7_7661_1[1]), .out(far_7_7661_2[1]));
    assign out[521] = far_7_7661_2[0] ^ far_7_7661_2[1]; 
    wire [1:0] far_7_7662_0;    relay_conn far_7_7662_0_a(.in(layer_6[478]), .out(far_7_7662_0[0]));    relay_conn far_7_7662_0_b(.in(layer_6[401]), .out(far_7_7662_0[1]));
    wire [1:0] far_7_7662_1;    relay_conn far_7_7662_1_a(.in(far_7_7662_0[0]), .out(far_7_7662_1[0]));    relay_conn far_7_7662_1_b(.in(far_7_7662_0[1]), .out(far_7_7662_1[1]));
    assign out[522] = far_7_7662_1[1] & ~far_7_7662_1[0]; 
    wire [1:0] far_7_7663_0;    relay_conn far_7_7663_0_a(.in(layer_6[633]), .out(far_7_7663_0[0]));    relay_conn far_7_7663_0_b(.in(layer_6[539]), .out(far_7_7663_0[1]));
    wire [1:0] far_7_7663_1;    relay_conn far_7_7663_1_a(.in(far_7_7663_0[0]), .out(far_7_7663_1[0]));    relay_conn far_7_7663_1_b(.in(far_7_7663_0[1]), .out(far_7_7663_1[1]));
    assign out[523] = far_7_7663_1[0] & ~far_7_7663_1[1]; 
    wire [1:0] far_7_7664_0;    relay_conn far_7_7664_0_a(.in(layer_6[575]), .out(far_7_7664_0[0]));    relay_conn far_7_7664_0_b(.in(layer_6[659]), .out(far_7_7664_0[1]));
    wire [1:0] far_7_7664_1;    relay_conn far_7_7664_1_a(.in(far_7_7664_0[0]), .out(far_7_7664_1[0]));    relay_conn far_7_7664_1_b(.in(far_7_7664_0[1]), .out(far_7_7664_1[1]));
    assign out[524] = ~far_7_7664_1[0]; 
    wire [1:0] far_7_7665_0;    relay_conn far_7_7665_0_a(.in(layer_6[157]), .out(far_7_7665_0[0]));    relay_conn far_7_7665_0_b(.in(layer_6[88]), .out(far_7_7665_0[1]));
    wire [1:0] far_7_7665_1;    relay_conn far_7_7665_1_a(.in(far_7_7665_0[0]), .out(far_7_7665_1[0]));    relay_conn far_7_7665_1_b(.in(far_7_7665_0[1]), .out(far_7_7665_1[1]));
    assign out[525] = far_7_7665_1[0]; 
    wire [1:0] far_7_7666_0;    relay_conn far_7_7666_0_a(.in(layer_6[930]), .out(far_7_7666_0[0]));    relay_conn far_7_7666_0_b(.in(layer_6[1008]), .out(far_7_7666_0[1]));
    wire [1:0] far_7_7666_1;    relay_conn far_7_7666_1_a(.in(far_7_7666_0[0]), .out(far_7_7666_1[0]));    relay_conn far_7_7666_1_b(.in(far_7_7666_0[1]), .out(far_7_7666_1[1]));
    assign out[526] = far_7_7666_1[1] & ~far_7_7666_1[0]; 
    assign out[527] = ~(layer_6[295] | layer_6[299]); 
    wire [1:0] far_7_7668_0;    relay_conn far_7_7668_0_a(.in(layer_6[883]), .out(far_7_7668_0[0]));    relay_conn far_7_7668_0_b(.in(layer_6[777]), .out(far_7_7668_0[1]));
    wire [1:0] far_7_7668_1;    relay_conn far_7_7668_1_a(.in(far_7_7668_0[0]), .out(far_7_7668_1[0]));    relay_conn far_7_7668_1_b(.in(far_7_7668_0[1]), .out(far_7_7668_1[1]));
    wire [1:0] far_7_7668_2;    relay_conn far_7_7668_2_a(.in(far_7_7668_1[0]), .out(far_7_7668_2[0]));    relay_conn far_7_7668_2_b(.in(far_7_7668_1[1]), .out(far_7_7668_2[1]));
    assign out[528] = far_7_7668_2[1] & ~far_7_7668_2[0]; 
    wire [1:0] far_7_7669_0;    relay_conn far_7_7669_0_a(.in(layer_6[376]), .out(far_7_7669_0[0]));    relay_conn far_7_7669_0_b(.in(layer_6[251]), .out(far_7_7669_0[1]));
    wire [1:0] far_7_7669_1;    relay_conn far_7_7669_1_a(.in(far_7_7669_0[0]), .out(far_7_7669_1[0]));    relay_conn far_7_7669_1_b(.in(far_7_7669_0[1]), .out(far_7_7669_1[1]));
    wire [1:0] far_7_7669_2;    relay_conn far_7_7669_2_a(.in(far_7_7669_1[0]), .out(far_7_7669_2[0]));    relay_conn far_7_7669_2_b(.in(far_7_7669_1[1]), .out(far_7_7669_2[1]));
    assign out[529] = far_7_7669_2[1]; 
    wire [1:0] far_7_7670_0;    relay_conn far_7_7670_0_a(.in(layer_6[394]), .out(far_7_7670_0[0]));    relay_conn far_7_7670_0_b(.in(layer_6[297]), .out(far_7_7670_0[1]));
    wire [1:0] far_7_7670_1;    relay_conn far_7_7670_1_a(.in(far_7_7670_0[0]), .out(far_7_7670_1[0]));    relay_conn far_7_7670_1_b(.in(far_7_7670_0[1]), .out(far_7_7670_1[1]));
    wire [1:0] far_7_7670_2;    relay_conn far_7_7670_2_a(.in(far_7_7670_1[0]), .out(far_7_7670_2[0]));    relay_conn far_7_7670_2_b(.in(far_7_7670_1[1]), .out(far_7_7670_2[1]));
    assign out[530] = far_7_7670_2[0] & far_7_7670_2[1]; 
    wire [1:0] far_7_7671_0;    relay_conn far_7_7671_0_a(.in(layer_6[557]), .out(far_7_7671_0[0]));    relay_conn far_7_7671_0_b(.in(layer_6[449]), .out(far_7_7671_0[1]));
    wire [1:0] far_7_7671_1;    relay_conn far_7_7671_1_a(.in(far_7_7671_0[0]), .out(far_7_7671_1[0]));    relay_conn far_7_7671_1_b(.in(far_7_7671_0[1]), .out(far_7_7671_1[1]));
    wire [1:0] far_7_7671_2;    relay_conn far_7_7671_2_a(.in(far_7_7671_1[0]), .out(far_7_7671_2[0]));    relay_conn far_7_7671_2_b(.in(far_7_7671_1[1]), .out(far_7_7671_2[1]));
    assign out[531] = ~(far_7_7671_2[0] ^ far_7_7671_2[1]); 
    wire [1:0] far_7_7672_0;    relay_conn far_7_7672_0_a(.in(layer_6[184]), .out(far_7_7672_0[0]));    relay_conn far_7_7672_0_b(.in(layer_6[91]), .out(far_7_7672_0[1]));
    wire [1:0] far_7_7672_1;    relay_conn far_7_7672_1_a(.in(far_7_7672_0[0]), .out(far_7_7672_1[0]));    relay_conn far_7_7672_1_b(.in(far_7_7672_0[1]), .out(far_7_7672_1[1]));
    assign out[532] = far_7_7672_1[1]; 
    wire [1:0] far_7_7673_0;    relay_conn far_7_7673_0_a(.in(layer_6[194]), .out(far_7_7673_0[0]));    relay_conn far_7_7673_0_b(.in(layer_6[255]), .out(far_7_7673_0[1]));
    assign out[533] = far_7_7673_0[0]; 
    wire [1:0] far_7_7674_0;    relay_conn far_7_7674_0_a(.in(layer_6[416]), .out(far_7_7674_0[0]));    relay_conn far_7_7674_0_b(.in(layer_6[489]), .out(far_7_7674_0[1]));
    wire [1:0] far_7_7674_1;    relay_conn far_7_7674_1_a(.in(far_7_7674_0[0]), .out(far_7_7674_1[0]));    relay_conn far_7_7674_1_b(.in(far_7_7674_0[1]), .out(far_7_7674_1[1]));
    assign out[534] = far_7_7674_1[0] & far_7_7674_1[1]; 
    wire [1:0] far_7_7675_0;    relay_conn far_7_7675_0_a(.in(layer_6[177]), .out(far_7_7675_0[0]));    relay_conn far_7_7675_0_b(.in(layer_6[273]), .out(far_7_7675_0[1]));
    wire [1:0] far_7_7675_1;    relay_conn far_7_7675_1_a(.in(far_7_7675_0[0]), .out(far_7_7675_1[0]));    relay_conn far_7_7675_1_b(.in(far_7_7675_0[1]), .out(far_7_7675_1[1]));
    wire [1:0] far_7_7675_2;    relay_conn far_7_7675_2_a(.in(far_7_7675_1[0]), .out(far_7_7675_2[0]));    relay_conn far_7_7675_2_b(.in(far_7_7675_1[1]), .out(far_7_7675_2[1]));
    assign out[535] = far_7_7675_2[1] & ~far_7_7675_2[0]; 
    wire [1:0] far_7_7676_0;    relay_conn far_7_7676_0_a(.in(layer_6[681]), .out(far_7_7676_0[0]));    relay_conn far_7_7676_0_b(.in(layer_6[585]), .out(far_7_7676_0[1]));
    wire [1:0] far_7_7676_1;    relay_conn far_7_7676_1_a(.in(far_7_7676_0[0]), .out(far_7_7676_1[0]));    relay_conn far_7_7676_1_b(.in(far_7_7676_0[1]), .out(far_7_7676_1[1]));
    wire [1:0] far_7_7676_2;    relay_conn far_7_7676_2_a(.in(far_7_7676_1[0]), .out(far_7_7676_2[0]));    relay_conn far_7_7676_2_b(.in(far_7_7676_1[1]), .out(far_7_7676_2[1]));
    assign out[536] = far_7_7676_2[1] & ~far_7_7676_2[0]; 
    wire [1:0] far_7_7677_0;    relay_conn far_7_7677_0_a(.in(layer_6[845]), .out(far_7_7677_0[0]));    relay_conn far_7_7677_0_b(.in(layer_6[718]), .out(far_7_7677_0[1]));
    wire [1:0] far_7_7677_1;    relay_conn far_7_7677_1_a(.in(far_7_7677_0[0]), .out(far_7_7677_1[0]));    relay_conn far_7_7677_1_b(.in(far_7_7677_0[1]), .out(far_7_7677_1[1]));
    wire [1:0] far_7_7677_2;    relay_conn far_7_7677_2_a(.in(far_7_7677_1[0]), .out(far_7_7677_2[0]));    relay_conn far_7_7677_2_b(.in(far_7_7677_1[1]), .out(far_7_7677_2[1]));
    assign out[537] = far_7_7677_2[0] & ~far_7_7677_2[1]; 
    wire [1:0] far_7_7678_0;    relay_conn far_7_7678_0_a(.in(layer_6[879]), .out(far_7_7678_0[0]));    relay_conn far_7_7678_0_b(.in(layer_6[760]), .out(far_7_7678_0[1]));
    wire [1:0] far_7_7678_1;    relay_conn far_7_7678_1_a(.in(far_7_7678_0[0]), .out(far_7_7678_1[0]));    relay_conn far_7_7678_1_b(.in(far_7_7678_0[1]), .out(far_7_7678_1[1]));
    wire [1:0] far_7_7678_2;    relay_conn far_7_7678_2_a(.in(far_7_7678_1[0]), .out(far_7_7678_2[0]));    relay_conn far_7_7678_2_b(.in(far_7_7678_1[1]), .out(far_7_7678_2[1]));
    assign out[538] = ~far_7_7678_2[0]; 
    wire [1:0] far_7_7679_0;    relay_conn far_7_7679_0_a(.in(layer_6[56]), .out(far_7_7679_0[0]));    relay_conn far_7_7679_0_b(.in(layer_6[180]), .out(far_7_7679_0[1]));
    wire [1:0] far_7_7679_1;    relay_conn far_7_7679_1_a(.in(far_7_7679_0[0]), .out(far_7_7679_1[0]));    relay_conn far_7_7679_1_b(.in(far_7_7679_0[1]), .out(far_7_7679_1[1]));
    wire [1:0] far_7_7679_2;    relay_conn far_7_7679_2_a(.in(far_7_7679_1[0]), .out(far_7_7679_2[0]));    relay_conn far_7_7679_2_b(.in(far_7_7679_1[1]), .out(far_7_7679_2[1]));
    assign out[539] = far_7_7679_2[0] & far_7_7679_2[1]; 
    wire [1:0] far_7_7680_0;    relay_conn far_7_7680_0_a(.in(layer_6[182]), .out(far_7_7680_0[0]));    relay_conn far_7_7680_0_b(.in(layer_6[72]), .out(far_7_7680_0[1]));
    wire [1:0] far_7_7680_1;    relay_conn far_7_7680_1_a(.in(far_7_7680_0[0]), .out(far_7_7680_1[0]));    relay_conn far_7_7680_1_b(.in(far_7_7680_0[1]), .out(far_7_7680_1[1]));
    wire [1:0] far_7_7680_2;    relay_conn far_7_7680_2_a(.in(far_7_7680_1[0]), .out(far_7_7680_2[0]));    relay_conn far_7_7680_2_b(.in(far_7_7680_1[1]), .out(far_7_7680_2[1]));
    assign out[540] = far_7_7680_2[0] & ~far_7_7680_2[1]; 
    assign out[541] = layer_6[558] & ~layer_6[539]; 
    wire [1:0] far_7_7682_0;    relay_conn far_7_7682_0_a(.in(layer_6[954]), .out(far_7_7682_0[0]));    relay_conn far_7_7682_0_b(.in(layer_6[884]), .out(far_7_7682_0[1]));
    wire [1:0] far_7_7682_1;    relay_conn far_7_7682_1_a(.in(far_7_7682_0[0]), .out(far_7_7682_1[0]));    relay_conn far_7_7682_1_b(.in(far_7_7682_0[1]), .out(far_7_7682_1[1]));
    assign out[542] = far_7_7682_1[0] & ~far_7_7682_1[1]; 
    assign out[543] = layer_6[40] & layer_6[64]; 
    wire [1:0] far_7_7684_0;    relay_conn far_7_7684_0_a(.in(layer_6[171]), .out(far_7_7684_0[0]));    relay_conn far_7_7684_0_b(.in(layer_6[299]), .out(far_7_7684_0[1]));
    wire [1:0] far_7_7684_1;    relay_conn far_7_7684_1_a(.in(far_7_7684_0[0]), .out(far_7_7684_1[0]));    relay_conn far_7_7684_1_b(.in(far_7_7684_0[1]), .out(far_7_7684_1[1]));
    wire [1:0] far_7_7684_2;    relay_conn far_7_7684_2_a(.in(far_7_7684_1[0]), .out(far_7_7684_2[0]));    relay_conn far_7_7684_2_b(.in(far_7_7684_1[1]), .out(far_7_7684_2[1]));
    wire [1:0] far_7_7684_3;    relay_conn far_7_7684_3_a(.in(far_7_7684_2[0]), .out(far_7_7684_3[0]));    relay_conn far_7_7684_3_b(.in(far_7_7684_2[1]), .out(far_7_7684_3[1]));
    assign out[544] = ~(far_7_7684_3[0] | far_7_7684_3[1]); 
    wire [1:0] far_7_7685_0;    relay_conn far_7_7685_0_a(.in(layer_6[142]), .out(far_7_7685_0[0]));    relay_conn far_7_7685_0_b(.in(layer_6[260]), .out(far_7_7685_0[1]));
    wire [1:0] far_7_7685_1;    relay_conn far_7_7685_1_a(.in(far_7_7685_0[0]), .out(far_7_7685_1[0]));    relay_conn far_7_7685_1_b(.in(far_7_7685_0[1]), .out(far_7_7685_1[1]));
    wire [1:0] far_7_7685_2;    relay_conn far_7_7685_2_a(.in(far_7_7685_1[0]), .out(far_7_7685_2[0]));    relay_conn far_7_7685_2_b(.in(far_7_7685_1[1]), .out(far_7_7685_2[1]));
    assign out[545] = far_7_7685_2[0] & ~far_7_7685_2[1]; 
    wire [1:0] far_7_7686_0;    relay_conn far_7_7686_0_a(.in(layer_6[230]), .out(far_7_7686_0[0]));    relay_conn far_7_7686_0_b(.in(layer_6[136]), .out(far_7_7686_0[1]));
    wire [1:0] far_7_7686_1;    relay_conn far_7_7686_1_a(.in(far_7_7686_0[0]), .out(far_7_7686_1[0]));    relay_conn far_7_7686_1_b(.in(far_7_7686_0[1]), .out(far_7_7686_1[1]));
    assign out[546] = far_7_7686_1[1] & ~far_7_7686_1[0]; 
    wire [1:0] far_7_7687_0;    relay_conn far_7_7687_0_a(.in(layer_6[456]), .out(far_7_7687_0[0]));    relay_conn far_7_7687_0_b(.in(layer_6[512]), .out(far_7_7687_0[1]));
    assign out[547] = far_7_7687_0[1]; 
    wire [1:0] far_7_7688_0;    relay_conn far_7_7688_0_a(.in(layer_6[197]), .out(far_7_7688_0[0]));    relay_conn far_7_7688_0_b(.in(layer_6[109]), .out(far_7_7688_0[1]));
    wire [1:0] far_7_7688_1;    relay_conn far_7_7688_1_a(.in(far_7_7688_0[0]), .out(far_7_7688_1[0]));    relay_conn far_7_7688_1_b(.in(far_7_7688_0[1]), .out(far_7_7688_1[1]));
    assign out[548] = ~(far_7_7688_1[0] | far_7_7688_1[1]); 
    wire [1:0] far_7_7689_0;    relay_conn far_7_7689_0_a(.in(layer_6[318]), .out(far_7_7689_0[0]));    relay_conn far_7_7689_0_b(.in(layer_6[253]), .out(far_7_7689_0[1]));
    wire [1:0] far_7_7689_1;    relay_conn far_7_7689_1_a(.in(far_7_7689_0[0]), .out(far_7_7689_1[0]));    relay_conn far_7_7689_1_b(.in(far_7_7689_0[1]), .out(far_7_7689_1[1]));
    assign out[549] = far_7_7689_1[0] & far_7_7689_1[1]; 
    wire [1:0] far_7_7690_0;    relay_conn far_7_7690_0_a(.in(layer_6[182]), .out(far_7_7690_0[0]));    relay_conn far_7_7690_0_b(.in(layer_6[100]), .out(far_7_7690_0[1]));
    wire [1:0] far_7_7690_1;    relay_conn far_7_7690_1_a(.in(far_7_7690_0[0]), .out(far_7_7690_1[0]));    relay_conn far_7_7690_1_b(.in(far_7_7690_0[1]), .out(far_7_7690_1[1]));
    assign out[550] = far_7_7690_1[0]; 
    wire [1:0] far_7_7691_0;    relay_conn far_7_7691_0_a(.in(layer_6[557]), .out(far_7_7691_0[0]));    relay_conn far_7_7691_0_b(.in(layer_6[596]), .out(far_7_7691_0[1]));
    assign out[551] = ~(far_7_7691_0[0] ^ far_7_7691_0[1]); 
    assign out[552] = layer_6[920] & ~layer_6[910]; 
    assign out[553] = layer_6[950] & ~layer_6[981]; 
    wire [1:0] far_7_7694_0;    relay_conn far_7_7694_0_a(.in(layer_6[208]), .out(far_7_7694_0[0]));    relay_conn far_7_7694_0_b(.in(layer_6[175]), .out(far_7_7694_0[1]));
    assign out[554] = far_7_7694_0[0] & far_7_7694_0[1]; 
    wire [1:0] far_7_7695_0;    relay_conn far_7_7695_0_a(.in(layer_6[356]), .out(far_7_7695_0[0]));    relay_conn far_7_7695_0_b(.in(layer_6[254]), .out(far_7_7695_0[1]));
    wire [1:0] far_7_7695_1;    relay_conn far_7_7695_1_a(.in(far_7_7695_0[0]), .out(far_7_7695_1[0]));    relay_conn far_7_7695_1_b(.in(far_7_7695_0[1]), .out(far_7_7695_1[1]));
    wire [1:0] far_7_7695_2;    relay_conn far_7_7695_2_a(.in(far_7_7695_1[0]), .out(far_7_7695_2[0]));    relay_conn far_7_7695_2_b(.in(far_7_7695_1[1]), .out(far_7_7695_2[1]));
    assign out[555] = far_7_7695_2[0] & ~far_7_7695_2[1]; 
    wire [1:0] far_7_7696_0;    relay_conn far_7_7696_0_a(.in(layer_6[620]), .out(far_7_7696_0[0]));    relay_conn far_7_7696_0_b(.in(layer_6[729]), .out(far_7_7696_0[1]));
    wire [1:0] far_7_7696_1;    relay_conn far_7_7696_1_a(.in(far_7_7696_0[0]), .out(far_7_7696_1[0]));    relay_conn far_7_7696_1_b(.in(far_7_7696_0[1]), .out(far_7_7696_1[1]));
    wire [1:0] far_7_7696_2;    relay_conn far_7_7696_2_a(.in(far_7_7696_1[0]), .out(far_7_7696_2[0]));    relay_conn far_7_7696_2_b(.in(far_7_7696_1[1]), .out(far_7_7696_2[1]));
    assign out[556] = ~far_7_7696_2[1]; 
    wire [1:0] far_7_7697_0;    relay_conn far_7_7697_0_a(.in(layer_6[913]), .out(far_7_7697_0[0]));    relay_conn far_7_7697_0_b(.in(layer_6[811]), .out(far_7_7697_0[1]));
    wire [1:0] far_7_7697_1;    relay_conn far_7_7697_1_a(.in(far_7_7697_0[0]), .out(far_7_7697_1[0]));    relay_conn far_7_7697_1_b(.in(far_7_7697_0[1]), .out(far_7_7697_1[1]));
    wire [1:0] far_7_7697_2;    relay_conn far_7_7697_2_a(.in(far_7_7697_1[0]), .out(far_7_7697_2[0]));    relay_conn far_7_7697_2_b(.in(far_7_7697_1[1]), .out(far_7_7697_2[1]));
    assign out[557] = ~far_7_7697_2[1]; 
    wire [1:0] far_7_7698_0;    relay_conn far_7_7698_0_a(.in(layer_6[478]), .out(far_7_7698_0[0]));    relay_conn far_7_7698_0_b(.in(layer_6[563]), .out(far_7_7698_0[1]));
    wire [1:0] far_7_7698_1;    relay_conn far_7_7698_1_a(.in(far_7_7698_0[0]), .out(far_7_7698_1[0]));    relay_conn far_7_7698_1_b(.in(far_7_7698_0[1]), .out(far_7_7698_1[1]));
    assign out[558] = ~(far_7_7698_1[0] | far_7_7698_1[1]); 
    wire [1:0] far_7_7699_0;    relay_conn far_7_7699_0_a(.in(layer_6[705]), .out(far_7_7699_0[0]));    relay_conn far_7_7699_0_b(.in(layer_6[615]), .out(far_7_7699_0[1]));
    wire [1:0] far_7_7699_1;    relay_conn far_7_7699_1_a(.in(far_7_7699_0[0]), .out(far_7_7699_1[0]));    relay_conn far_7_7699_1_b(.in(far_7_7699_0[1]), .out(far_7_7699_1[1]));
    assign out[559] = far_7_7699_1[1]; 
    wire [1:0] far_7_7700_0;    relay_conn far_7_7700_0_a(.in(layer_6[376]), .out(far_7_7700_0[0]));    relay_conn far_7_7700_0_b(.in(layer_6[498]), .out(far_7_7700_0[1]));
    wire [1:0] far_7_7700_1;    relay_conn far_7_7700_1_a(.in(far_7_7700_0[0]), .out(far_7_7700_1[0]));    relay_conn far_7_7700_1_b(.in(far_7_7700_0[1]), .out(far_7_7700_1[1]));
    wire [1:0] far_7_7700_2;    relay_conn far_7_7700_2_a(.in(far_7_7700_1[0]), .out(far_7_7700_2[0]));    relay_conn far_7_7700_2_b(.in(far_7_7700_1[1]), .out(far_7_7700_2[1]));
    assign out[560] = far_7_7700_2[0] & far_7_7700_2[1]; 
    wire [1:0] far_7_7701_0;    relay_conn far_7_7701_0_a(.in(layer_6[397]), .out(far_7_7701_0[0]));    relay_conn far_7_7701_0_b(.in(layer_6[307]), .out(far_7_7701_0[1]));
    wire [1:0] far_7_7701_1;    relay_conn far_7_7701_1_a(.in(far_7_7701_0[0]), .out(far_7_7701_1[0]));    relay_conn far_7_7701_1_b(.in(far_7_7701_0[1]), .out(far_7_7701_1[1]));
    assign out[561] = far_7_7701_1[1] & ~far_7_7701_1[0]; 
    wire [1:0] far_7_7702_0;    relay_conn far_7_7702_0_a(.in(layer_6[222]), .out(far_7_7702_0[0]));    relay_conn far_7_7702_0_b(.in(layer_6[290]), .out(far_7_7702_0[1]));
    wire [1:0] far_7_7702_1;    relay_conn far_7_7702_1_a(.in(far_7_7702_0[0]), .out(far_7_7702_1[0]));    relay_conn far_7_7702_1_b(.in(far_7_7702_0[1]), .out(far_7_7702_1[1]));
    assign out[562] = ~(far_7_7702_1[0] | far_7_7702_1[1]); 
    wire [1:0] far_7_7703_0;    relay_conn far_7_7703_0_a(.in(layer_6[208]), .out(far_7_7703_0[0]));    relay_conn far_7_7703_0_b(.in(layer_6[315]), .out(far_7_7703_0[1]));
    wire [1:0] far_7_7703_1;    relay_conn far_7_7703_1_a(.in(far_7_7703_0[0]), .out(far_7_7703_1[0]));    relay_conn far_7_7703_1_b(.in(far_7_7703_0[1]), .out(far_7_7703_1[1]));
    wire [1:0] far_7_7703_2;    relay_conn far_7_7703_2_a(.in(far_7_7703_1[0]), .out(far_7_7703_2[0]));    relay_conn far_7_7703_2_b(.in(far_7_7703_1[1]), .out(far_7_7703_2[1]));
    assign out[563] = far_7_7703_2[0]; 
    wire [1:0] far_7_7704_0;    relay_conn far_7_7704_0_a(.in(layer_6[732]), .out(far_7_7704_0[0]));    relay_conn far_7_7704_0_b(.in(layer_6[659]), .out(far_7_7704_0[1]));
    wire [1:0] far_7_7704_1;    relay_conn far_7_7704_1_a(.in(far_7_7704_0[0]), .out(far_7_7704_1[0]));    relay_conn far_7_7704_1_b(.in(far_7_7704_0[1]), .out(far_7_7704_1[1]));
    assign out[564] = ~(far_7_7704_1[0] | far_7_7704_1[1]); 
    wire [1:0] far_7_7705_0;    relay_conn far_7_7705_0_a(.in(layer_6[1008]), .out(far_7_7705_0[0]));    relay_conn far_7_7705_0_b(.in(layer_6[881]), .out(far_7_7705_0[1]));
    wire [1:0] far_7_7705_1;    relay_conn far_7_7705_1_a(.in(far_7_7705_0[0]), .out(far_7_7705_1[0]));    relay_conn far_7_7705_1_b(.in(far_7_7705_0[1]), .out(far_7_7705_1[1]));
    wire [1:0] far_7_7705_2;    relay_conn far_7_7705_2_a(.in(far_7_7705_1[0]), .out(far_7_7705_2[0]));    relay_conn far_7_7705_2_b(.in(far_7_7705_1[1]), .out(far_7_7705_2[1]));
    assign out[565] = far_7_7705_2[0]; 
    wire [1:0] far_7_7706_0;    relay_conn far_7_7706_0_a(.in(layer_6[591]), .out(far_7_7706_0[0]));    relay_conn far_7_7706_0_b(.in(layer_6[659]), .out(far_7_7706_0[1]));
    wire [1:0] far_7_7706_1;    relay_conn far_7_7706_1_a(.in(far_7_7706_0[0]), .out(far_7_7706_1[0]));    relay_conn far_7_7706_1_b(.in(far_7_7706_0[1]), .out(far_7_7706_1[1]));
    assign out[566] = far_7_7706_1[0] & ~far_7_7706_1[1]; 
    assign out[567] = ~(layer_6[271] | layer_6[299]); 
    wire [1:0] far_7_7708_0;    relay_conn far_7_7708_0_a(.in(layer_6[128]), .out(far_7_7708_0[0]));    relay_conn far_7_7708_0_b(.in(layer_6[181]), .out(far_7_7708_0[1]));
    assign out[568] = far_7_7708_0[0] & far_7_7708_0[1]; 
    wire [1:0] far_7_7709_0;    relay_conn far_7_7709_0_a(.in(layer_6[649]), .out(far_7_7709_0[0]));    relay_conn far_7_7709_0_b(.in(layer_6[539]), .out(far_7_7709_0[1]));
    wire [1:0] far_7_7709_1;    relay_conn far_7_7709_1_a(.in(far_7_7709_0[0]), .out(far_7_7709_1[0]));    relay_conn far_7_7709_1_b(.in(far_7_7709_0[1]), .out(far_7_7709_1[1]));
    wire [1:0] far_7_7709_2;    relay_conn far_7_7709_2_a(.in(far_7_7709_1[0]), .out(far_7_7709_2[0]));    relay_conn far_7_7709_2_b(.in(far_7_7709_1[1]), .out(far_7_7709_2[1]));
    assign out[569] = far_7_7709_2[0] & ~far_7_7709_2[1]; 
    wire [1:0] far_7_7710_0;    relay_conn far_7_7710_0_a(.in(layer_6[565]), .out(far_7_7710_0[0]));    relay_conn far_7_7710_0_b(.in(layer_6[471]), .out(far_7_7710_0[1]));
    wire [1:0] far_7_7710_1;    relay_conn far_7_7710_1_a(.in(far_7_7710_0[0]), .out(far_7_7710_1[0]));    relay_conn far_7_7710_1_b(.in(far_7_7710_0[1]), .out(far_7_7710_1[1]));
    assign out[570] = ~(far_7_7710_1[0] | far_7_7710_1[1]); 
    assign out[571] = layer_6[455]; 
    assign out[572] = layer_6[150]; 
    wire [1:0] far_7_7713_0;    relay_conn far_7_7713_0_a(.in(layer_6[773]), .out(far_7_7713_0[0]));    relay_conn far_7_7713_0_b(.in(layer_6[718]), .out(far_7_7713_0[1]));
    assign out[573] = ~(far_7_7713_0[0] | far_7_7713_0[1]); 
    assign out[574] = layer_6[573] & ~layer_6[550]; 
    wire [1:0] far_7_7715_0;    relay_conn far_7_7715_0_a(.in(layer_6[966]), .out(far_7_7715_0[0]));    relay_conn far_7_7715_0_b(.in(layer_6[1008]), .out(far_7_7715_0[1]));
    assign out[575] = far_7_7715_0[0] & far_7_7715_0[1]; 
    assign out[576] = layer_6[932]; 
    assign out[577] = ~(layer_6[744] | layer_6[767]); 
    wire [1:0] far_7_7718_0;    relay_conn far_7_7718_0_a(.in(layer_6[29]), .out(far_7_7718_0[0]));    relay_conn far_7_7718_0_b(.in(layer_6[124]), .out(far_7_7718_0[1]));
    wire [1:0] far_7_7718_1;    relay_conn far_7_7718_1_a(.in(far_7_7718_0[0]), .out(far_7_7718_1[0]));    relay_conn far_7_7718_1_b(.in(far_7_7718_0[1]), .out(far_7_7718_1[1]));
    assign out[578] = far_7_7718_1[0]; 
    wire [1:0] far_7_7719_0;    relay_conn far_7_7719_0_a(.in(layer_6[261]), .out(far_7_7719_0[0]));    relay_conn far_7_7719_0_b(.in(layer_6[350]), .out(far_7_7719_0[1]));
    wire [1:0] far_7_7719_1;    relay_conn far_7_7719_1_a(.in(far_7_7719_0[0]), .out(far_7_7719_1[0]));    relay_conn far_7_7719_1_b(.in(far_7_7719_0[1]), .out(far_7_7719_1[1]));
    assign out[579] = far_7_7719_1[1] & ~far_7_7719_1[0]; 
    assign out[580] = ~layer_6[913] | (layer_6[913] & layer_6[917]); 
    wire [1:0] far_7_7721_0;    relay_conn far_7_7721_0_a(.in(layer_6[361]), .out(far_7_7721_0[0]));    relay_conn far_7_7721_0_b(.in(layer_6[437]), .out(far_7_7721_0[1]));
    wire [1:0] far_7_7721_1;    relay_conn far_7_7721_1_a(.in(far_7_7721_0[0]), .out(far_7_7721_1[0]));    relay_conn far_7_7721_1_b(.in(far_7_7721_0[1]), .out(far_7_7721_1[1]));
    assign out[581] = far_7_7721_1[0] & far_7_7721_1[1]; 
    wire [1:0] far_7_7722_0;    relay_conn far_7_7722_0_a(.in(layer_6[60]), .out(far_7_7722_0[0]));    relay_conn far_7_7722_0_b(.in(layer_6[119]), .out(far_7_7722_0[1]));
    assign out[582] = ~far_7_7722_0[0]; 
    assign out[583] = layer_6[966] & ~layer_6[994]; 
    assign out[584] = layer_6[742] & ~layer_6[763]; 
    assign out[585] = layer_6[393] & layer_6[394]; 
    assign out[586] = ~(layer_6[647] | layer_6[656]); 
    assign out[587] = layer_6[485] & ~layer_6[510]; 
    assign out[588] = layer_6[788] & ~layer_6[799]; 
    assign out[589] = layer_6[37] & ~layer_6[60]; 
    wire [1:0] far_7_7730_0;    relay_conn far_7_7730_0_a(.in(layer_6[42]), .out(far_7_7730_0[0]));    relay_conn far_7_7730_0_b(.in(layer_6[97]), .out(far_7_7730_0[1]));
    assign out[590] = far_7_7730_0[1]; 
    wire [1:0] far_7_7731_0;    relay_conn far_7_7731_0_a(.in(layer_6[571]), .out(far_7_7731_0[0]));    relay_conn far_7_7731_0_b(.in(layer_6[632]), .out(far_7_7731_0[1]));
    assign out[591] = ~far_7_7731_0[0]; 
    wire [1:0] far_7_7732_0;    relay_conn far_7_7732_0_a(.in(layer_6[543]), .out(far_7_7732_0[0]));    relay_conn far_7_7732_0_b(.in(layer_6[475]), .out(far_7_7732_0[1]));
    wire [1:0] far_7_7732_1;    relay_conn far_7_7732_1_a(.in(far_7_7732_0[0]), .out(far_7_7732_1[0]));    relay_conn far_7_7732_1_b(.in(far_7_7732_0[1]), .out(far_7_7732_1[1]));
    assign out[592] = far_7_7732_1[0] & far_7_7732_1[1]; 
    assign out[593] = ~layer_6[755]; 
    assign out[594] = layer_6[470] & layer_6[460]; 
    assign out[595] = ~layer_6[404]; 
    assign out[596] = layer_6[742] & ~layer_6[763]; 
    wire [1:0] far_7_7737_0;    relay_conn far_7_7737_0_a(.in(layer_6[416]), .out(far_7_7737_0[0]));    relay_conn far_7_7737_0_b(.in(layer_6[491]), .out(far_7_7737_0[1]));
    wire [1:0] far_7_7737_1;    relay_conn far_7_7737_1_a(.in(far_7_7737_0[0]), .out(far_7_7737_1[0]));    relay_conn far_7_7737_1_b(.in(far_7_7737_0[1]), .out(far_7_7737_1[1]));
    assign out[597] = ~(far_7_7737_1[0] ^ far_7_7737_1[1]); 
    wire [1:0] far_7_7738_0;    relay_conn far_7_7738_0_a(.in(layer_6[372]), .out(far_7_7738_0[0]));    relay_conn far_7_7738_0_b(.in(layer_6[329]), .out(far_7_7738_0[1]));
    assign out[598] = far_7_7738_0[0] & far_7_7738_0[1]; 
    wire [1:0] far_7_7739_0;    relay_conn far_7_7739_0_a(.in(layer_6[569]), .out(far_7_7739_0[0]));    relay_conn far_7_7739_0_b(.in(layer_6[602]), .out(far_7_7739_0[1]));
    assign out[599] = far_7_7739_0[0] & far_7_7739_0[1]; 
    wire [1:0] far_7_7740_0;    relay_conn far_7_7740_0_a(.in(layer_6[400]), .out(far_7_7740_0[0]));    relay_conn far_7_7740_0_b(.in(layer_6[476]), .out(far_7_7740_0[1]));
    wire [1:0] far_7_7740_1;    relay_conn far_7_7740_1_a(.in(far_7_7740_0[0]), .out(far_7_7740_1[0]));    relay_conn far_7_7740_1_b(.in(far_7_7740_0[1]), .out(far_7_7740_1[1]));
    assign out[600] = far_7_7740_1[0] & ~far_7_7740_1[1]; 
    wire [1:0] far_7_7741_0;    relay_conn far_7_7741_0_a(.in(layer_6[981]), .out(far_7_7741_0[0]));    relay_conn far_7_7741_0_b(.in(layer_6[919]), .out(far_7_7741_0[1]));
    assign out[601] = far_7_7741_0[1] & ~far_7_7741_0[0]; 
    wire [1:0] far_7_7742_0;    relay_conn far_7_7742_0_a(.in(layer_6[342]), .out(far_7_7742_0[0]));    relay_conn far_7_7742_0_b(.in(layer_6[404]), .out(far_7_7742_0[1]));
    assign out[602] = ~far_7_7742_0[1]; 
    assign out[603] = ~(layer_6[404] & layer_6[412]); 
    wire [1:0] far_7_7744_0;    relay_conn far_7_7744_0_a(.in(layer_6[481]), .out(far_7_7744_0[0]));    relay_conn far_7_7744_0_b(.in(layer_6[449]), .out(far_7_7744_0[1]));
    assign out[604] = ~far_7_7744_0[0] | (far_7_7744_0[0] & far_7_7744_0[1]); 
    assign out[605] = layer_6[731]; 
    assign out[606] = layer_6[490]; 
    wire [1:0] far_7_7747_0;    relay_conn far_7_7747_0_a(.in(layer_6[924]), .out(far_7_7747_0[0]));    relay_conn far_7_7747_0_b(.in(layer_6[990]), .out(far_7_7747_0[1]));
    wire [1:0] far_7_7747_1;    relay_conn far_7_7747_1_a(.in(far_7_7747_0[0]), .out(far_7_7747_1[0]));    relay_conn far_7_7747_1_b(.in(far_7_7747_0[1]), .out(far_7_7747_1[1]));
    assign out[607] = ~far_7_7747_1[1]; 
    wire [1:0] far_7_7748_0;    relay_conn far_7_7748_0_a(.in(layer_6[210]), .out(far_7_7748_0[0]));    relay_conn far_7_7748_0_b(.in(layer_6[96]), .out(far_7_7748_0[1]));
    wire [1:0] far_7_7748_1;    relay_conn far_7_7748_1_a(.in(far_7_7748_0[0]), .out(far_7_7748_1[0]));    relay_conn far_7_7748_1_b(.in(far_7_7748_0[1]), .out(far_7_7748_1[1]));
    wire [1:0] far_7_7748_2;    relay_conn far_7_7748_2_a(.in(far_7_7748_1[0]), .out(far_7_7748_2[0]));    relay_conn far_7_7748_2_b(.in(far_7_7748_1[1]), .out(far_7_7748_2[1]));
    assign out[608] = ~(far_7_7748_2[0] | far_7_7748_2[1]); 
    assign out[609] = layer_6[240]; 
    wire [1:0] far_7_7750_0;    relay_conn far_7_7750_0_a(.in(layer_6[663]), .out(far_7_7750_0[0]));    relay_conn far_7_7750_0_b(.in(layer_6[737]), .out(far_7_7750_0[1]));
    wire [1:0] far_7_7750_1;    relay_conn far_7_7750_1_a(.in(far_7_7750_0[0]), .out(far_7_7750_1[0]));    relay_conn far_7_7750_1_b(.in(far_7_7750_0[1]), .out(far_7_7750_1[1]));
    assign out[610] = far_7_7750_1[1] & ~far_7_7750_1[0]; 
    assign out[611] = layer_6[970] ^ layer_6[942]; 
    wire [1:0] far_7_7752_0;    relay_conn far_7_7752_0_a(.in(layer_6[908]), .out(far_7_7752_0[0]));    relay_conn far_7_7752_0_b(.in(layer_6[971]), .out(far_7_7752_0[1]));
    assign out[612] = ~(far_7_7752_0[0] & far_7_7752_0[1]); 
    wire [1:0] far_7_7753_0;    relay_conn far_7_7753_0_a(.in(layer_6[306]), .out(far_7_7753_0[0]));    relay_conn far_7_7753_0_b(.in(layer_6[202]), .out(far_7_7753_0[1]));
    wire [1:0] far_7_7753_1;    relay_conn far_7_7753_1_a(.in(far_7_7753_0[0]), .out(far_7_7753_1[0]));    relay_conn far_7_7753_1_b(.in(far_7_7753_0[1]), .out(far_7_7753_1[1]));
    wire [1:0] far_7_7753_2;    relay_conn far_7_7753_2_a(.in(far_7_7753_1[0]), .out(far_7_7753_2[0]));    relay_conn far_7_7753_2_b(.in(far_7_7753_1[1]), .out(far_7_7753_2[1]));
    assign out[613] = far_7_7753_2[0]; 
    wire [1:0] far_7_7754_0;    relay_conn far_7_7754_0_a(.in(layer_6[837]), .out(far_7_7754_0[0]));    relay_conn far_7_7754_0_b(.in(layer_6[737]), .out(far_7_7754_0[1]));
    wire [1:0] far_7_7754_1;    relay_conn far_7_7754_1_a(.in(far_7_7754_0[0]), .out(far_7_7754_1[0]));    relay_conn far_7_7754_1_b(.in(far_7_7754_0[1]), .out(far_7_7754_1[1]));
    wire [1:0] far_7_7754_2;    relay_conn far_7_7754_2_a(.in(far_7_7754_1[0]), .out(far_7_7754_2[0]));    relay_conn far_7_7754_2_b(.in(far_7_7754_1[1]), .out(far_7_7754_2[1]));
    assign out[614] = ~far_7_7754_2[1]; 
    assign out[615] = ~(layer_6[416] ^ layer_6[424]); 
    wire [1:0] far_7_7756_0;    relay_conn far_7_7756_0_a(.in(layer_6[617]), .out(far_7_7756_0[0]));    relay_conn far_7_7756_0_b(.in(layer_6[681]), .out(far_7_7756_0[1]));
    wire [1:0] far_7_7756_1;    relay_conn far_7_7756_1_a(.in(far_7_7756_0[0]), .out(far_7_7756_1[0]));    relay_conn far_7_7756_1_b(.in(far_7_7756_0[1]), .out(far_7_7756_1[1]));
    assign out[616] = far_7_7756_1[1]; 
    wire [1:0] far_7_7757_0;    relay_conn far_7_7757_0_a(.in(layer_6[408]), .out(far_7_7757_0[0]));    relay_conn far_7_7757_0_b(.in(layer_6[511]), .out(far_7_7757_0[1]));
    wire [1:0] far_7_7757_1;    relay_conn far_7_7757_1_a(.in(far_7_7757_0[0]), .out(far_7_7757_1[0]));    relay_conn far_7_7757_1_b(.in(far_7_7757_0[1]), .out(far_7_7757_1[1]));
    wire [1:0] far_7_7757_2;    relay_conn far_7_7757_2_a(.in(far_7_7757_1[0]), .out(far_7_7757_2[0]));    relay_conn far_7_7757_2_b(.in(far_7_7757_1[1]), .out(far_7_7757_2[1]));
    assign out[617] = far_7_7757_2[0]; 
    wire [1:0] far_7_7758_0;    relay_conn far_7_7758_0_a(.in(layer_6[956]), .out(far_7_7758_0[0]));    relay_conn far_7_7758_0_b(.in(layer_6[995]), .out(far_7_7758_0[1]));
    assign out[618] = far_7_7758_0[0] ^ far_7_7758_0[1]; 
    wire [1:0] far_7_7759_0;    relay_conn far_7_7759_0_a(.in(layer_6[56]), .out(far_7_7759_0[0]));    relay_conn far_7_7759_0_b(.in(layer_6[146]), .out(far_7_7759_0[1]));
    wire [1:0] far_7_7759_1;    relay_conn far_7_7759_1_a(.in(far_7_7759_0[0]), .out(far_7_7759_1[0]));    relay_conn far_7_7759_1_b(.in(far_7_7759_0[1]), .out(far_7_7759_1[1]));
    assign out[619] = far_7_7759_1[0] | far_7_7759_1[1]; 
    wire [1:0] far_7_7760_0;    relay_conn far_7_7760_0_a(.in(layer_6[924]), .out(far_7_7760_0[0]));    relay_conn far_7_7760_0_b(.in(layer_6[1015]), .out(far_7_7760_0[1]));
    wire [1:0] far_7_7760_1;    relay_conn far_7_7760_1_a(.in(far_7_7760_0[0]), .out(far_7_7760_1[0]));    relay_conn far_7_7760_1_b(.in(far_7_7760_0[1]), .out(far_7_7760_1[1]));
    assign out[620] = ~(far_7_7760_1[0] ^ far_7_7760_1[1]); 
    wire [1:0] far_7_7761_0;    relay_conn far_7_7761_0_a(.in(layer_6[499]), .out(far_7_7761_0[0]));    relay_conn far_7_7761_0_b(.in(layer_6[424]), .out(far_7_7761_0[1]));
    wire [1:0] far_7_7761_1;    relay_conn far_7_7761_1_a(.in(far_7_7761_0[0]), .out(far_7_7761_1[0]));    relay_conn far_7_7761_1_b(.in(far_7_7761_0[1]), .out(far_7_7761_1[1]));
    assign out[621] = ~(far_7_7761_1[0] ^ far_7_7761_1[1]); 
    wire [1:0] far_7_7762_0;    relay_conn far_7_7762_0_a(.in(layer_6[491]), .out(far_7_7762_0[0]));    relay_conn far_7_7762_0_b(.in(layer_6[396]), .out(far_7_7762_0[1]));
    wire [1:0] far_7_7762_1;    relay_conn far_7_7762_1_a(.in(far_7_7762_0[0]), .out(far_7_7762_1[0]));    relay_conn far_7_7762_1_b(.in(far_7_7762_0[1]), .out(far_7_7762_1[1]));
    assign out[622] = ~(far_7_7762_1[0] ^ far_7_7762_1[1]); 
    wire [1:0] far_7_7763_0;    relay_conn far_7_7763_0_a(.in(layer_6[629]), .out(far_7_7763_0[0]));    relay_conn far_7_7763_0_b(.in(layer_6[539]), .out(far_7_7763_0[1]));
    wire [1:0] far_7_7763_1;    relay_conn far_7_7763_1_a(.in(far_7_7763_0[0]), .out(far_7_7763_1[0]));    relay_conn far_7_7763_1_b(.in(far_7_7763_0[1]), .out(far_7_7763_1[1]));
    assign out[623] = ~(far_7_7763_1[0] | far_7_7763_1[1]); 
    assign out[624] = layer_6[779] & ~layer_6[759]; 
    assign out[625] = ~(layer_6[867] ^ layer_6[874]); 
    wire [1:0] far_7_7766_0;    relay_conn far_7_7766_0_a(.in(layer_6[273]), .out(far_7_7766_0[0]));    relay_conn far_7_7766_0_b(.in(layer_6[310]), .out(far_7_7766_0[1]));
    assign out[626] = far_7_7766_0[0] & far_7_7766_0[1]; 
    wire [1:0] far_7_7767_0;    relay_conn far_7_7767_0_a(.in(layer_6[871]), .out(far_7_7767_0[0]));    relay_conn far_7_7767_0_b(.in(layer_6[822]), .out(far_7_7767_0[1]));
    assign out[627] = ~(far_7_7767_0[0] ^ far_7_7767_0[1]); 
    wire [1:0] far_7_7768_0;    relay_conn far_7_7768_0_a(.in(layer_6[996]), .out(far_7_7768_0[0]));    relay_conn far_7_7768_0_b(.in(layer_6[919]), .out(far_7_7768_0[1]));
    wire [1:0] far_7_7768_1;    relay_conn far_7_7768_1_a(.in(far_7_7768_0[0]), .out(far_7_7768_1[0]));    relay_conn far_7_7768_1_b(.in(far_7_7768_0[1]), .out(far_7_7768_1[1]));
    assign out[628] = far_7_7768_1[0]; 
    wire [1:0] far_7_7769_0;    relay_conn far_7_7769_0_a(.in(layer_6[451]), .out(far_7_7769_0[0]));    relay_conn far_7_7769_0_b(.in(layer_6[338]), .out(far_7_7769_0[1]));
    wire [1:0] far_7_7769_1;    relay_conn far_7_7769_1_a(.in(far_7_7769_0[0]), .out(far_7_7769_1[0]));    relay_conn far_7_7769_1_b(.in(far_7_7769_0[1]), .out(far_7_7769_1[1]));
    wire [1:0] far_7_7769_2;    relay_conn far_7_7769_2_a(.in(far_7_7769_1[0]), .out(far_7_7769_2[0]));    relay_conn far_7_7769_2_b(.in(far_7_7769_1[1]), .out(far_7_7769_2[1]));
    assign out[629] = ~(far_7_7769_2[0] | far_7_7769_2[1]); 
    assign out[630] = ~layer_6[687]; 
    wire [1:0] far_7_7771_0;    relay_conn far_7_7771_0_a(.in(layer_6[557]), .out(far_7_7771_0[0]));    relay_conn far_7_7771_0_b(.in(layer_6[511]), .out(far_7_7771_0[1]));
    assign out[631] = far_7_7771_0[0] & far_7_7771_0[1]; 
    assign out[632] = layer_6[475] & ~layer_6[497]; 
    wire [1:0] far_7_7773_0;    relay_conn far_7_7773_0_a(.in(layer_6[672]), .out(far_7_7773_0[0]));    relay_conn far_7_7773_0_b(.in(layer_6[737]), .out(far_7_7773_0[1]));
    wire [1:0] far_7_7773_1;    relay_conn far_7_7773_1_a(.in(far_7_7773_0[0]), .out(far_7_7773_1[0]));    relay_conn far_7_7773_1_b(.in(far_7_7773_0[1]), .out(far_7_7773_1[1]));
    assign out[633] = ~far_7_7773_1[1]; 
    wire [1:0] far_7_7774_0;    relay_conn far_7_7774_0_a(.in(layer_6[229]), .out(far_7_7774_0[0]));    relay_conn far_7_7774_0_b(.in(layer_6[197]), .out(far_7_7774_0[1]));
    assign out[634] = ~far_7_7774_0[0]; 
    assign out[635] = layer_6[648]; 
    wire [1:0] far_7_7776_0;    relay_conn far_7_7776_0_a(.in(layer_6[416]), .out(far_7_7776_0[0]));    relay_conn far_7_7776_0_b(.in(layer_6[324]), .out(far_7_7776_0[1]));
    wire [1:0] far_7_7776_1;    relay_conn far_7_7776_1_a(.in(far_7_7776_0[0]), .out(far_7_7776_1[0]));    relay_conn far_7_7776_1_b(.in(far_7_7776_0[1]), .out(far_7_7776_1[1]));
    assign out[636] = ~far_7_7776_1[1]; 
    wire [1:0] far_7_7777_0;    relay_conn far_7_7777_0_a(.in(layer_6[845]), .out(far_7_7777_0[0]));    relay_conn far_7_7777_0_b(.in(layer_6[730]), .out(far_7_7777_0[1]));
    wire [1:0] far_7_7777_1;    relay_conn far_7_7777_1_a(.in(far_7_7777_0[0]), .out(far_7_7777_1[0]));    relay_conn far_7_7777_1_b(.in(far_7_7777_0[1]), .out(far_7_7777_1[1]));
    wire [1:0] far_7_7777_2;    relay_conn far_7_7777_2_a(.in(far_7_7777_1[0]), .out(far_7_7777_2[0]));    relay_conn far_7_7777_2_b(.in(far_7_7777_1[1]), .out(far_7_7777_2[1]));
    assign out[637] = ~far_7_7777_2[0] | (far_7_7777_2[0] & far_7_7777_2[1]); 
    wire [1:0] far_7_7778_0;    relay_conn far_7_7778_0_a(.in(layer_6[775]), .out(far_7_7778_0[0]));    relay_conn far_7_7778_0_b(.in(layer_6[681]), .out(far_7_7778_0[1]));
    wire [1:0] far_7_7778_1;    relay_conn far_7_7778_1_a(.in(far_7_7778_0[0]), .out(far_7_7778_1[0]));    relay_conn far_7_7778_1_b(.in(far_7_7778_0[1]), .out(far_7_7778_1[1]));
    assign out[638] = far_7_7778_1[1]; 
    wire [1:0] far_7_7779_0;    relay_conn far_7_7779_0_a(.in(layer_6[404]), .out(far_7_7779_0[0]));    relay_conn far_7_7779_0_b(.in(layer_6[476]), .out(far_7_7779_0[1]));
    wire [1:0] far_7_7779_1;    relay_conn far_7_7779_1_a(.in(far_7_7779_0[0]), .out(far_7_7779_1[0]));    relay_conn far_7_7779_1_b(.in(far_7_7779_0[1]), .out(far_7_7779_1[1]));
    assign out[639] = far_7_7779_1[0] & far_7_7779_1[1]; 
    wire [1:0] far_7_7780_0;    relay_conn far_7_7780_0_a(.in(layer_6[306]), .out(far_7_7780_0[0]));    relay_conn far_7_7780_0_b(.in(layer_6[203]), .out(far_7_7780_0[1]));
    wire [1:0] far_7_7780_1;    relay_conn far_7_7780_1_a(.in(far_7_7780_0[0]), .out(far_7_7780_1[0]));    relay_conn far_7_7780_1_b(.in(far_7_7780_0[1]), .out(far_7_7780_1[1]));
    wire [1:0] far_7_7780_2;    relay_conn far_7_7780_2_a(.in(far_7_7780_1[0]), .out(far_7_7780_2[0]));    relay_conn far_7_7780_2_b(.in(far_7_7780_1[1]), .out(far_7_7780_2[1]));
    assign out[640] = far_7_7780_2[0]; 
    assign out[641] = layer_6[646] & layer_6[615]; 
    wire [1:0] far_7_7782_0;    relay_conn far_7_7782_0_a(.in(layer_6[237]), .out(far_7_7782_0[0]));    relay_conn far_7_7782_0_b(.in(layer_6[139]), .out(far_7_7782_0[1]));
    wire [1:0] far_7_7782_1;    relay_conn far_7_7782_1_a(.in(far_7_7782_0[0]), .out(far_7_7782_1[0]));    relay_conn far_7_7782_1_b(.in(far_7_7782_0[1]), .out(far_7_7782_1[1]));
    wire [1:0] far_7_7782_2;    relay_conn far_7_7782_2_a(.in(far_7_7782_1[0]), .out(far_7_7782_2[0]));    relay_conn far_7_7782_2_b(.in(far_7_7782_1[1]), .out(far_7_7782_2[1]));
    assign out[642] = ~(far_7_7782_2[0] | far_7_7782_2[1]); 
    assign out[643] = layer_6[919] & ~layer_6[950]; 
    wire [1:0] far_7_7784_0;    relay_conn far_7_7784_0_a(.in(layer_6[799]), .out(far_7_7784_0[0]));    relay_conn far_7_7784_0_b(.in(layer_6[676]), .out(far_7_7784_0[1]));
    wire [1:0] far_7_7784_1;    relay_conn far_7_7784_1_a(.in(far_7_7784_0[0]), .out(far_7_7784_1[0]));    relay_conn far_7_7784_1_b(.in(far_7_7784_0[1]), .out(far_7_7784_1[1]));
    wire [1:0] far_7_7784_2;    relay_conn far_7_7784_2_a(.in(far_7_7784_1[0]), .out(far_7_7784_2[0]));    relay_conn far_7_7784_2_b(.in(far_7_7784_1[1]), .out(far_7_7784_2[1]));
    assign out[644] = far_7_7784_2[0] & ~far_7_7784_2[1]; 
    wire [1:0] far_7_7785_0;    relay_conn far_7_7785_0_a(.in(layer_6[931]), .out(far_7_7785_0[0]));    relay_conn far_7_7785_0_b(.in(layer_6[888]), .out(far_7_7785_0[1]));
    assign out[645] = far_7_7785_0[1] & ~far_7_7785_0[0]; 
    assign out[646] = layer_6[116]; 
    wire [1:0] far_7_7787_0;    relay_conn far_7_7787_0_a(.in(layer_6[100]), .out(far_7_7787_0[0]));    relay_conn far_7_7787_0_b(.in(layer_6[141]), .out(far_7_7787_0[1]));
    assign out[647] = far_7_7787_0[0]; 
    wire [1:0] far_7_7788_0;    relay_conn far_7_7788_0_a(.in(layer_6[580]), .out(far_7_7788_0[0]));    relay_conn far_7_7788_0_b(.in(layer_6[685]), .out(far_7_7788_0[1]));
    wire [1:0] far_7_7788_1;    relay_conn far_7_7788_1_a(.in(far_7_7788_0[0]), .out(far_7_7788_1[0]));    relay_conn far_7_7788_1_b(.in(far_7_7788_0[1]), .out(far_7_7788_1[1]));
    wire [1:0] far_7_7788_2;    relay_conn far_7_7788_2_a(.in(far_7_7788_1[0]), .out(far_7_7788_2[0]));    relay_conn far_7_7788_2_b(.in(far_7_7788_1[1]), .out(far_7_7788_2[1]));
    assign out[648] = far_7_7788_2[0] ^ far_7_7788_2[1]; 
    wire [1:0] far_7_7789_0;    relay_conn far_7_7789_0_a(.in(layer_6[763]), .out(far_7_7789_0[0]));    relay_conn far_7_7789_0_b(.in(layer_6[649]), .out(far_7_7789_0[1]));
    wire [1:0] far_7_7789_1;    relay_conn far_7_7789_1_a(.in(far_7_7789_0[0]), .out(far_7_7789_1[0]));    relay_conn far_7_7789_1_b(.in(far_7_7789_0[1]), .out(far_7_7789_1[1]));
    wire [1:0] far_7_7789_2;    relay_conn far_7_7789_2_a(.in(far_7_7789_1[0]), .out(far_7_7789_2[0]));    relay_conn far_7_7789_2_b(.in(far_7_7789_1[1]), .out(far_7_7789_2[1]));
    assign out[649] = far_7_7789_2[0] ^ far_7_7789_2[1]; 
    wire [1:0] far_7_7790_0;    relay_conn far_7_7790_0_a(.in(layer_6[268]), .out(far_7_7790_0[0]));    relay_conn far_7_7790_0_b(.in(layer_6[186]), .out(far_7_7790_0[1]));
    wire [1:0] far_7_7790_1;    relay_conn far_7_7790_1_a(.in(far_7_7790_0[0]), .out(far_7_7790_1[0]));    relay_conn far_7_7790_1_b(.in(far_7_7790_0[1]), .out(far_7_7790_1[1]));
    assign out[650] = far_7_7790_1[0] & far_7_7790_1[1]; 
    wire [1:0] far_7_7791_0;    relay_conn far_7_7791_0_a(.in(layer_6[435]), .out(far_7_7791_0[0]));    relay_conn far_7_7791_0_b(.in(layer_6[315]), .out(far_7_7791_0[1]));
    wire [1:0] far_7_7791_1;    relay_conn far_7_7791_1_a(.in(far_7_7791_0[0]), .out(far_7_7791_1[0]));    relay_conn far_7_7791_1_b(.in(far_7_7791_0[1]), .out(far_7_7791_1[1]));
    wire [1:0] far_7_7791_2;    relay_conn far_7_7791_2_a(.in(far_7_7791_1[0]), .out(far_7_7791_2[0]));    relay_conn far_7_7791_2_b(.in(far_7_7791_1[1]), .out(far_7_7791_2[1]));
    assign out[651] = ~far_7_7791_2[0]; 
    assign out[652] = layer_6[765] & ~layer_6[760]; 
    wire [1:0] far_7_7793_0;    relay_conn far_7_7793_0_a(.in(layer_6[220]), .out(far_7_7793_0[0]));    relay_conn far_7_7793_0_b(.in(layer_6[339]), .out(far_7_7793_0[1]));
    wire [1:0] far_7_7793_1;    relay_conn far_7_7793_1_a(.in(far_7_7793_0[0]), .out(far_7_7793_1[0]));    relay_conn far_7_7793_1_b(.in(far_7_7793_0[1]), .out(far_7_7793_1[1]));
    wire [1:0] far_7_7793_2;    relay_conn far_7_7793_2_a(.in(far_7_7793_1[0]), .out(far_7_7793_2[0]));    relay_conn far_7_7793_2_b(.in(far_7_7793_1[1]), .out(far_7_7793_2[1]));
    assign out[653] = ~(far_7_7793_2[0] | far_7_7793_2[1]); 
    assign out[654] = layer_6[897] & ~layer_6[866]; 
    wire [1:0] far_7_7795_0;    relay_conn far_7_7795_0_a(.in(layer_6[190]), .out(far_7_7795_0[0]));    relay_conn far_7_7795_0_b(.in(layer_6[297]), .out(far_7_7795_0[1]));
    wire [1:0] far_7_7795_1;    relay_conn far_7_7795_1_a(.in(far_7_7795_0[0]), .out(far_7_7795_1[0]));    relay_conn far_7_7795_1_b(.in(far_7_7795_0[1]), .out(far_7_7795_1[1]));
    wire [1:0] far_7_7795_2;    relay_conn far_7_7795_2_a(.in(far_7_7795_1[0]), .out(far_7_7795_2[0]));    relay_conn far_7_7795_2_b(.in(far_7_7795_1[1]), .out(far_7_7795_2[1]));
    assign out[655] = ~far_7_7795_2[0]; 
    assign out[656] = ~(layer_6[310] ^ layer_6[317]); 
    assign out[657] = layer_6[94] & layer_6[67]; 
    wire [1:0] far_7_7798_0;    relay_conn far_7_7798_0_a(.in(layer_6[663]), .out(far_7_7798_0[0]));    relay_conn far_7_7798_0_b(.in(layer_6[614]), .out(far_7_7798_0[1]));
    assign out[658] = ~far_7_7798_0[1]; 
    wire [1:0] far_7_7799_0;    relay_conn far_7_7799_0_a(.in(layer_6[944]), .out(far_7_7799_0[0]));    relay_conn far_7_7799_0_b(.in(layer_6[860]), .out(far_7_7799_0[1]));
    wire [1:0] far_7_7799_1;    relay_conn far_7_7799_1_a(.in(far_7_7799_0[0]), .out(far_7_7799_1[0]));    relay_conn far_7_7799_1_b(.in(far_7_7799_0[1]), .out(far_7_7799_1[1]));
    assign out[659] = ~far_7_7799_1[1]; 
    wire [1:0] far_7_7800_0;    relay_conn far_7_7800_0_a(.in(layer_6[313]), .out(far_7_7800_0[0]));    relay_conn far_7_7800_0_b(.in(layer_6[418]), .out(far_7_7800_0[1]));
    wire [1:0] far_7_7800_1;    relay_conn far_7_7800_1_a(.in(far_7_7800_0[0]), .out(far_7_7800_1[0]));    relay_conn far_7_7800_1_b(.in(far_7_7800_0[1]), .out(far_7_7800_1[1]));
    wire [1:0] far_7_7800_2;    relay_conn far_7_7800_2_a(.in(far_7_7800_1[0]), .out(far_7_7800_2[0]));    relay_conn far_7_7800_2_b(.in(far_7_7800_1[1]), .out(far_7_7800_2[1]));
    assign out[660] = far_7_7800_2[1] & ~far_7_7800_2[0]; 
    wire [1:0] far_7_7801_0;    relay_conn far_7_7801_0_a(.in(layer_6[100]), .out(far_7_7801_0[0]));    relay_conn far_7_7801_0_b(.in(layer_6[136]), .out(far_7_7801_0[1]));
    assign out[661] = far_7_7801_0[0] & far_7_7801_0[1]; 
    assign out[662] = ~(layer_6[451] | layer_6[472]); 
    assign out[663] = layer_6[489]; 
    wire [1:0] far_7_7804_0;    relay_conn far_7_7804_0_a(.in(layer_6[607]), .out(far_7_7804_0[0]));    relay_conn far_7_7804_0_b(.in(layer_6[541]), .out(far_7_7804_0[1]));
    wire [1:0] far_7_7804_1;    relay_conn far_7_7804_1_a(.in(far_7_7804_0[0]), .out(far_7_7804_1[0]));    relay_conn far_7_7804_1_b(.in(far_7_7804_0[1]), .out(far_7_7804_1[1]));
    assign out[664] = far_7_7804_1[1]; 
    assign out[665] = layer_6[251]; 
    wire [1:0] far_7_7806_0;    relay_conn far_7_7806_0_a(.in(layer_6[230]), .out(far_7_7806_0[0]));    relay_conn far_7_7806_0_b(.in(layer_6[321]), .out(far_7_7806_0[1]));
    wire [1:0] far_7_7806_1;    relay_conn far_7_7806_1_a(.in(far_7_7806_0[0]), .out(far_7_7806_1[0]));    relay_conn far_7_7806_1_b(.in(far_7_7806_0[1]), .out(far_7_7806_1[1]));
    assign out[666] = ~(far_7_7806_1[0] | far_7_7806_1[1]); 
    wire [1:0] far_7_7807_0;    relay_conn far_7_7807_0_a(.in(layer_6[632]), .out(far_7_7807_0[0]));    relay_conn far_7_7807_0_b(.in(layer_6[531]), .out(far_7_7807_0[1]));
    wire [1:0] far_7_7807_1;    relay_conn far_7_7807_1_a(.in(far_7_7807_0[0]), .out(far_7_7807_1[0]));    relay_conn far_7_7807_1_b(.in(far_7_7807_0[1]), .out(far_7_7807_1[1]));
    wire [1:0] far_7_7807_2;    relay_conn far_7_7807_2_a(.in(far_7_7807_1[0]), .out(far_7_7807_2[0]));    relay_conn far_7_7807_2_b(.in(far_7_7807_1[1]), .out(far_7_7807_2[1]));
    assign out[667] = far_7_7807_2[1]; 
    assign out[668] = layer_6[923]; 
    wire [1:0] far_7_7809_0;    relay_conn far_7_7809_0_a(.in(layer_6[228]), .out(far_7_7809_0[0]));    relay_conn far_7_7809_0_b(.in(layer_6[295]), .out(far_7_7809_0[1]));
    wire [1:0] far_7_7809_1;    relay_conn far_7_7809_1_a(.in(far_7_7809_0[0]), .out(far_7_7809_1[0]));    relay_conn far_7_7809_1_b(.in(far_7_7809_0[1]), .out(far_7_7809_1[1]));
    assign out[669] = far_7_7809_1[1]; 
    assign out[670] = ~(layer_6[191] ^ layer_6[165]); 
    assign out[671] = layer_6[155]; 
    assign out[672] = ~layer_6[497]; 
    wire [1:0] far_7_7813_0;    relay_conn far_7_7813_0_a(.in(layer_6[778]), .out(far_7_7813_0[0]));    relay_conn far_7_7813_0_b(.in(layer_6[845]), .out(far_7_7813_0[1]));
    wire [1:0] far_7_7813_1;    relay_conn far_7_7813_1_a(.in(far_7_7813_0[0]), .out(far_7_7813_1[0]));    relay_conn far_7_7813_1_b(.in(far_7_7813_0[1]), .out(far_7_7813_1[1]));
    assign out[673] = ~far_7_7813_1[1]; 
    wire [1:0] far_7_7814_0;    relay_conn far_7_7814_0_a(.in(layer_6[1018]), .out(far_7_7814_0[0]));    relay_conn far_7_7814_0_b(.in(layer_6[971]), .out(far_7_7814_0[1]));
    assign out[674] = far_7_7814_0[0]; 
    wire [1:0] far_7_7815_0;    relay_conn far_7_7815_0_a(.in(layer_6[826]), .out(far_7_7815_0[0]));    relay_conn far_7_7815_0_b(.in(layer_6[931]), .out(far_7_7815_0[1]));
    wire [1:0] far_7_7815_1;    relay_conn far_7_7815_1_a(.in(far_7_7815_0[0]), .out(far_7_7815_1[0]));    relay_conn far_7_7815_1_b(.in(far_7_7815_0[1]), .out(far_7_7815_1[1]));
    wire [1:0] far_7_7815_2;    relay_conn far_7_7815_2_a(.in(far_7_7815_1[0]), .out(far_7_7815_2[0]));    relay_conn far_7_7815_2_b(.in(far_7_7815_1[1]), .out(far_7_7815_2[1]));
    assign out[675] = ~far_7_7815_2[1]; 
    assign out[676] = ~layer_6[388] | (layer_6[388] & layer_6[416]); 
    assign out[677] = layer_6[35] & layer_6[54]; 
    assign out[678] = ~layer_6[950]; 
    wire [1:0] far_7_7819_0;    relay_conn far_7_7819_0_a(.in(layer_6[178]), .out(far_7_7819_0[0]));    relay_conn far_7_7819_0_b(.in(layer_6[94]), .out(far_7_7819_0[1]));
    wire [1:0] far_7_7819_1;    relay_conn far_7_7819_1_a(.in(far_7_7819_0[0]), .out(far_7_7819_1[0]));    relay_conn far_7_7819_1_b(.in(far_7_7819_0[1]), .out(far_7_7819_1[1]));
    assign out[679] = far_7_7819_1[1]; 
    wire [1:0] far_7_7820_0;    relay_conn far_7_7820_0_a(.in(layer_6[737]), .out(far_7_7820_0[0]));    relay_conn far_7_7820_0_b(.in(layer_6[839]), .out(far_7_7820_0[1]));
    wire [1:0] far_7_7820_1;    relay_conn far_7_7820_1_a(.in(far_7_7820_0[0]), .out(far_7_7820_1[0]));    relay_conn far_7_7820_1_b(.in(far_7_7820_0[1]), .out(far_7_7820_1[1]));
    wire [1:0] far_7_7820_2;    relay_conn far_7_7820_2_a(.in(far_7_7820_1[0]), .out(far_7_7820_2[0]));    relay_conn far_7_7820_2_b(.in(far_7_7820_1[1]), .out(far_7_7820_2[1]));
    assign out[680] = ~far_7_7820_2[0]; 
    assign out[681] = layer_6[516] & ~layer_6[539]; 
    wire [1:0] far_7_7822_0;    relay_conn far_7_7822_0_a(.in(layer_6[76]), .out(far_7_7822_0[0]));    relay_conn far_7_7822_0_b(.in(layer_6[30]), .out(far_7_7822_0[1]));
    assign out[682] = far_7_7822_0[0] ^ far_7_7822_0[1]; 
    wire [1:0] far_7_7823_0;    relay_conn far_7_7823_0_a(.in(layer_6[499]), .out(far_7_7823_0[0]));    relay_conn far_7_7823_0_b(.in(layer_6[454]), .out(far_7_7823_0[1]));
    assign out[683] = ~far_7_7823_0[1]; 
    wire [1:0] far_7_7824_0;    relay_conn far_7_7824_0_a(.in(layer_6[573]), .out(far_7_7824_0[0]));    relay_conn far_7_7824_0_b(.in(layer_6[513]), .out(far_7_7824_0[1]));
    assign out[684] = ~far_7_7824_0[0]; 
    wire [1:0] far_7_7825_0;    relay_conn far_7_7825_0_a(.in(layer_6[953]), .out(far_7_7825_0[0]));    relay_conn far_7_7825_0_b(.in(layer_6[851]), .out(far_7_7825_0[1]));
    wire [1:0] far_7_7825_1;    relay_conn far_7_7825_1_a(.in(far_7_7825_0[0]), .out(far_7_7825_1[0]));    relay_conn far_7_7825_1_b(.in(far_7_7825_0[1]), .out(far_7_7825_1[1]));
    wire [1:0] far_7_7825_2;    relay_conn far_7_7825_2_a(.in(far_7_7825_1[0]), .out(far_7_7825_2[0]));    relay_conn far_7_7825_2_b(.in(far_7_7825_1[1]), .out(far_7_7825_2[1]));
    assign out[685] = far_7_7825_2[1] & ~far_7_7825_2[0]; 
    assign out[686] = layer_6[21] & layer_6[29]; 
    wire [1:0] far_7_7827_0;    relay_conn far_7_7827_0_a(.in(layer_6[552]), .out(far_7_7827_0[0]));    relay_conn far_7_7827_0_b(.in(layer_6[489]), .out(far_7_7827_0[1]));
    assign out[687] = far_7_7827_0[0] & far_7_7827_0[1]; 
    wire [1:0] far_7_7828_0;    relay_conn far_7_7828_0_a(.in(layer_6[267]), .out(far_7_7828_0[0]));    relay_conn far_7_7828_0_b(.in(layer_6[152]), .out(far_7_7828_0[1]));
    wire [1:0] far_7_7828_1;    relay_conn far_7_7828_1_a(.in(far_7_7828_0[0]), .out(far_7_7828_1[0]));    relay_conn far_7_7828_1_b(.in(far_7_7828_0[1]), .out(far_7_7828_1[1]));
    wire [1:0] far_7_7828_2;    relay_conn far_7_7828_2_a(.in(far_7_7828_1[0]), .out(far_7_7828_2[0]));    relay_conn far_7_7828_2_b(.in(far_7_7828_1[1]), .out(far_7_7828_2[1]));
    assign out[688] = ~far_7_7828_2[1]; 
    wire [1:0] far_7_7829_0;    relay_conn far_7_7829_0_a(.in(layer_6[487]), .out(far_7_7829_0[0]));    relay_conn far_7_7829_0_b(.in(layer_6[542]), .out(far_7_7829_0[1]));
    assign out[689] = ~far_7_7829_0[1]; 
    wire [1:0] far_7_7830_0;    relay_conn far_7_7830_0_a(.in(layer_6[778]), .out(far_7_7830_0[0]));    relay_conn far_7_7830_0_b(.in(layer_6[835]), .out(far_7_7830_0[1]));
    assign out[690] = far_7_7830_0[0]; 
    wire [1:0] far_7_7831_0;    relay_conn far_7_7831_0_a(.in(layer_6[43]), .out(far_7_7831_0[0]));    relay_conn far_7_7831_0_b(.in(layer_6[7]), .out(far_7_7831_0[1]));
    assign out[691] = ~far_7_7831_0[1]; 
    wire [1:0] far_7_7832_0;    relay_conn far_7_7832_0_a(.in(layer_6[507]), .out(far_7_7832_0[0]));    relay_conn far_7_7832_0_b(.in(layer_6[435]), .out(far_7_7832_0[1]));
    wire [1:0] far_7_7832_1;    relay_conn far_7_7832_1_a(.in(far_7_7832_0[0]), .out(far_7_7832_1[0]));    relay_conn far_7_7832_1_b(.in(far_7_7832_0[1]), .out(far_7_7832_1[1]));
    assign out[692] = ~far_7_7832_1[1]; 
    wire [1:0] far_7_7833_0;    relay_conn far_7_7833_0_a(.in(layer_6[507]), .out(far_7_7833_0[0]));    relay_conn far_7_7833_0_b(.in(layer_6[455]), .out(far_7_7833_0[1]));
    assign out[693] = far_7_7833_0[1]; 
    wire [1:0] far_7_7834_0;    relay_conn far_7_7834_0_a(.in(layer_6[762]), .out(far_7_7834_0[0]));    relay_conn far_7_7834_0_b(.in(layer_6[659]), .out(far_7_7834_0[1]));
    wire [1:0] far_7_7834_1;    relay_conn far_7_7834_1_a(.in(far_7_7834_0[0]), .out(far_7_7834_1[0]));    relay_conn far_7_7834_1_b(.in(far_7_7834_0[1]), .out(far_7_7834_1[1]));
    wire [1:0] far_7_7834_2;    relay_conn far_7_7834_2_a(.in(far_7_7834_1[0]), .out(far_7_7834_2[0]));    relay_conn far_7_7834_2_b(.in(far_7_7834_1[1]), .out(far_7_7834_2[1]));
    assign out[694] = far_7_7834_2[1] & ~far_7_7834_2[0]; 
    wire [1:0] far_7_7835_0;    relay_conn far_7_7835_0_a(.in(layer_6[599]), .out(far_7_7835_0[0]));    relay_conn far_7_7835_0_b(.in(layer_6[691]), .out(far_7_7835_0[1]));
    wire [1:0] far_7_7835_1;    relay_conn far_7_7835_1_a(.in(far_7_7835_0[0]), .out(far_7_7835_1[0]));    relay_conn far_7_7835_1_b(.in(far_7_7835_0[1]), .out(far_7_7835_1[1]));
    assign out[695] = far_7_7835_1[1] & ~far_7_7835_1[0]; 
    wire [1:0] far_7_7836_0;    relay_conn far_7_7836_0_a(.in(layer_6[364]), .out(far_7_7836_0[0]));    relay_conn far_7_7836_0_b(.in(layer_6[295]), .out(far_7_7836_0[1]));
    wire [1:0] far_7_7836_1;    relay_conn far_7_7836_1_a(.in(far_7_7836_0[0]), .out(far_7_7836_1[0]));    relay_conn far_7_7836_1_b(.in(far_7_7836_0[1]), .out(far_7_7836_1[1]));
    assign out[696] = far_7_7836_1[0] & far_7_7836_1[1]; 
    wire [1:0] far_7_7837_0;    relay_conn far_7_7837_0_a(.in(layer_6[171]), .out(far_7_7837_0[0]));    relay_conn far_7_7837_0_b(.in(layer_6[229]), .out(far_7_7837_0[1]));
    assign out[697] = ~(far_7_7837_0[0] ^ far_7_7837_0[1]); 
    wire [1:0] far_7_7838_0;    relay_conn far_7_7838_0_a(.in(layer_6[896]), .out(far_7_7838_0[0]));    relay_conn far_7_7838_0_b(.in(layer_6[814]), .out(far_7_7838_0[1]));
    wire [1:0] far_7_7838_1;    relay_conn far_7_7838_1_a(.in(far_7_7838_0[0]), .out(far_7_7838_1[0]));    relay_conn far_7_7838_1_b(.in(far_7_7838_0[1]), .out(far_7_7838_1[1]));
    assign out[698] = ~(far_7_7838_1[0] ^ far_7_7838_1[1]); 
    wire [1:0] far_7_7839_0;    relay_conn far_7_7839_0_a(.in(layer_6[766]), .out(far_7_7839_0[0]));    relay_conn far_7_7839_0_b(.in(layer_6[683]), .out(far_7_7839_0[1]));
    wire [1:0] far_7_7839_1;    relay_conn far_7_7839_1_a(.in(far_7_7839_0[0]), .out(far_7_7839_1[0]));    relay_conn far_7_7839_1_b(.in(far_7_7839_0[1]), .out(far_7_7839_1[1]));
    assign out[699] = far_7_7839_1[0] & far_7_7839_1[1]; 
    wire [1:0] far_7_7840_0;    relay_conn far_7_7840_0_a(.in(layer_6[395]), .out(far_7_7840_0[0]));    relay_conn far_7_7840_0_b(.in(layer_6[330]), .out(far_7_7840_0[1]));
    wire [1:0] far_7_7840_1;    relay_conn far_7_7840_1_a(.in(far_7_7840_0[0]), .out(far_7_7840_1[0]));    relay_conn far_7_7840_1_b(.in(far_7_7840_0[1]), .out(far_7_7840_1[1]));
    assign out[700] = far_7_7840_1[1] & ~far_7_7840_1[0]; 
    assign out[701] = layer_6[917]; 
    wire [1:0] far_7_7842_0;    relay_conn far_7_7842_0_a(.in(layer_6[730]), .out(far_7_7842_0[0]));    relay_conn far_7_7842_0_b(.in(layer_6[675]), .out(far_7_7842_0[1]));
    assign out[702] = far_7_7842_0[0] & ~far_7_7842_0[1]; 
    wire [1:0] far_7_7843_0;    relay_conn far_7_7843_0_a(.in(layer_6[260]), .out(far_7_7843_0[0]));    relay_conn far_7_7843_0_b(.in(layer_6[160]), .out(far_7_7843_0[1]));
    wire [1:0] far_7_7843_1;    relay_conn far_7_7843_1_a(.in(far_7_7843_0[0]), .out(far_7_7843_1[0]));    relay_conn far_7_7843_1_b(.in(far_7_7843_0[1]), .out(far_7_7843_1[1]));
    wire [1:0] far_7_7843_2;    relay_conn far_7_7843_2_a(.in(far_7_7843_1[0]), .out(far_7_7843_2[0]));    relay_conn far_7_7843_2_b(.in(far_7_7843_1[1]), .out(far_7_7843_2[1]));
    assign out[703] = ~far_7_7843_2[1]; 
    wire [1:0] far_7_7844_0;    relay_conn far_7_7844_0_a(.in(layer_6[913]), .out(far_7_7844_0[0]));    relay_conn far_7_7844_0_b(.in(layer_6[827]), .out(far_7_7844_0[1]));
    wire [1:0] far_7_7844_1;    relay_conn far_7_7844_1_a(.in(far_7_7844_0[0]), .out(far_7_7844_1[0]));    relay_conn far_7_7844_1_b(.in(far_7_7844_0[1]), .out(far_7_7844_1[1]));
    assign out[704] = ~far_7_7844_1[0] | (far_7_7844_1[0] & far_7_7844_1[1]); 
    wire [1:0] far_7_7845_0;    relay_conn far_7_7845_0_a(.in(layer_6[884]), .out(far_7_7845_0[0]));    relay_conn far_7_7845_0_b(.in(layer_6[935]), .out(far_7_7845_0[1]));
    assign out[705] = ~(far_7_7845_0[0] | far_7_7845_0[1]); 
    wire [1:0] far_7_7846_0;    relay_conn far_7_7846_0_a(.in(layer_6[741]), .out(far_7_7846_0[0]));    relay_conn far_7_7846_0_b(.in(layer_6[811]), .out(far_7_7846_0[1]));
    wire [1:0] far_7_7846_1;    relay_conn far_7_7846_1_a(.in(far_7_7846_0[0]), .out(far_7_7846_1[0]));    relay_conn far_7_7846_1_b(.in(far_7_7846_0[1]), .out(far_7_7846_1[1]));
    assign out[706] = far_7_7846_1[0] | far_7_7846_1[1]; 
    wire [1:0] far_7_7847_0;    relay_conn far_7_7847_0_a(.in(layer_6[315]), .out(far_7_7847_0[0]));    relay_conn far_7_7847_0_b(.in(layer_6[229]), .out(far_7_7847_0[1]));
    wire [1:0] far_7_7847_1;    relay_conn far_7_7847_1_a(.in(far_7_7847_0[0]), .out(far_7_7847_1[0]));    relay_conn far_7_7847_1_b(.in(far_7_7847_0[1]), .out(far_7_7847_1[1]));
    assign out[707] = ~far_7_7847_1[1]; 
    wire [1:0] far_7_7848_0;    relay_conn far_7_7848_0_a(.in(layer_6[777]), .out(far_7_7848_0[0]));    relay_conn far_7_7848_0_b(.in(layer_6[743]), .out(far_7_7848_0[1]));
    assign out[708] = ~far_7_7848_0[1]; 
    wire [1:0] far_7_7849_0;    relay_conn far_7_7849_0_a(.in(layer_6[456]), .out(far_7_7849_0[0]));    relay_conn far_7_7849_0_b(.in(layer_6[550]), .out(far_7_7849_0[1]));
    wire [1:0] far_7_7849_1;    relay_conn far_7_7849_1_a(.in(far_7_7849_0[0]), .out(far_7_7849_1[0]));    relay_conn far_7_7849_1_b(.in(far_7_7849_0[1]), .out(far_7_7849_1[1]));
    assign out[709] = ~(far_7_7849_1[0] ^ far_7_7849_1[1]); 
    wire [1:0] far_7_7850_0;    relay_conn far_7_7850_0_a(.in(layer_6[972]), .out(far_7_7850_0[0]));    relay_conn far_7_7850_0_b(.in(layer_6[896]), .out(far_7_7850_0[1]));
    wire [1:0] far_7_7850_1;    relay_conn far_7_7850_1_a(.in(far_7_7850_0[0]), .out(far_7_7850_1[0]));    relay_conn far_7_7850_1_b(.in(far_7_7850_0[1]), .out(far_7_7850_1[1]));
    assign out[710] = far_7_7850_1[0] ^ far_7_7850_1[1]; 
    assign out[711] = ~layer_6[422]; 
    assign out[712] = ~(layer_6[919] ^ layer_6[920]); 
    wire [1:0] far_7_7853_0;    relay_conn far_7_7853_0_a(.in(layer_6[358]), .out(far_7_7853_0[0]));    relay_conn far_7_7853_0_b(.in(layer_6[477]), .out(far_7_7853_0[1]));
    wire [1:0] far_7_7853_1;    relay_conn far_7_7853_1_a(.in(far_7_7853_0[0]), .out(far_7_7853_1[0]));    relay_conn far_7_7853_1_b(.in(far_7_7853_0[1]), .out(far_7_7853_1[1]));
    wire [1:0] far_7_7853_2;    relay_conn far_7_7853_2_a(.in(far_7_7853_1[0]), .out(far_7_7853_2[0]));    relay_conn far_7_7853_2_b(.in(far_7_7853_1[1]), .out(far_7_7853_2[1]));
    assign out[713] = far_7_7853_2[0] & ~far_7_7853_2[1]; 
    wire [1:0] far_7_7854_0;    relay_conn far_7_7854_0_a(.in(layer_6[737]), .out(far_7_7854_0[0]));    relay_conn far_7_7854_0_b(.in(layer_6[808]), .out(far_7_7854_0[1]));
    wire [1:0] far_7_7854_1;    relay_conn far_7_7854_1_a(.in(far_7_7854_0[0]), .out(far_7_7854_1[0]));    relay_conn far_7_7854_1_b(.in(far_7_7854_0[1]), .out(far_7_7854_1[1]));
    assign out[714] = far_7_7854_1[0] & far_7_7854_1[1]; 
    assign out[715] = ~layer_6[619]; 
    wire [1:0] far_7_7856_0;    relay_conn far_7_7856_0_a(.in(layer_6[453]), .out(far_7_7856_0[0]));    relay_conn far_7_7856_0_b(.in(layer_6[512]), .out(far_7_7856_0[1]));
    assign out[716] = ~(far_7_7856_0[0] | far_7_7856_0[1]); 
    wire [1:0] far_7_7857_0;    relay_conn far_7_7857_0_a(.in(layer_6[54]), .out(far_7_7857_0[0]));    relay_conn far_7_7857_0_b(.in(layer_6[110]), .out(far_7_7857_0[1]));
    assign out[717] = ~far_7_7857_0[1]; 
    wire [1:0] far_7_7858_0;    relay_conn far_7_7858_0_a(.in(layer_6[524]), .out(far_7_7858_0[0]));    relay_conn far_7_7858_0_b(.in(layer_6[404]), .out(far_7_7858_0[1]));
    wire [1:0] far_7_7858_1;    relay_conn far_7_7858_1_a(.in(far_7_7858_0[0]), .out(far_7_7858_1[0]));    relay_conn far_7_7858_1_b(.in(far_7_7858_0[1]), .out(far_7_7858_1[1]));
    wire [1:0] far_7_7858_2;    relay_conn far_7_7858_2_a(.in(far_7_7858_1[0]), .out(far_7_7858_2[0]));    relay_conn far_7_7858_2_b(.in(far_7_7858_1[1]), .out(far_7_7858_2[1]));
    assign out[718] = ~far_7_7858_2[0]; 
    wire [1:0] far_7_7859_0;    relay_conn far_7_7859_0_a(.in(layer_6[486]), .out(far_7_7859_0[0]));    relay_conn far_7_7859_0_b(.in(layer_6[610]), .out(far_7_7859_0[1]));
    wire [1:0] far_7_7859_1;    relay_conn far_7_7859_1_a(.in(far_7_7859_0[0]), .out(far_7_7859_1[0]));    relay_conn far_7_7859_1_b(.in(far_7_7859_0[1]), .out(far_7_7859_1[1]));
    wire [1:0] far_7_7859_2;    relay_conn far_7_7859_2_a(.in(far_7_7859_1[0]), .out(far_7_7859_2[0]));    relay_conn far_7_7859_2_b(.in(far_7_7859_1[1]), .out(far_7_7859_2[1]));
    assign out[719] = far_7_7859_2[0]; 
    wire [1:0] far_7_7860_0;    relay_conn far_7_7860_0_a(.in(layer_6[136]), .out(far_7_7860_0[0]));    relay_conn far_7_7860_0_b(.in(layer_6[230]), .out(far_7_7860_0[1]));
    wire [1:0] far_7_7860_1;    relay_conn far_7_7860_1_a(.in(far_7_7860_0[0]), .out(far_7_7860_1[0]));    relay_conn far_7_7860_1_b(.in(far_7_7860_0[1]), .out(far_7_7860_1[1]));
    assign out[720] = ~far_7_7860_1[1]; 
    wire [1:0] far_7_7861_0;    relay_conn far_7_7861_0_a(.in(layer_6[773]), .out(far_7_7861_0[0]));    relay_conn far_7_7861_0_b(.in(layer_6[685]), .out(far_7_7861_0[1]));
    wire [1:0] far_7_7861_1;    relay_conn far_7_7861_1_a(.in(far_7_7861_0[0]), .out(far_7_7861_1[0]));    relay_conn far_7_7861_1_b(.in(far_7_7861_0[1]), .out(far_7_7861_1[1]));
    assign out[721] = far_7_7861_1[0] ^ far_7_7861_1[1]; 
    wire [1:0] far_7_7862_0;    relay_conn far_7_7862_0_a(.in(layer_6[941]), .out(far_7_7862_0[0]));    relay_conn far_7_7862_0_b(.in(layer_6[825]), .out(far_7_7862_0[1]));
    wire [1:0] far_7_7862_1;    relay_conn far_7_7862_1_a(.in(far_7_7862_0[0]), .out(far_7_7862_1[0]));    relay_conn far_7_7862_1_b(.in(far_7_7862_0[1]), .out(far_7_7862_1[1]));
    wire [1:0] far_7_7862_2;    relay_conn far_7_7862_2_a(.in(far_7_7862_1[0]), .out(far_7_7862_2[0]));    relay_conn far_7_7862_2_b(.in(far_7_7862_1[1]), .out(far_7_7862_2[1]));
    assign out[722] = ~far_7_7862_2[1]; 
    assign out[723] = layer_6[30] & ~layer_6[2]; 
    wire [1:0] far_7_7864_0;    relay_conn far_7_7864_0_a(.in(layer_6[566]), .out(far_7_7864_0[0]));    relay_conn far_7_7864_0_b(.in(layer_6[632]), .out(far_7_7864_0[1]));
    wire [1:0] far_7_7864_1;    relay_conn far_7_7864_1_a(.in(far_7_7864_0[0]), .out(far_7_7864_1[0]));    relay_conn far_7_7864_1_b(.in(far_7_7864_0[1]), .out(far_7_7864_1[1]));
    assign out[724] = ~(far_7_7864_1[0] | far_7_7864_1[1]); 
    wire [1:0] far_7_7865_0;    relay_conn far_7_7865_0_a(.in(layer_6[504]), .out(far_7_7865_0[0]));    relay_conn far_7_7865_0_b(.in(layer_6[574]), .out(far_7_7865_0[1]));
    wire [1:0] far_7_7865_1;    relay_conn far_7_7865_1_a(.in(far_7_7865_0[0]), .out(far_7_7865_1[0]));    relay_conn far_7_7865_1_b(.in(far_7_7865_0[1]), .out(far_7_7865_1[1]));
    assign out[725] = far_7_7865_1[0]; 
    assign out[726] = ~(layer_6[142] & layer_6[140]); 
    wire [1:0] far_7_7867_0;    relay_conn far_7_7867_0_a(.in(layer_6[857]), .out(far_7_7867_0[0]));    relay_conn far_7_7867_0_b(.in(layer_6[967]), .out(far_7_7867_0[1]));
    wire [1:0] far_7_7867_1;    relay_conn far_7_7867_1_a(.in(far_7_7867_0[0]), .out(far_7_7867_1[0]));    relay_conn far_7_7867_1_b(.in(far_7_7867_0[1]), .out(far_7_7867_1[1]));
    wire [1:0] far_7_7867_2;    relay_conn far_7_7867_2_a(.in(far_7_7867_1[0]), .out(far_7_7867_2[0]));    relay_conn far_7_7867_2_b(.in(far_7_7867_1[1]), .out(far_7_7867_2[1]));
    assign out[727] = ~far_7_7867_2[1]; 
    assign out[728] = ~(layer_6[928] & layer_6[923]); 
    assign out[729] = layer_6[465]; 
    assign out[730] = layer_6[98] & ~layer_6[128]; 
    wire [1:0] far_7_7871_0;    relay_conn far_7_7871_0_a(.in(layer_6[397]), .out(far_7_7871_0[0]));    relay_conn far_7_7871_0_b(.in(layer_6[525]), .out(far_7_7871_0[1]));
    wire [1:0] far_7_7871_1;    relay_conn far_7_7871_1_a(.in(far_7_7871_0[0]), .out(far_7_7871_1[0]));    relay_conn far_7_7871_1_b(.in(far_7_7871_0[1]), .out(far_7_7871_1[1]));
    wire [1:0] far_7_7871_2;    relay_conn far_7_7871_2_a(.in(far_7_7871_1[0]), .out(far_7_7871_2[0]));    relay_conn far_7_7871_2_b(.in(far_7_7871_1[1]), .out(far_7_7871_2[1]));
    wire [1:0] far_7_7871_3;    relay_conn far_7_7871_3_a(.in(far_7_7871_2[0]), .out(far_7_7871_3[0]));    relay_conn far_7_7871_3_b(.in(far_7_7871_2[1]), .out(far_7_7871_3[1]));
    assign out[731] = far_7_7871_3[1]; 
    assign out[732] = ~layer_6[100]; 
    assign out[733] = layer_6[337]; 
    wire [1:0] far_7_7874_0;    relay_conn far_7_7874_0_a(.in(layer_6[9]), .out(far_7_7874_0[0]));    relay_conn far_7_7874_0_b(.in(layer_6[71]), .out(far_7_7874_0[1]));
    assign out[734] = far_7_7874_0[1] & ~far_7_7874_0[0]; 
    wire [1:0] far_7_7875_0;    relay_conn far_7_7875_0_a(.in(layer_6[605]), .out(far_7_7875_0[0]));    relay_conn far_7_7875_0_b(.in(layer_6[652]), .out(far_7_7875_0[1]));
    assign out[735] = far_7_7875_0[0] | far_7_7875_0[1]; 
    wire [1:0] far_7_7876_0;    relay_conn far_7_7876_0_a(.in(layer_6[422]), .out(far_7_7876_0[0]));    relay_conn far_7_7876_0_b(.in(layer_6[512]), .out(far_7_7876_0[1]));
    wire [1:0] far_7_7876_1;    relay_conn far_7_7876_1_a(.in(far_7_7876_0[0]), .out(far_7_7876_1[0]));    relay_conn far_7_7876_1_b(.in(far_7_7876_0[1]), .out(far_7_7876_1[1]));
    assign out[736] = far_7_7876_1[0] & ~far_7_7876_1[1]; 
    assign out[737] = layer_6[68]; 
    assign out[738] = layer_6[913]; 
    wire [1:0] far_7_7879_0;    relay_conn far_7_7879_0_a(.in(layer_6[1019]), .out(far_7_7879_0[0]));    relay_conn far_7_7879_0_b(.in(layer_6[931]), .out(far_7_7879_0[1]));
    wire [1:0] far_7_7879_1;    relay_conn far_7_7879_1_a(.in(far_7_7879_0[0]), .out(far_7_7879_1[0]));    relay_conn far_7_7879_1_b(.in(far_7_7879_0[1]), .out(far_7_7879_1[1]));
    assign out[739] = far_7_7879_1[0] & far_7_7879_1[1]; 
    assign out[740] = layer_6[643] | layer_6[629]; 
    wire [1:0] far_7_7881_0;    relay_conn far_7_7881_0_a(.in(layer_6[730]), .out(far_7_7881_0[0]));    relay_conn far_7_7881_0_b(.in(layer_6[816]), .out(far_7_7881_0[1]));
    wire [1:0] far_7_7881_1;    relay_conn far_7_7881_1_a(.in(far_7_7881_0[0]), .out(far_7_7881_1[0]));    relay_conn far_7_7881_1_b(.in(far_7_7881_0[1]), .out(far_7_7881_1[1]));
    assign out[741] = ~(far_7_7881_1[0] | far_7_7881_1[1]); 
    assign out[742] = ~layer_6[825]; 
    assign out[743] = ~layer_6[642]; 
    wire [1:0] far_7_7884_0;    relay_conn far_7_7884_0_a(.in(layer_6[392]), .out(far_7_7884_0[0]));    relay_conn far_7_7884_0_b(.in(layer_6[320]), .out(far_7_7884_0[1]));
    wire [1:0] far_7_7884_1;    relay_conn far_7_7884_1_a(.in(far_7_7884_0[0]), .out(far_7_7884_1[0]));    relay_conn far_7_7884_1_b(.in(far_7_7884_0[1]), .out(far_7_7884_1[1]));
    assign out[744] = far_7_7884_1[1]; 
    assign out[745] = ~(layer_6[296] ^ layer_6[270]); 
    wire [1:0] far_7_7886_0;    relay_conn far_7_7886_0_a(.in(layer_6[623]), .out(far_7_7886_0[0]));    relay_conn far_7_7886_0_b(.in(layer_6[681]), .out(far_7_7886_0[1]));
    assign out[746] = ~(far_7_7886_0[0] ^ far_7_7886_0[1]); 
    wire [1:0] far_7_7887_0;    relay_conn far_7_7887_0_a(.in(layer_6[132]), .out(far_7_7887_0[0]));    relay_conn far_7_7887_0_b(.in(layer_6[56]), .out(far_7_7887_0[1]));
    wire [1:0] far_7_7887_1;    relay_conn far_7_7887_1_a(.in(far_7_7887_0[0]), .out(far_7_7887_1[0]));    relay_conn far_7_7887_1_b(.in(far_7_7887_0[1]), .out(far_7_7887_1[1]));
    assign out[747] = far_7_7887_1[1] & ~far_7_7887_1[0]; 
    wire [1:0] far_7_7888_0;    relay_conn far_7_7888_0_a(.in(layer_6[453]), .out(far_7_7888_0[0]));    relay_conn far_7_7888_0_b(.in(layer_6[343]), .out(far_7_7888_0[1]));
    wire [1:0] far_7_7888_1;    relay_conn far_7_7888_1_a(.in(far_7_7888_0[0]), .out(far_7_7888_1[0]));    relay_conn far_7_7888_1_b(.in(far_7_7888_0[1]), .out(far_7_7888_1[1]));
    wire [1:0] far_7_7888_2;    relay_conn far_7_7888_2_a(.in(far_7_7888_1[0]), .out(far_7_7888_2[0]));    relay_conn far_7_7888_2_b(.in(far_7_7888_1[1]), .out(far_7_7888_2[1]));
    assign out[748] = ~(far_7_7888_2[0] | far_7_7888_2[1]); 
    assign out[749] = layer_6[612] & ~layer_6[603]; 
    wire [1:0] far_7_7890_0;    relay_conn far_7_7890_0_a(.in(layer_6[130]), .out(far_7_7890_0[0]));    relay_conn far_7_7890_0_b(.in(layer_6[80]), .out(far_7_7890_0[1]));
    assign out[750] = ~far_7_7890_0[0]; 
    wire [1:0] far_7_7891_0;    relay_conn far_7_7891_0_a(.in(layer_6[257]), .out(far_7_7891_0[0]));    relay_conn far_7_7891_0_b(.in(layer_6[192]), .out(far_7_7891_0[1]));
    wire [1:0] far_7_7891_1;    relay_conn far_7_7891_1_a(.in(far_7_7891_0[0]), .out(far_7_7891_1[0]));    relay_conn far_7_7891_1_b(.in(far_7_7891_0[1]), .out(far_7_7891_1[1]));
    assign out[751] = far_7_7891_1[0] & ~far_7_7891_1[1]; 
    wire [1:0] far_7_7892_0;    relay_conn far_7_7892_0_a(.in(layer_6[200]), .out(far_7_7892_0[0]));    relay_conn far_7_7892_0_b(.in(layer_6[315]), .out(far_7_7892_0[1]));
    wire [1:0] far_7_7892_1;    relay_conn far_7_7892_1_a(.in(far_7_7892_0[0]), .out(far_7_7892_1[0]));    relay_conn far_7_7892_1_b(.in(far_7_7892_0[1]), .out(far_7_7892_1[1]));
    wire [1:0] far_7_7892_2;    relay_conn far_7_7892_2_a(.in(far_7_7892_1[0]), .out(far_7_7892_2[0]));    relay_conn far_7_7892_2_b(.in(far_7_7892_1[1]), .out(far_7_7892_2[1]));
    assign out[752] = ~(far_7_7892_2[0] ^ far_7_7892_2[1]); 
    assign out[753] = ~layer_6[181]; 
    wire [1:0] far_7_7894_0;    relay_conn far_7_7894_0_a(.in(layer_6[896]), .out(far_7_7894_0[0]));    relay_conn far_7_7894_0_b(.in(layer_6[799]), .out(far_7_7894_0[1]));
    wire [1:0] far_7_7894_1;    relay_conn far_7_7894_1_a(.in(far_7_7894_0[0]), .out(far_7_7894_1[0]));    relay_conn far_7_7894_1_b(.in(far_7_7894_0[1]), .out(far_7_7894_1[1]));
    wire [1:0] far_7_7894_2;    relay_conn far_7_7894_2_a(.in(far_7_7894_1[0]), .out(far_7_7894_2[0]));    relay_conn far_7_7894_2_b(.in(far_7_7894_1[1]), .out(far_7_7894_2[1]));
    assign out[754] = far_7_7894_2[1] & ~far_7_7894_2[0]; 
    wire [1:0] far_7_7895_0;    relay_conn far_7_7895_0_a(.in(layer_6[766]), .out(far_7_7895_0[0]));    relay_conn far_7_7895_0_b(.in(layer_6[821]), .out(far_7_7895_0[1]));
    assign out[755] = far_7_7895_0[1]; 
    wire [1:0] far_7_7896_0;    relay_conn far_7_7896_0_a(.in(layer_6[971]), .out(far_7_7896_0[0]));    relay_conn far_7_7896_0_b(.in(layer_6[935]), .out(far_7_7896_0[1]));
    assign out[756] = ~(far_7_7896_0[0] ^ far_7_7896_0[1]); 
    wire [1:0] far_7_7897_0;    relay_conn far_7_7897_0_a(.in(layer_6[390]), .out(far_7_7897_0[0]));    relay_conn far_7_7897_0_b(.in(layer_6[278]), .out(far_7_7897_0[1]));
    wire [1:0] far_7_7897_1;    relay_conn far_7_7897_1_a(.in(far_7_7897_0[0]), .out(far_7_7897_1[0]));    relay_conn far_7_7897_1_b(.in(far_7_7897_0[1]), .out(far_7_7897_1[1]));
    wire [1:0] far_7_7897_2;    relay_conn far_7_7897_2_a(.in(far_7_7897_1[0]), .out(far_7_7897_2[0]));    relay_conn far_7_7897_2_b(.in(far_7_7897_1[1]), .out(far_7_7897_2[1]));
    assign out[757] = ~(far_7_7897_2[0] ^ far_7_7897_2[1]); 
    assign out[758] = ~layer_6[691]; 
    wire [1:0] far_7_7899_0;    relay_conn far_7_7899_0_a(.in(layer_6[1016]), .out(far_7_7899_0[0]));    relay_conn far_7_7899_0_b(.in(layer_6[904]), .out(far_7_7899_0[1]));
    wire [1:0] far_7_7899_1;    relay_conn far_7_7899_1_a(.in(far_7_7899_0[0]), .out(far_7_7899_1[0]));    relay_conn far_7_7899_1_b(.in(far_7_7899_0[1]), .out(far_7_7899_1[1]));
    wire [1:0] far_7_7899_2;    relay_conn far_7_7899_2_a(.in(far_7_7899_1[0]), .out(far_7_7899_2[0]));    relay_conn far_7_7899_2_b(.in(far_7_7899_1[1]), .out(far_7_7899_2[1]));
    assign out[759] = far_7_7899_2[0] & ~far_7_7899_2[1]; 
    wire [1:0] far_7_7900_0;    relay_conn far_7_7900_0_a(.in(layer_6[538]), .out(far_7_7900_0[0]));    relay_conn far_7_7900_0_b(.in(layer_6[623]), .out(far_7_7900_0[1]));
    wire [1:0] far_7_7900_1;    relay_conn far_7_7900_1_a(.in(far_7_7900_0[0]), .out(far_7_7900_1[0]));    relay_conn far_7_7900_1_b(.in(far_7_7900_0[1]), .out(far_7_7900_1[1]));
    assign out[760] = far_7_7900_1[0] ^ far_7_7900_1[1]; 
    wire [1:0] far_7_7901_0;    relay_conn far_7_7901_0_a(.in(layer_6[413]), .out(far_7_7901_0[0]));    relay_conn far_7_7901_0_b(.in(layer_6[460]), .out(far_7_7901_0[1]));
    assign out[761] = ~far_7_7901_0[1]; 
    wire [1:0] far_7_7902_0;    relay_conn far_7_7902_0_a(.in(layer_6[493]), .out(far_7_7902_0[0]));    relay_conn far_7_7902_0_b(.in(layer_6[404]), .out(far_7_7902_0[1]));
    wire [1:0] far_7_7902_1;    relay_conn far_7_7902_1_a(.in(far_7_7902_0[0]), .out(far_7_7902_1[0]));    relay_conn far_7_7902_1_b(.in(far_7_7902_0[1]), .out(far_7_7902_1[1]));
    assign out[762] = ~(far_7_7902_1[0] ^ far_7_7902_1[1]); 
    wire [1:0] far_7_7903_0;    relay_conn far_7_7903_0_a(.in(layer_6[483]), .out(far_7_7903_0[0]));    relay_conn far_7_7903_0_b(.in(layer_6[424]), .out(far_7_7903_0[1]));
    assign out[763] = ~far_7_7903_0[0]; 
    wire [1:0] far_7_7904_0;    relay_conn far_7_7904_0_a(.in(layer_6[61]), .out(far_7_7904_0[0]));    relay_conn far_7_7904_0_b(.in(layer_6[148]), .out(far_7_7904_0[1]));
    wire [1:0] far_7_7904_1;    relay_conn far_7_7904_1_a(.in(far_7_7904_0[0]), .out(far_7_7904_1[0]));    relay_conn far_7_7904_1_b(.in(far_7_7904_0[1]), .out(far_7_7904_1[1]));
    assign out[764] = ~far_7_7904_1[1]; 
    wire [1:0] far_7_7905_0;    relay_conn far_7_7905_0_a(.in(layer_6[995]), .out(far_7_7905_0[0]));    relay_conn far_7_7905_0_b(.in(layer_6[959]), .out(far_7_7905_0[1]));
    assign out[765] = far_7_7905_0[0]; 
    assign out[766] = ~(layer_6[254] & layer_6[255]); 
    wire [1:0] far_7_7907_0;    relay_conn far_7_7907_0_a(.in(layer_6[404]), .out(far_7_7907_0[0]));    relay_conn far_7_7907_0_b(.in(layer_6[439]), .out(far_7_7907_0[1]));
    assign out[767] = far_7_7907_0[0]; 
    wire [1:0] far_7_7908_0;    relay_conn far_7_7908_0_a(.in(layer_6[574]), .out(far_7_7908_0[0]));    relay_conn far_7_7908_0_b(.in(layer_6[531]), .out(far_7_7908_0[1]));
    assign out[768] = ~(far_7_7908_0[0] | far_7_7908_0[1]); 
    assign out[769] = ~layer_6[923] | (layer_6[925] & layer_6[923]); 
    assign out[770] = layer_6[995] & layer_6[972]; 
    wire [1:0] far_7_7911_0;    relay_conn far_7_7911_0_a(.in(layer_6[215]), .out(far_7_7911_0[0]));    relay_conn far_7_7911_0_b(.in(layer_6[324]), .out(far_7_7911_0[1]));
    wire [1:0] far_7_7911_1;    relay_conn far_7_7911_1_a(.in(far_7_7911_0[0]), .out(far_7_7911_1[0]));    relay_conn far_7_7911_1_b(.in(far_7_7911_0[1]), .out(far_7_7911_1[1]));
    wire [1:0] far_7_7911_2;    relay_conn far_7_7911_2_a(.in(far_7_7911_1[0]), .out(far_7_7911_2[0]));    relay_conn far_7_7911_2_b(.in(far_7_7911_1[1]), .out(far_7_7911_2[1]));
    assign out[771] = ~(far_7_7911_2[0] | far_7_7911_2[1]); 
    wire [1:0] far_7_7912_0;    relay_conn far_7_7912_0_a(.in(layer_6[191]), .out(far_7_7912_0[0]));    relay_conn far_7_7912_0_b(.in(layer_6[285]), .out(far_7_7912_0[1]));
    wire [1:0] far_7_7912_1;    relay_conn far_7_7912_1_a(.in(far_7_7912_0[0]), .out(far_7_7912_1[0]));    relay_conn far_7_7912_1_b(.in(far_7_7912_0[1]), .out(far_7_7912_1[1]));
    assign out[772] = far_7_7912_1[1]; 
    assign out[773] = layer_6[126]; 
    wire [1:0] far_7_7914_0;    relay_conn far_7_7914_0_a(.in(layer_6[60]), .out(far_7_7914_0[0]));    relay_conn far_7_7914_0_b(.in(layer_6[144]), .out(far_7_7914_0[1]));
    wire [1:0] far_7_7914_1;    relay_conn far_7_7914_1_a(.in(far_7_7914_0[0]), .out(far_7_7914_1[0]));    relay_conn far_7_7914_1_b(.in(far_7_7914_0[1]), .out(far_7_7914_1[1]));
    assign out[774] = far_7_7914_1[0] & ~far_7_7914_1[1]; 
    wire [1:0] far_7_7915_0;    relay_conn far_7_7915_0_a(.in(layer_6[757]), .out(far_7_7915_0[0]));    relay_conn far_7_7915_0_b(.in(layer_6[837]), .out(far_7_7915_0[1]));
    wire [1:0] far_7_7915_1;    relay_conn far_7_7915_1_a(.in(far_7_7915_0[0]), .out(far_7_7915_1[0]));    relay_conn far_7_7915_1_b(.in(far_7_7915_0[1]), .out(far_7_7915_1[1]));
    assign out[775] = far_7_7915_1[1]; 
    wire [1:0] far_7_7916_0;    relay_conn far_7_7916_0_a(.in(layer_6[157]), .out(far_7_7916_0[0]));    relay_conn far_7_7916_0_b(.in(layer_6[247]), .out(far_7_7916_0[1]));
    wire [1:0] far_7_7916_1;    relay_conn far_7_7916_1_a(.in(far_7_7916_0[0]), .out(far_7_7916_1[0]));    relay_conn far_7_7916_1_b(.in(far_7_7916_0[1]), .out(far_7_7916_1[1]));
    assign out[776] = ~far_7_7916_1[0]; 
    wire [1:0] far_7_7917_0;    relay_conn far_7_7917_0_a(.in(layer_6[331]), .out(far_7_7917_0[0]));    relay_conn far_7_7917_0_b(.in(layer_6[388]), .out(far_7_7917_0[1]));
    assign out[777] = ~far_7_7917_0[0]; 
    wire [1:0] far_7_7918_0;    relay_conn far_7_7918_0_a(.in(layer_6[542]), .out(far_7_7918_0[0]));    relay_conn far_7_7918_0_b(.in(layer_6[475]), .out(far_7_7918_0[1]));
    wire [1:0] far_7_7918_1;    relay_conn far_7_7918_1_a(.in(far_7_7918_0[0]), .out(far_7_7918_1[0]));    relay_conn far_7_7918_1_b(.in(far_7_7918_0[1]), .out(far_7_7918_1[1]));
    assign out[778] = far_7_7918_1[0] & ~far_7_7918_1[1]; 
    wire [1:0] far_7_7919_0;    relay_conn far_7_7919_0_a(.in(layer_6[991]), .out(far_7_7919_0[0]));    relay_conn far_7_7919_0_b(.in(layer_6[950]), .out(far_7_7919_0[1]));
    assign out[779] = far_7_7919_0[1] & ~far_7_7919_0[0]; 
    wire [1:0] far_7_7920_0;    relay_conn far_7_7920_0_a(.in(layer_6[763]), .out(far_7_7920_0[0]));    relay_conn far_7_7920_0_b(.in(layer_6[638]), .out(far_7_7920_0[1]));
    wire [1:0] far_7_7920_1;    relay_conn far_7_7920_1_a(.in(far_7_7920_0[0]), .out(far_7_7920_1[0]));    relay_conn far_7_7920_1_b(.in(far_7_7920_0[1]), .out(far_7_7920_1[1]));
    wire [1:0] far_7_7920_2;    relay_conn far_7_7920_2_a(.in(far_7_7920_1[0]), .out(far_7_7920_2[0]));    relay_conn far_7_7920_2_b(.in(far_7_7920_1[1]), .out(far_7_7920_2[1]));
    assign out[780] = far_7_7920_2[0] & far_7_7920_2[1]; 
    assign out[781] = layer_6[720] & ~layer_6[732]; 
    wire [1:0] far_7_7922_0;    relay_conn far_7_7922_0_a(.in(layer_6[499]), .out(far_7_7922_0[0]));    relay_conn far_7_7922_0_b(.in(layer_6[614]), .out(far_7_7922_0[1]));
    wire [1:0] far_7_7922_1;    relay_conn far_7_7922_1_a(.in(far_7_7922_0[0]), .out(far_7_7922_1[0]));    relay_conn far_7_7922_1_b(.in(far_7_7922_0[1]), .out(far_7_7922_1[1]));
    wire [1:0] far_7_7922_2;    relay_conn far_7_7922_2_a(.in(far_7_7922_1[0]), .out(far_7_7922_2[0]));    relay_conn far_7_7922_2_b(.in(far_7_7922_1[1]), .out(far_7_7922_2[1]));
    assign out[782] = ~(far_7_7922_2[0] | far_7_7922_2[1]); 
    wire [1:0] far_7_7923_0;    relay_conn far_7_7923_0_a(.in(layer_6[312]), .out(far_7_7923_0[0]));    relay_conn far_7_7923_0_b(.in(layer_6[360]), .out(far_7_7923_0[1]));
    assign out[783] = ~(far_7_7923_0[0] | far_7_7923_0[1]); 
    assign out[784] = ~(layer_6[40] ^ layer_6[51]); 
    wire [1:0] far_7_7925_0;    relay_conn far_7_7925_0_a(.in(layer_6[994]), .out(far_7_7925_0[0]));    relay_conn far_7_7925_0_b(.in(layer_6[891]), .out(far_7_7925_0[1]));
    wire [1:0] far_7_7925_1;    relay_conn far_7_7925_1_a(.in(far_7_7925_0[0]), .out(far_7_7925_1[0]));    relay_conn far_7_7925_1_b(.in(far_7_7925_0[1]), .out(far_7_7925_1[1]));
    wire [1:0] far_7_7925_2;    relay_conn far_7_7925_2_a(.in(far_7_7925_1[0]), .out(far_7_7925_2[0]));    relay_conn far_7_7925_2_b(.in(far_7_7925_1[1]), .out(far_7_7925_2[1]));
    assign out[785] = ~(far_7_7925_2[0] | far_7_7925_2[1]); 
    wire [1:0] far_7_7926_0;    relay_conn far_7_7926_0_a(.in(layer_6[720]), .out(far_7_7926_0[0]));    relay_conn far_7_7926_0_b(.in(layer_6[845]), .out(far_7_7926_0[1]));
    wire [1:0] far_7_7926_1;    relay_conn far_7_7926_1_a(.in(far_7_7926_0[0]), .out(far_7_7926_1[0]));    relay_conn far_7_7926_1_b(.in(far_7_7926_0[1]), .out(far_7_7926_1[1]));
    wire [1:0] far_7_7926_2;    relay_conn far_7_7926_2_a(.in(far_7_7926_1[0]), .out(far_7_7926_2[0]));    relay_conn far_7_7926_2_b(.in(far_7_7926_1[1]), .out(far_7_7926_2[1]));
    assign out[786] = far_7_7926_2[0] & far_7_7926_2[1]; 
    wire [1:0] far_7_7927_0;    relay_conn far_7_7927_0_a(.in(layer_6[741]), .out(far_7_7927_0[0]));    relay_conn far_7_7927_0_b(.in(layer_6[821]), .out(far_7_7927_0[1]));
    wire [1:0] far_7_7927_1;    relay_conn far_7_7927_1_a(.in(far_7_7927_0[0]), .out(far_7_7927_1[0]));    relay_conn far_7_7927_1_b(.in(far_7_7927_0[1]), .out(far_7_7927_1[1]));
    assign out[787] = far_7_7927_1[1]; 
    wire [1:0] far_7_7928_0;    relay_conn far_7_7928_0_a(.in(layer_6[624]), .out(far_7_7928_0[0]));    relay_conn far_7_7928_0_b(.in(layer_6[511]), .out(far_7_7928_0[1]));
    wire [1:0] far_7_7928_1;    relay_conn far_7_7928_1_a(.in(far_7_7928_0[0]), .out(far_7_7928_1[0]));    relay_conn far_7_7928_1_b(.in(far_7_7928_0[1]), .out(far_7_7928_1[1]));
    wire [1:0] far_7_7928_2;    relay_conn far_7_7928_2_a(.in(far_7_7928_1[0]), .out(far_7_7928_2[0]));    relay_conn far_7_7928_2_b(.in(far_7_7928_1[1]), .out(far_7_7928_2[1]));
    assign out[788] = ~far_7_7928_2[1]; 
    wire [1:0] far_7_7929_0;    relay_conn far_7_7929_0_a(.in(layer_6[677]), .out(far_7_7929_0[0]));    relay_conn far_7_7929_0_b(.in(layer_6[605]), .out(far_7_7929_0[1]));
    wire [1:0] far_7_7929_1;    relay_conn far_7_7929_1_a(.in(far_7_7929_0[0]), .out(far_7_7929_1[0]));    relay_conn far_7_7929_1_b(.in(far_7_7929_0[1]), .out(far_7_7929_1[1]));
    assign out[789] = far_7_7929_1[0] & far_7_7929_1[1]; 
    assign out[790] = layer_6[169] & ~layer_6[167]; 
    wire [1:0] far_7_7931_0;    relay_conn far_7_7931_0_a(.in(layer_6[428]), .out(far_7_7931_0[0]));    relay_conn far_7_7931_0_b(.in(layer_6[329]), .out(far_7_7931_0[1]));
    wire [1:0] far_7_7931_1;    relay_conn far_7_7931_1_a(.in(far_7_7931_0[0]), .out(far_7_7931_1[0]));    relay_conn far_7_7931_1_b(.in(far_7_7931_0[1]), .out(far_7_7931_1[1]));
    wire [1:0] far_7_7931_2;    relay_conn far_7_7931_2_a(.in(far_7_7931_1[0]), .out(far_7_7931_2[0]));    relay_conn far_7_7931_2_b(.in(far_7_7931_1[1]), .out(far_7_7931_2[1]));
    assign out[791] = far_7_7931_2[0]; 
    wire [1:0] far_7_7932_0;    relay_conn far_7_7932_0_a(.in(layer_6[995]), .out(far_7_7932_0[0]));    relay_conn far_7_7932_0_b(.in(layer_6[920]), .out(far_7_7932_0[1]));
    wire [1:0] far_7_7932_1;    relay_conn far_7_7932_1_a(.in(far_7_7932_0[0]), .out(far_7_7932_1[0]));    relay_conn far_7_7932_1_b(.in(far_7_7932_0[1]), .out(far_7_7932_1[1]));
    assign out[792] = far_7_7932_1[0]; 
    wire [1:0] far_7_7933_0;    relay_conn far_7_7933_0_a(.in(layer_6[706]), .out(far_7_7933_0[0]));    relay_conn far_7_7933_0_b(.in(layer_6[648]), .out(far_7_7933_0[1]));
    assign out[793] = far_7_7933_0[0] ^ far_7_7933_0[1]; 
    wire [1:0] far_7_7934_0;    relay_conn far_7_7934_0_a(.in(layer_6[94]), .out(far_7_7934_0[0]));    relay_conn far_7_7934_0_b(.in(layer_6[220]), .out(far_7_7934_0[1]));
    wire [1:0] far_7_7934_1;    relay_conn far_7_7934_1_a(.in(far_7_7934_0[0]), .out(far_7_7934_1[0]));    relay_conn far_7_7934_1_b(.in(far_7_7934_0[1]), .out(far_7_7934_1[1]));
    wire [1:0] far_7_7934_2;    relay_conn far_7_7934_2_a(.in(far_7_7934_1[0]), .out(far_7_7934_2[0]));    relay_conn far_7_7934_2_b(.in(far_7_7934_1[1]), .out(far_7_7934_2[1]));
    assign out[794] = far_7_7934_2[1] & ~far_7_7934_2[0]; 
    wire [1:0] far_7_7935_0;    relay_conn far_7_7935_0_a(.in(layer_6[955]), .out(far_7_7935_0[0]));    relay_conn far_7_7935_0_b(.in(layer_6[999]), .out(far_7_7935_0[1]));
    assign out[795] = far_7_7935_0[1]; 
    wire [1:0] far_7_7936_0;    relay_conn far_7_7936_0_a(.in(layer_6[210]), .out(far_7_7936_0[0]));    relay_conn far_7_7936_0_b(.in(layer_6[270]), .out(far_7_7936_0[1]));
    assign out[796] = ~(far_7_7936_0[0] | far_7_7936_0[1]); 
    wire [1:0] far_7_7937_0;    relay_conn far_7_7937_0_a(.in(layer_6[540]), .out(far_7_7937_0[0]));    relay_conn far_7_7937_0_b(.in(layer_6[643]), .out(far_7_7937_0[1]));
    wire [1:0] far_7_7937_1;    relay_conn far_7_7937_1_a(.in(far_7_7937_0[0]), .out(far_7_7937_1[0]));    relay_conn far_7_7937_1_b(.in(far_7_7937_0[1]), .out(far_7_7937_1[1]));
    wire [1:0] far_7_7937_2;    relay_conn far_7_7937_2_a(.in(far_7_7937_1[0]), .out(far_7_7937_2[0]));    relay_conn far_7_7937_2_b(.in(far_7_7937_1[1]), .out(far_7_7937_2[1]));
    assign out[797] = ~far_7_7937_2[0]; 
    wire [1:0] far_7_7938_0;    relay_conn far_7_7938_0_a(.in(layer_6[14]), .out(far_7_7938_0[0]));    relay_conn far_7_7938_0_b(.in(layer_6[116]), .out(far_7_7938_0[1]));
    wire [1:0] far_7_7938_1;    relay_conn far_7_7938_1_a(.in(far_7_7938_0[0]), .out(far_7_7938_1[0]));    relay_conn far_7_7938_1_b(.in(far_7_7938_0[1]), .out(far_7_7938_1[1]));
    wire [1:0] far_7_7938_2;    relay_conn far_7_7938_2_a(.in(far_7_7938_1[0]), .out(far_7_7938_2[0]));    relay_conn far_7_7938_2_b(.in(far_7_7938_1[1]), .out(far_7_7938_2[1]));
    assign out[798] = ~(far_7_7938_2[0] | far_7_7938_2[1]); 
    wire [1:0] far_7_7939_0;    relay_conn far_7_7939_0_a(.in(layer_6[260]), .out(far_7_7939_0[0]));    relay_conn far_7_7939_0_b(.in(layer_6[155]), .out(far_7_7939_0[1]));
    wire [1:0] far_7_7939_1;    relay_conn far_7_7939_1_a(.in(far_7_7939_0[0]), .out(far_7_7939_1[0]));    relay_conn far_7_7939_1_b(.in(far_7_7939_0[1]), .out(far_7_7939_1[1]));
    wire [1:0] far_7_7939_2;    relay_conn far_7_7939_2_a(.in(far_7_7939_1[0]), .out(far_7_7939_2[0]));    relay_conn far_7_7939_2_b(.in(far_7_7939_1[1]), .out(far_7_7939_2[1]));
    assign out[799] = far_7_7939_2[1]; 
    wire [1:0] far_7_7940_0;    relay_conn far_7_7940_0_a(.in(layer_6[766]), .out(far_7_7940_0[0]));    relay_conn far_7_7940_0_b(.in(layer_6[730]), .out(far_7_7940_0[1]));
    assign out[800] = ~(far_7_7940_0[0] & far_7_7940_0[1]); 
    wire [1:0] far_7_7941_0;    relay_conn far_7_7941_0_a(.in(layer_6[874]), .out(far_7_7941_0[0]));    relay_conn far_7_7941_0_b(.in(layer_6[758]), .out(far_7_7941_0[1]));
    wire [1:0] far_7_7941_1;    relay_conn far_7_7941_1_a(.in(far_7_7941_0[0]), .out(far_7_7941_1[0]));    relay_conn far_7_7941_1_b(.in(far_7_7941_0[1]), .out(far_7_7941_1[1]));
    wire [1:0] far_7_7941_2;    relay_conn far_7_7941_2_a(.in(far_7_7941_1[0]), .out(far_7_7941_2[0]));    relay_conn far_7_7941_2_b(.in(far_7_7941_1[1]), .out(far_7_7941_2[1]));
    assign out[801] = ~(far_7_7941_2[0] & far_7_7941_2[1]); 
    wire [1:0] far_7_7942_0;    relay_conn far_7_7942_0_a(.in(layer_6[644]), .out(far_7_7942_0[0]));    relay_conn far_7_7942_0_b(.in(layer_6[768]), .out(far_7_7942_0[1]));
    wire [1:0] far_7_7942_1;    relay_conn far_7_7942_1_a(.in(far_7_7942_0[0]), .out(far_7_7942_1[0]));    relay_conn far_7_7942_1_b(.in(far_7_7942_0[1]), .out(far_7_7942_1[1]));
    wire [1:0] far_7_7942_2;    relay_conn far_7_7942_2_a(.in(far_7_7942_1[0]), .out(far_7_7942_2[0]));    relay_conn far_7_7942_2_b(.in(far_7_7942_1[1]), .out(far_7_7942_2[1]));
    assign out[802] = far_7_7942_2[1] & ~far_7_7942_2[0]; 
    wire [1:0] far_7_7943_0;    relay_conn far_7_7943_0_a(.in(layer_6[456]), .out(far_7_7943_0[0]));    relay_conn far_7_7943_0_b(.in(layer_6[561]), .out(far_7_7943_0[1]));
    wire [1:0] far_7_7943_1;    relay_conn far_7_7943_1_a(.in(far_7_7943_0[0]), .out(far_7_7943_1[0]));    relay_conn far_7_7943_1_b(.in(far_7_7943_0[1]), .out(far_7_7943_1[1]));
    wire [1:0] far_7_7943_2;    relay_conn far_7_7943_2_a(.in(far_7_7943_1[0]), .out(far_7_7943_2[0]));    relay_conn far_7_7943_2_b(.in(far_7_7943_1[1]), .out(far_7_7943_2[1]));
    assign out[803] = ~far_7_7943_2[1]; 
    assign out[804] = ~(layer_6[117] | layer_6[96]); 
    wire [1:0] far_7_7945_0;    relay_conn far_7_7945_0_a(.in(layer_6[198]), .out(far_7_7945_0[0]));    relay_conn far_7_7945_0_b(.in(layer_6[157]), .out(far_7_7945_0[1]));
    assign out[805] = far_7_7945_0[0] & ~far_7_7945_0[1]; 
    wire [1:0] far_7_7946_0;    relay_conn far_7_7946_0_a(.in(layer_6[924]), .out(far_7_7946_0[0]));    relay_conn far_7_7946_0_b(.in(layer_6[814]), .out(far_7_7946_0[1]));
    wire [1:0] far_7_7946_1;    relay_conn far_7_7946_1_a(.in(far_7_7946_0[0]), .out(far_7_7946_1[0]));    relay_conn far_7_7946_1_b(.in(far_7_7946_0[1]), .out(far_7_7946_1[1]));
    wire [1:0] far_7_7946_2;    relay_conn far_7_7946_2_a(.in(far_7_7946_1[0]), .out(far_7_7946_2[0]));    relay_conn far_7_7946_2_b(.in(far_7_7946_1[1]), .out(far_7_7946_2[1]));
    assign out[806] = ~(far_7_7946_2[0] ^ far_7_7946_2[1]); 
    wire [1:0] far_7_7947_0;    relay_conn far_7_7947_0_a(.in(layer_6[1016]), .out(far_7_7947_0[0]));    relay_conn far_7_7947_0_b(.in(layer_6[888]), .out(far_7_7947_0[1]));
    wire [1:0] far_7_7947_1;    relay_conn far_7_7947_1_a(.in(far_7_7947_0[0]), .out(far_7_7947_1[0]));    relay_conn far_7_7947_1_b(.in(far_7_7947_0[1]), .out(far_7_7947_1[1]));
    wire [1:0] far_7_7947_2;    relay_conn far_7_7947_2_a(.in(far_7_7947_1[0]), .out(far_7_7947_2[0]));    relay_conn far_7_7947_2_b(.in(far_7_7947_1[1]), .out(far_7_7947_2[1]));
    wire [1:0] far_7_7947_3;    relay_conn far_7_7947_3_a(.in(far_7_7947_2[0]), .out(far_7_7947_3[0]));    relay_conn far_7_7947_3_b(.in(far_7_7947_2[1]), .out(far_7_7947_3[1]));
    assign out[807] = far_7_7947_3[0] & ~far_7_7947_3[1]; 
    wire [1:0] far_7_7948_0;    relay_conn far_7_7948_0_a(.in(layer_6[268]), .out(far_7_7948_0[0]));    relay_conn far_7_7948_0_b(.in(layer_6[320]), .out(far_7_7948_0[1]));
    assign out[808] = far_7_7948_0[0] & far_7_7948_0[1]; 
    assign out[809] = layer_6[575] & ~layer_6[566]; 
    assign out[810] = layer_6[425] & ~layer_6[394]; 
    wire [1:0] far_7_7951_0;    relay_conn far_7_7951_0_a(.in(layer_6[649]), .out(far_7_7951_0[0]));    relay_conn far_7_7951_0_b(.in(layer_6[753]), .out(far_7_7951_0[1]));
    wire [1:0] far_7_7951_1;    relay_conn far_7_7951_1_a(.in(far_7_7951_0[0]), .out(far_7_7951_1[0]));    relay_conn far_7_7951_1_b(.in(far_7_7951_0[1]), .out(far_7_7951_1[1]));
    wire [1:0] far_7_7951_2;    relay_conn far_7_7951_2_a(.in(far_7_7951_1[0]), .out(far_7_7951_2[0]));    relay_conn far_7_7951_2_b(.in(far_7_7951_1[1]), .out(far_7_7951_2[1]));
    assign out[811] = ~far_7_7951_2[1]; 
    wire [1:0] far_7_7952_0;    relay_conn far_7_7952_0_a(.in(layer_6[273]), .out(far_7_7952_0[0]));    relay_conn far_7_7952_0_b(.in(layer_6[238]), .out(far_7_7952_0[1]));
    assign out[812] = ~far_7_7952_0[1]; 
    wire [1:0] far_7_7953_0;    relay_conn far_7_7953_0_a(.in(layer_6[101]), .out(far_7_7953_0[0]));    relay_conn far_7_7953_0_b(.in(layer_6[160]), .out(far_7_7953_0[1]));
    assign out[813] = far_7_7953_0[1] & ~far_7_7953_0[0]; 
    wire [1:0] far_7_7954_0;    relay_conn far_7_7954_0_a(.in(layer_6[236]), .out(far_7_7954_0[0]));    relay_conn far_7_7954_0_b(.in(layer_6[128]), .out(far_7_7954_0[1]));
    wire [1:0] far_7_7954_1;    relay_conn far_7_7954_1_a(.in(far_7_7954_0[0]), .out(far_7_7954_1[0]));    relay_conn far_7_7954_1_b(.in(far_7_7954_0[1]), .out(far_7_7954_1[1]));
    wire [1:0] far_7_7954_2;    relay_conn far_7_7954_2_a(.in(far_7_7954_1[0]), .out(far_7_7954_2[0]));    relay_conn far_7_7954_2_b(.in(far_7_7954_1[1]), .out(far_7_7954_2[1]));
    assign out[814] = ~far_7_7954_2[1]; 
    wire [1:0] far_7_7955_0;    relay_conn far_7_7955_0_a(.in(layer_6[292]), .out(far_7_7955_0[0]));    relay_conn far_7_7955_0_b(.in(layer_6[192]), .out(far_7_7955_0[1]));
    wire [1:0] far_7_7955_1;    relay_conn far_7_7955_1_a(.in(far_7_7955_0[0]), .out(far_7_7955_1[0]));    relay_conn far_7_7955_1_b(.in(far_7_7955_0[1]), .out(far_7_7955_1[1]));
    wire [1:0] far_7_7955_2;    relay_conn far_7_7955_2_a(.in(far_7_7955_1[0]), .out(far_7_7955_2[0]));    relay_conn far_7_7955_2_b(.in(far_7_7955_1[1]), .out(far_7_7955_2[1]));
    assign out[815] = ~far_7_7955_2[0]; 
    wire [1:0] far_7_7956_0;    relay_conn far_7_7956_0_a(.in(layer_6[57]), .out(far_7_7956_0[0]));    relay_conn far_7_7956_0_b(.in(layer_6[128]), .out(far_7_7956_0[1]));
    wire [1:0] far_7_7956_1;    relay_conn far_7_7956_1_a(.in(far_7_7956_0[0]), .out(far_7_7956_1[0]));    relay_conn far_7_7956_1_b(.in(far_7_7956_0[1]), .out(far_7_7956_1[1]));
    assign out[816] = far_7_7956_1[0] & far_7_7956_1[1]; 
    wire [1:0] far_7_7957_0;    relay_conn far_7_7957_0_a(.in(layer_6[906]), .out(far_7_7957_0[0]));    relay_conn far_7_7957_0_b(.in(layer_6[1008]), .out(far_7_7957_0[1]));
    wire [1:0] far_7_7957_1;    relay_conn far_7_7957_1_a(.in(far_7_7957_0[0]), .out(far_7_7957_1[0]));    relay_conn far_7_7957_1_b(.in(far_7_7957_0[1]), .out(far_7_7957_1[1]));
    wire [1:0] far_7_7957_2;    relay_conn far_7_7957_2_a(.in(far_7_7957_1[0]), .out(far_7_7957_2[0]));    relay_conn far_7_7957_2_b(.in(far_7_7957_1[1]), .out(far_7_7957_2[1]));
    assign out[817] = far_7_7957_2[0] & ~far_7_7957_2[1]; 
    wire [1:0] far_7_7958_0;    relay_conn far_7_7958_0_a(.in(layer_6[923]), .out(far_7_7958_0[0]));    relay_conn far_7_7958_0_b(.in(layer_6[859]), .out(far_7_7958_0[1]));
    wire [1:0] far_7_7958_1;    relay_conn far_7_7958_1_a(.in(far_7_7958_0[0]), .out(far_7_7958_1[0]));    relay_conn far_7_7958_1_b(.in(far_7_7958_0[1]), .out(far_7_7958_1[1]));
    assign out[818] = far_7_7958_1[1] & ~far_7_7958_1[0]; 
    wire [1:0] far_7_7959_0;    relay_conn far_7_7959_0_a(.in(layer_6[732]), .out(far_7_7959_0[0]));    relay_conn far_7_7959_0_b(.in(layer_6[774]), .out(far_7_7959_0[1]));
    assign out[819] = far_7_7959_0[0]; 
    assign out[820] = layer_6[345] & ~layer_6[337]; 
    wire [1:0] far_7_7961_0;    relay_conn far_7_7961_0_a(.in(layer_6[369]), .out(far_7_7961_0[0]));    relay_conn far_7_7961_0_b(.in(layer_6[468]), .out(far_7_7961_0[1]));
    wire [1:0] far_7_7961_1;    relay_conn far_7_7961_1_a(.in(far_7_7961_0[0]), .out(far_7_7961_1[0]));    relay_conn far_7_7961_1_b(.in(far_7_7961_0[1]), .out(far_7_7961_1[1]));
    wire [1:0] far_7_7961_2;    relay_conn far_7_7961_2_a(.in(far_7_7961_1[0]), .out(far_7_7961_2[0]));    relay_conn far_7_7961_2_b(.in(far_7_7961_1[1]), .out(far_7_7961_2[1]));
    assign out[821] = far_7_7961_2[0] & ~far_7_7961_2[1]; 
    wire [1:0] far_7_7962_0;    relay_conn far_7_7962_0_a(.in(layer_6[534]), .out(far_7_7962_0[0]));    relay_conn far_7_7962_0_b(.in(layer_6[456]), .out(far_7_7962_0[1]));
    wire [1:0] far_7_7962_1;    relay_conn far_7_7962_1_a(.in(far_7_7962_0[0]), .out(far_7_7962_1[0]));    relay_conn far_7_7962_1_b(.in(far_7_7962_0[1]), .out(far_7_7962_1[1]));
    assign out[822] = far_7_7962_1[0] & far_7_7962_1[1]; 
    wire [1:0] far_7_7963_0;    relay_conn far_7_7963_0_a(.in(layer_6[30]), .out(far_7_7963_0[0]));    relay_conn far_7_7963_0_b(.in(layer_6[127]), .out(far_7_7963_0[1]));
    wire [1:0] far_7_7963_1;    relay_conn far_7_7963_1_a(.in(far_7_7963_0[0]), .out(far_7_7963_1[0]));    relay_conn far_7_7963_1_b(.in(far_7_7963_0[1]), .out(far_7_7963_1[1]));
    wire [1:0] far_7_7963_2;    relay_conn far_7_7963_2_a(.in(far_7_7963_1[0]), .out(far_7_7963_2[0]));    relay_conn far_7_7963_2_b(.in(far_7_7963_1[1]), .out(far_7_7963_2[1]));
    assign out[823] = ~far_7_7963_2[1]; 
    wire [1:0] far_7_7964_0;    relay_conn far_7_7964_0_a(.in(layer_6[583]), .out(far_7_7964_0[0]));    relay_conn far_7_7964_0_b(.in(layer_6[497]), .out(far_7_7964_0[1]));
    wire [1:0] far_7_7964_1;    relay_conn far_7_7964_1_a(.in(far_7_7964_0[0]), .out(far_7_7964_1[0]));    relay_conn far_7_7964_1_b(.in(far_7_7964_0[1]), .out(far_7_7964_1[1]));
    assign out[824] = far_7_7964_1[1] & ~far_7_7964_1[0]; 
    wire [1:0] far_7_7965_0;    relay_conn far_7_7965_0_a(.in(layer_6[786]), .out(far_7_7965_0[0]));    relay_conn far_7_7965_0_b(.in(layer_6[892]), .out(far_7_7965_0[1]));
    wire [1:0] far_7_7965_1;    relay_conn far_7_7965_1_a(.in(far_7_7965_0[0]), .out(far_7_7965_1[0]));    relay_conn far_7_7965_1_b(.in(far_7_7965_0[1]), .out(far_7_7965_1[1]));
    wire [1:0] far_7_7965_2;    relay_conn far_7_7965_2_a(.in(far_7_7965_1[0]), .out(far_7_7965_2[0]));    relay_conn far_7_7965_2_b(.in(far_7_7965_1[1]), .out(far_7_7965_2[1]));
    assign out[825] = ~far_7_7965_2[1]; 
    assign out[826] = ~layer_6[348]; 
    wire [1:0] far_7_7967_0;    relay_conn far_7_7967_0_a(.in(layer_6[63]), .out(far_7_7967_0[0]));    relay_conn far_7_7967_0_b(.in(layer_6[134]), .out(far_7_7967_0[1]));
    wire [1:0] far_7_7967_1;    relay_conn far_7_7967_1_a(.in(far_7_7967_0[0]), .out(far_7_7967_1[0]));    relay_conn far_7_7967_1_b(.in(far_7_7967_0[1]), .out(far_7_7967_1[1]));
    assign out[827] = ~far_7_7967_1[0]; 
    wire [1:0] far_7_7968_0;    relay_conn far_7_7968_0_a(.in(layer_6[196]), .out(far_7_7968_0[0]));    relay_conn far_7_7968_0_b(.in(layer_6[128]), .out(far_7_7968_0[1]));
    wire [1:0] far_7_7968_1;    relay_conn far_7_7968_1_a(.in(far_7_7968_0[0]), .out(far_7_7968_1[0]));    relay_conn far_7_7968_1_b(.in(far_7_7968_0[1]), .out(far_7_7968_1[1]));
    assign out[828] = far_7_7968_1[1] & ~far_7_7968_1[0]; 
    wire [1:0] far_7_7969_0;    relay_conn far_7_7969_0_a(.in(layer_6[799]), .out(far_7_7969_0[0]));    relay_conn far_7_7969_0_b(.in(layer_6[917]), .out(far_7_7969_0[1]));
    wire [1:0] far_7_7969_1;    relay_conn far_7_7969_1_a(.in(far_7_7969_0[0]), .out(far_7_7969_1[0]));    relay_conn far_7_7969_1_b(.in(far_7_7969_0[1]), .out(far_7_7969_1[1]));
    wire [1:0] far_7_7969_2;    relay_conn far_7_7969_2_a(.in(far_7_7969_1[0]), .out(far_7_7969_2[0]));    relay_conn far_7_7969_2_b(.in(far_7_7969_1[1]), .out(far_7_7969_2[1]));
    assign out[829] = far_7_7969_2[1]; 
    assign out[830] = ~layer_6[780]; 
    wire [1:0] far_7_7971_0;    relay_conn far_7_7971_0_a(.in(layer_6[883]), .out(far_7_7971_0[0]));    relay_conn far_7_7971_0_b(.in(layer_6[777]), .out(far_7_7971_0[1]));
    wire [1:0] far_7_7971_1;    relay_conn far_7_7971_1_a(.in(far_7_7971_0[0]), .out(far_7_7971_1[0]));    relay_conn far_7_7971_1_b(.in(far_7_7971_0[1]), .out(far_7_7971_1[1]));
    wire [1:0] far_7_7971_2;    relay_conn far_7_7971_2_a(.in(far_7_7971_1[0]), .out(far_7_7971_2[0]));    relay_conn far_7_7971_2_b(.in(far_7_7971_1[1]), .out(far_7_7971_2[1]));
    assign out[831] = ~far_7_7971_2[0]; 
    wire [1:0] far_7_7972_0;    relay_conn far_7_7972_0_a(.in(layer_6[404]), .out(far_7_7972_0[0]));    relay_conn far_7_7972_0_b(.in(layer_6[464]), .out(far_7_7972_0[1]));
    assign out[832] = far_7_7972_0[0] & ~far_7_7972_0[1]; 
    wire [1:0] far_7_7973_0;    relay_conn far_7_7973_0_a(.in(layer_6[699]), .out(far_7_7973_0[0]));    relay_conn far_7_7973_0_b(.in(layer_6[614]), .out(far_7_7973_0[1]));
    wire [1:0] far_7_7973_1;    relay_conn far_7_7973_1_a(.in(far_7_7973_0[0]), .out(far_7_7973_1[0]));    relay_conn far_7_7973_1_b(.in(far_7_7973_0[1]), .out(far_7_7973_1[1]));
    assign out[833] = ~far_7_7973_1[1]; 
    assign out[834] = layer_6[601]; 
    wire [1:0] far_7_7975_0;    relay_conn far_7_7975_0_a(.in(layer_6[993]), .out(far_7_7975_0[0]));    relay_conn far_7_7975_0_b(.in(layer_6[923]), .out(far_7_7975_0[1]));
    wire [1:0] far_7_7975_1;    relay_conn far_7_7975_1_a(.in(far_7_7975_0[0]), .out(far_7_7975_1[0]));    relay_conn far_7_7975_1_b(.in(far_7_7975_0[1]), .out(far_7_7975_1[1]));
    assign out[835] = ~(far_7_7975_1[0] | far_7_7975_1[1]); 
    wire [1:0] far_7_7976_0;    relay_conn far_7_7976_0_a(.in(layer_6[678]), .out(far_7_7976_0[0]));    relay_conn far_7_7976_0_b(.in(layer_6[779]), .out(far_7_7976_0[1]));
    wire [1:0] far_7_7976_1;    relay_conn far_7_7976_1_a(.in(far_7_7976_0[0]), .out(far_7_7976_1[0]));    relay_conn far_7_7976_1_b(.in(far_7_7976_0[1]), .out(far_7_7976_1[1]));
    wire [1:0] far_7_7976_2;    relay_conn far_7_7976_2_a(.in(far_7_7976_1[0]), .out(far_7_7976_2[0]));    relay_conn far_7_7976_2_b(.in(far_7_7976_1[1]), .out(far_7_7976_2[1]));
    assign out[836] = far_7_7976_2[1] & ~far_7_7976_2[0]; 
    wire [1:0] far_7_7977_0;    relay_conn far_7_7977_0_a(.in(layer_6[387]), .out(far_7_7977_0[0]));    relay_conn far_7_7977_0_b(.in(layer_6[332]), .out(far_7_7977_0[1]));
    assign out[837] = far_7_7977_0[0] & ~far_7_7977_0[1]; 
    assign out[838] = layer_6[667] ^ layer_6[665]; 
    wire [1:0] far_7_7979_0;    relay_conn far_7_7979_0_a(.in(layer_6[916]), .out(far_7_7979_0[0]));    relay_conn far_7_7979_0_b(.in(layer_6[799]), .out(far_7_7979_0[1]));
    wire [1:0] far_7_7979_1;    relay_conn far_7_7979_1_a(.in(far_7_7979_0[0]), .out(far_7_7979_1[0]));    relay_conn far_7_7979_1_b(.in(far_7_7979_0[1]), .out(far_7_7979_1[1]));
    wire [1:0] far_7_7979_2;    relay_conn far_7_7979_2_a(.in(far_7_7979_1[0]), .out(far_7_7979_2[0]));    relay_conn far_7_7979_2_b(.in(far_7_7979_1[1]), .out(far_7_7979_2[1]));
    assign out[839] = ~far_7_7979_2[0]; 
    wire [1:0] far_7_7980_0;    relay_conn far_7_7980_0_a(.in(layer_6[837]), .out(far_7_7980_0[0]));    relay_conn far_7_7980_0_b(.in(layer_6[799]), .out(far_7_7980_0[1]));
    assign out[840] = ~(far_7_7980_0[0] | far_7_7980_0[1]); 
    assign out[841] = layer_6[815] ^ layer_6[794]; 
    wire [1:0] far_7_7982_0;    relay_conn far_7_7982_0_a(.in(layer_6[976]), .out(far_7_7982_0[0]));    relay_conn far_7_7982_0_b(.in(layer_6[1017]), .out(far_7_7982_0[1]));
    assign out[842] = far_7_7982_0[0] & ~far_7_7982_0[1]; 
    wire [1:0] far_7_7983_0;    relay_conn far_7_7983_0_a(.in(layer_6[189]), .out(far_7_7983_0[0]));    relay_conn far_7_7983_0_b(.in(layer_6[267]), .out(far_7_7983_0[1]));
    wire [1:0] far_7_7983_1;    relay_conn far_7_7983_1_a(.in(far_7_7983_0[0]), .out(far_7_7983_1[0]));    relay_conn far_7_7983_1_b(.in(far_7_7983_0[1]), .out(far_7_7983_1[1]));
    assign out[843] = ~(far_7_7983_1[0] ^ far_7_7983_1[1]); 
    assign out[844] = layer_6[788] & layer_6[789]; 
    wire [1:0] far_7_7985_0;    relay_conn far_7_7985_0_a(.in(layer_6[395]), .out(far_7_7985_0[0]));    relay_conn far_7_7985_0_b(.in(layer_6[503]), .out(far_7_7985_0[1]));
    wire [1:0] far_7_7985_1;    relay_conn far_7_7985_1_a(.in(far_7_7985_0[0]), .out(far_7_7985_1[0]));    relay_conn far_7_7985_1_b(.in(far_7_7985_0[1]), .out(far_7_7985_1[1]));
    wire [1:0] far_7_7985_2;    relay_conn far_7_7985_2_a(.in(far_7_7985_1[0]), .out(far_7_7985_2[0]));    relay_conn far_7_7985_2_b(.in(far_7_7985_1[1]), .out(far_7_7985_2[1]));
    assign out[845] = far_7_7985_2[0] & far_7_7985_2[1]; 
    wire [1:0] far_7_7986_0;    relay_conn far_7_7986_0_a(.in(layer_6[831]), .out(far_7_7986_0[0]));    relay_conn far_7_7986_0_b(.in(layer_6[930]), .out(far_7_7986_0[1]));
    wire [1:0] far_7_7986_1;    relay_conn far_7_7986_1_a(.in(far_7_7986_0[0]), .out(far_7_7986_1[0]));    relay_conn far_7_7986_1_b(.in(far_7_7986_0[1]), .out(far_7_7986_1[1]));
    wire [1:0] far_7_7986_2;    relay_conn far_7_7986_2_a(.in(far_7_7986_1[0]), .out(far_7_7986_2[0]));    relay_conn far_7_7986_2_b(.in(far_7_7986_1[1]), .out(far_7_7986_2[1]));
    assign out[846] = far_7_7986_2[0] & ~far_7_7986_2[1]; 
    assign out[847] = layer_6[550] & ~layer_6[523]; 
    wire [1:0] far_7_7988_0;    relay_conn far_7_7988_0_a(.in(layer_6[845]), .out(far_7_7988_0[0]));    relay_conn far_7_7988_0_b(.in(layer_6[778]), .out(far_7_7988_0[1]));
    wire [1:0] far_7_7988_1;    relay_conn far_7_7988_1_a(.in(far_7_7988_0[0]), .out(far_7_7988_1[0]));    relay_conn far_7_7988_1_b(.in(far_7_7988_0[1]), .out(far_7_7988_1[1]));
    assign out[848] = far_7_7988_1[0] & far_7_7988_1[1]; 
    wire [1:0] far_7_7989_0;    relay_conn far_7_7989_0_a(.in(layer_6[718]), .out(far_7_7989_0[0]));    relay_conn far_7_7989_0_b(.in(layer_6[835]), .out(far_7_7989_0[1]));
    wire [1:0] far_7_7989_1;    relay_conn far_7_7989_1_a(.in(far_7_7989_0[0]), .out(far_7_7989_1[0]));    relay_conn far_7_7989_1_b(.in(far_7_7989_0[1]), .out(far_7_7989_1[1]));
    wire [1:0] far_7_7989_2;    relay_conn far_7_7989_2_a(.in(far_7_7989_1[0]), .out(far_7_7989_2[0]));    relay_conn far_7_7989_2_b(.in(far_7_7989_1[1]), .out(far_7_7989_2[1]));
    assign out[849] = far_7_7989_2[1]; 
    wire [1:0] far_7_7990_0;    relay_conn far_7_7990_0_a(.in(layer_6[254]), .out(far_7_7990_0[0]));    relay_conn far_7_7990_0_b(.in(layer_6[192]), .out(far_7_7990_0[1]));
    assign out[850] = ~far_7_7990_0[0]; 
    assign out[851] = layer_6[950]; 
    wire [1:0] far_7_7992_0;    relay_conn far_7_7992_0_a(.in(layer_6[971]), .out(far_7_7992_0[0]));    relay_conn far_7_7992_0_b(.in(layer_6[884]), .out(far_7_7992_0[1]));
    wire [1:0] far_7_7992_1;    relay_conn far_7_7992_1_a(.in(far_7_7992_0[0]), .out(far_7_7992_1[0]));    relay_conn far_7_7992_1_b(.in(far_7_7992_0[1]), .out(far_7_7992_1[1]));
    assign out[852] = far_7_7992_1[0] ^ far_7_7992_1[1]; 
    assign out[853] = layer_6[226] ^ layer_6[227]; 
    wire [1:0] far_7_7994_0;    relay_conn far_7_7994_0_a(.in(layer_6[415]), .out(far_7_7994_0[0]));    relay_conn far_7_7994_0_b(.in(layer_6[469]), .out(far_7_7994_0[1]));
    assign out[854] = far_7_7994_0[0] & ~far_7_7994_0[1]; 
    wire [1:0] far_7_7995_0;    relay_conn far_7_7995_0_a(.in(layer_6[778]), .out(far_7_7995_0[0]));    relay_conn far_7_7995_0_b(.in(layer_6[824]), .out(far_7_7995_0[1]));
    assign out[855] = far_7_7995_0[0]; 
    wire [1:0] far_7_7996_0;    relay_conn far_7_7996_0_a(.in(layer_6[120]), .out(far_7_7996_0[0]));    relay_conn far_7_7996_0_b(.in(layer_6[66]), .out(far_7_7996_0[1]));
    assign out[856] = ~far_7_7996_0[1]; 
    wire [1:0] far_7_7997_0;    relay_conn far_7_7997_0_a(.in(layer_6[773]), .out(far_7_7997_0[0]));    relay_conn far_7_7997_0_b(.in(layer_6[839]), .out(far_7_7997_0[1]));
    wire [1:0] far_7_7997_1;    relay_conn far_7_7997_1_a(.in(far_7_7997_0[0]), .out(far_7_7997_1[0]));    relay_conn far_7_7997_1_b(.in(far_7_7997_0[1]), .out(far_7_7997_1[1]));
    assign out[857] = far_7_7997_1[1]; 
    wire [1:0] far_7_7998_0;    relay_conn far_7_7998_0_a(.in(layer_6[799]), .out(far_7_7998_0[0]));    relay_conn far_7_7998_0_b(.in(layer_6[870]), .out(far_7_7998_0[1]));
    wire [1:0] far_7_7998_1;    relay_conn far_7_7998_1_a(.in(far_7_7998_0[0]), .out(far_7_7998_1[0]));    relay_conn far_7_7998_1_b(.in(far_7_7998_0[1]), .out(far_7_7998_1[1]));
    assign out[858] = far_7_7998_1[1] & ~far_7_7998_1[0]; 
    wire [1:0] far_7_7999_0;    relay_conn far_7_7999_0_a(.in(layer_6[396]), .out(far_7_7999_0[0]));    relay_conn far_7_7999_0_b(.in(layer_6[497]), .out(far_7_7999_0[1]));
    wire [1:0] far_7_7999_1;    relay_conn far_7_7999_1_a(.in(far_7_7999_0[0]), .out(far_7_7999_1[0]));    relay_conn far_7_7999_1_b(.in(far_7_7999_0[1]), .out(far_7_7999_1[1]));
    wire [1:0] far_7_7999_2;    relay_conn far_7_7999_2_a(.in(far_7_7999_1[0]), .out(far_7_7999_2[0]));    relay_conn far_7_7999_2_b(.in(far_7_7999_1[1]), .out(far_7_7999_2[1]));
    assign out[859] = far_7_7999_2[0] & far_7_7999_2[1]; 
    assign out[860] = ~layer_6[916]; 
    wire [1:0] far_7_8001_0;    relay_conn far_7_8001_0_a(.in(layer_6[470]), .out(far_7_8001_0[0]));    relay_conn far_7_8001_0_b(.in(layer_6[393]), .out(far_7_8001_0[1]));
    wire [1:0] far_7_8001_1;    relay_conn far_7_8001_1_a(.in(far_7_8001_0[0]), .out(far_7_8001_1[0]));    relay_conn far_7_8001_1_b(.in(far_7_8001_0[1]), .out(far_7_8001_1[1]));
    assign out[861] = ~(far_7_8001_1[0] ^ far_7_8001_1[1]); 
    wire [1:0] far_7_8002_0;    relay_conn far_7_8002_0_a(.in(layer_6[226]), .out(far_7_8002_0[0]));    relay_conn far_7_8002_0_b(.in(layer_6[339]), .out(far_7_8002_0[1]));
    wire [1:0] far_7_8002_1;    relay_conn far_7_8002_1_a(.in(far_7_8002_0[0]), .out(far_7_8002_1[0]));    relay_conn far_7_8002_1_b(.in(far_7_8002_0[1]), .out(far_7_8002_1[1]));
    wire [1:0] far_7_8002_2;    relay_conn far_7_8002_2_a(.in(far_7_8002_1[0]), .out(far_7_8002_2[0]));    relay_conn far_7_8002_2_b(.in(far_7_8002_1[1]), .out(far_7_8002_2[1]));
    assign out[862] = far_7_8002_2[1]; 
    wire [1:0] far_7_8003_0;    relay_conn far_7_8003_0_a(.in(layer_6[428]), .out(far_7_8003_0[0]));    relay_conn far_7_8003_0_b(.in(layer_6[503]), .out(far_7_8003_0[1]));
    wire [1:0] far_7_8003_1;    relay_conn far_7_8003_1_a(.in(far_7_8003_0[0]), .out(far_7_8003_1[0]));    relay_conn far_7_8003_1_b(.in(far_7_8003_0[1]), .out(far_7_8003_1[1]));
    assign out[863] = ~far_7_8003_1[0]; 
    wire [1:0] far_7_8004_0;    relay_conn far_7_8004_0_a(.in(layer_6[737]), .out(far_7_8004_0[0]));    relay_conn far_7_8004_0_b(.in(layer_6[793]), .out(far_7_8004_0[1]));
    assign out[864] = far_7_8004_0[0] & ~far_7_8004_0[1]; 
    wire [1:0] far_7_8005_0;    relay_conn far_7_8005_0_a(.in(layer_6[952]), .out(far_7_8005_0[0]));    relay_conn far_7_8005_0_b(.in(layer_6[845]), .out(far_7_8005_0[1]));
    wire [1:0] far_7_8005_1;    relay_conn far_7_8005_1_a(.in(far_7_8005_0[0]), .out(far_7_8005_1[0]));    relay_conn far_7_8005_1_b(.in(far_7_8005_0[1]), .out(far_7_8005_1[1]));
    wire [1:0] far_7_8005_2;    relay_conn far_7_8005_2_a(.in(far_7_8005_1[0]), .out(far_7_8005_2[0]));    relay_conn far_7_8005_2_b(.in(far_7_8005_1[1]), .out(far_7_8005_2[1]));
    assign out[865] = far_7_8005_2[0] ^ far_7_8005_2[1]; 
    wire [1:0] far_7_8006_0;    relay_conn far_7_8006_0_a(.in(layer_6[721]), .out(far_7_8006_0[0]));    relay_conn far_7_8006_0_b(.in(layer_6[678]), .out(far_7_8006_0[1]));
    assign out[866] = far_7_8006_0[0] & ~far_7_8006_0[1]; 
    wire [1:0] far_7_8007_0;    relay_conn far_7_8007_0_a(.in(layer_6[229]), .out(far_7_8007_0[0]));    relay_conn far_7_8007_0_b(.in(layer_6[126]), .out(far_7_8007_0[1]));
    wire [1:0] far_7_8007_1;    relay_conn far_7_8007_1_a(.in(far_7_8007_0[0]), .out(far_7_8007_1[0]));    relay_conn far_7_8007_1_b(.in(far_7_8007_0[1]), .out(far_7_8007_1[1]));
    wire [1:0] far_7_8007_2;    relay_conn far_7_8007_2_a(.in(far_7_8007_1[0]), .out(far_7_8007_2[0]));    relay_conn far_7_8007_2_b(.in(far_7_8007_1[1]), .out(far_7_8007_2[1]));
    assign out[867] = ~(far_7_8007_2[0] | far_7_8007_2[1]); 
    wire [1:0] far_7_8008_0;    relay_conn far_7_8008_0_a(.in(layer_6[899]), .out(far_7_8008_0[0]));    relay_conn far_7_8008_0_b(.in(layer_6[947]), .out(far_7_8008_0[1]));
    assign out[868] = far_7_8008_0[0]; 
    wire [1:0] far_7_8009_0;    relay_conn far_7_8009_0_a(.in(layer_6[51]), .out(far_7_8009_0[0]));    relay_conn far_7_8009_0_b(.in(layer_6[119]), .out(far_7_8009_0[1]));
    wire [1:0] far_7_8009_1;    relay_conn far_7_8009_1_a(.in(far_7_8009_0[0]), .out(far_7_8009_1[0]));    relay_conn far_7_8009_1_b(.in(far_7_8009_0[1]), .out(far_7_8009_1[1]));
    assign out[869] = ~far_7_8009_1[0]; 
    assign out[870] = ~(layer_6[173] | layer_6[171]); 
    wire [1:0] far_7_8011_0;    relay_conn far_7_8011_0_a(.in(layer_6[789]), .out(far_7_8011_0[0]));    relay_conn far_7_8011_0_b(.in(layer_6[704]), .out(far_7_8011_0[1]));
    wire [1:0] far_7_8011_1;    relay_conn far_7_8011_1_a(.in(far_7_8011_0[0]), .out(far_7_8011_1[0]));    relay_conn far_7_8011_1_b(.in(far_7_8011_0[1]), .out(far_7_8011_1[1]));
    assign out[871] = far_7_8011_1[1]; 
    wire [1:0] far_7_8012_0;    relay_conn far_7_8012_0_a(.in(layer_6[281]), .out(far_7_8012_0[0]));    relay_conn far_7_8012_0_b(.in(layer_6[219]), .out(far_7_8012_0[1]));
    assign out[872] = far_7_8012_0[0] & ~far_7_8012_0[1]; 
    wire [1:0] far_7_8013_0;    relay_conn far_7_8013_0_a(.in(layer_6[595]), .out(far_7_8013_0[0]));    relay_conn far_7_8013_0_b(.in(layer_6[517]), .out(far_7_8013_0[1]));
    wire [1:0] far_7_8013_1;    relay_conn far_7_8013_1_a(.in(far_7_8013_0[0]), .out(far_7_8013_1[0]));    relay_conn far_7_8013_1_b(.in(far_7_8013_0[1]), .out(far_7_8013_1[1]));
    assign out[873] = ~(far_7_8013_1[0] | far_7_8013_1[1]); 
    wire [1:0] far_7_8014_0;    relay_conn far_7_8014_0_a(.in(layer_6[71]), .out(far_7_8014_0[0]));    relay_conn far_7_8014_0_b(.in(layer_6[197]), .out(far_7_8014_0[1]));
    wire [1:0] far_7_8014_1;    relay_conn far_7_8014_1_a(.in(far_7_8014_0[0]), .out(far_7_8014_1[0]));    relay_conn far_7_8014_1_b(.in(far_7_8014_0[1]), .out(far_7_8014_1[1]));
    wire [1:0] far_7_8014_2;    relay_conn far_7_8014_2_a(.in(far_7_8014_1[0]), .out(far_7_8014_2[0]));    relay_conn far_7_8014_2_b(.in(far_7_8014_1[1]), .out(far_7_8014_2[1]));
    assign out[874] = far_7_8014_2[0] & far_7_8014_2[1]; 
    wire [1:0] far_7_8015_0;    relay_conn far_7_8015_0_a(.in(layer_6[499]), .out(far_7_8015_0[0]));    relay_conn far_7_8015_0_b(.in(layer_6[453]), .out(far_7_8015_0[1]));
    assign out[875] = ~far_7_8015_0[0]; 
    wire [1:0] far_7_8016_0;    relay_conn far_7_8016_0_a(.in(layer_6[459]), .out(far_7_8016_0[0]));    relay_conn far_7_8016_0_b(.in(layer_6[404]), .out(far_7_8016_0[1]));
    assign out[876] = ~far_7_8016_0[0]; 
    wire [1:0] far_7_8017_0;    relay_conn far_7_8017_0_a(.in(layer_6[478]), .out(far_7_8017_0[0]));    relay_conn far_7_8017_0_b(.in(layer_6[391]), .out(far_7_8017_0[1]));
    wire [1:0] far_7_8017_1;    relay_conn far_7_8017_1_a(.in(far_7_8017_0[0]), .out(far_7_8017_1[0]));    relay_conn far_7_8017_1_b(.in(far_7_8017_0[1]), .out(far_7_8017_1[1]));
    assign out[877] = ~(far_7_8017_1[0] ^ far_7_8017_1[1]); 
    assign out[878] = ~layer_6[42] | (layer_6[42] & layer_6[19]); 
    assign out[879] = ~layer_6[199]; 
    assign out[880] = ~(layer_6[585] ^ layer_6[605]); 
    assign out[881] = layer_6[421] & ~layer_6[429]; 
    wire [1:0] far_7_8022_0;    relay_conn far_7_8022_0_a(.in(layer_6[678]), .out(far_7_8022_0[0]));    relay_conn far_7_8022_0_b(.in(layer_6[614]), .out(far_7_8022_0[1]));
    wire [1:0] far_7_8022_1;    relay_conn far_7_8022_1_a(.in(far_7_8022_0[0]), .out(far_7_8022_1[0]));    relay_conn far_7_8022_1_b(.in(far_7_8022_0[1]), .out(far_7_8022_1[1]));
    assign out[882] = ~far_7_8022_1[0]; 
    assign out[883] = layer_6[128]; 
    wire [1:0] far_7_8024_0;    relay_conn far_7_8024_0_a(.in(layer_6[418]), .out(far_7_8024_0[0]));    relay_conn far_7_8024_0_b(.in(layer_6[310]), .out(far_7_8024_0[1]));
    wire [1:0] far_7_8024_1;    relay_conn far_7_8024_1_a(.in(far_7_8024_0[0]), .out(far_7_8024_1[0]));    relay_conn far_7_8024_1_b(.in(far_7_8024_0[1]), .out(far_7_8024_1[1]));
    wire [1:0] far_7_8024_2;    relay_conn far_7_8024_2_a(.in(far_7_8024_1[0]), .out(far_7_8024_2[0]));    relay_conn far_7_8024_2_b(.in(far_7_8024_1[1]), .out(far_7_8024_2[1]));
    assign out[884] = ~far_7_8024_2[0]; 
    wire [1:0] far_7_8025_0;    relay_conn far_7_8025_0_a(.in(layer_6[198]), .out(far_7_8025_0[0]));    relay_conn far_7_8025_0_b(.in(layer_6[101]), .out(far_7_8025_0[1]));
    wire [1:0] far_7_8025_1;    relay_conn far_7_8025_1_a(.in(far_7_8025_0[0]), .out(far_7_8025_1[0]));    relay_conn far_7_8025_1_b(.in(far_7_8025_0[1]), .out(far_7_8025_1[1]));
    wire [1:0] far_7_8025_2;    relay_conn far_7_8025_2_a(.in(far_7_8025_1[0]), .out(far_7_8025_2[0]));    relay_conn far_7_8025_2_b(.in(far_7_8025_1[1]), .out(far_7_8025_2[1]));
    assign out[885] = ~far_7_8025_2[1]; 
    wire [1:0] far_7_8026_0;    relay_conn far_7_8026_0_a(.in(layer_6[715]), .out(far_7_8026_0[0]));    relay_conn far_7_8026_0_b(.in(layer_6[652]), .out(far_7_8026_0[1]));
    assign out[886] = ~far_7_8026_0[0]; 
    wire [1:0] far_7_8027_0;    relay_conn far_7_8027_0_a(.in(layer_6[191]), .out(far_7_8027_0[0]));    relay_conn far_7_8027_0_b(.in(layer_6[260]), .out(far_7_8027_0[1]));
    wire [1:0] far_7_8027_1;    relay_conn far_7_8027_1_a(.in(far_7_8027_0[0]), .out(far_7_8027_1[0]));    relay_conn far_7_8027_1_b(.in(far_7_8027_0[1]), .out(far_7_8027_1[1]));
    assign out[887] = ~far_7_8027_1[0]; 
    wire [1:0] far_7_8028_0;    relay_conn far_7_8028_0_a(.in(layer_6[821]), .out(far_7_8028_0[0]));    relay_conn far_7_8028_0_b(.in(layer_6[737]), .out(far_7_8028_0[1]));
    wire [1:0] far_7_8028_1;    relay_conn far_7_8028_1_a(.in(far_7_8028_0[0]), .out(far_7_8028_1[0]));    relay_conn far_7_8028_1_b(.in(far_7_8028_0[1]), .out(far_7_8028_1[1]));
    assign out[888] = far_7_8028_1[1] & ~far_7_8028_1[0]; 
    wire [1:0] far_7_8029_0;    relay_conn far_7_8029_0_a(.in(layer_6[440]), .out(far_7_8029_0[0]));    relay_conn far_7_8029_0_b(.in(layer_6[387]), .out(far_7_8029_0[1]));
    assign out[889] = far_7_8029_0[1]; 
    wire [1:0] far_7_8030_0;    relay_conn far_7_8030_0_a(.in(layer_6[317]), .out(far_7_8030_0[0]));    relay_conn far_7_8030_0_b(.in(layer_6[353]), .out(far_7_8030_0[1]));
    assign out[890] = far_7_8030_0[0] & ~far_7_8030_0[1]; 
    assign out[891] = ~(layer_6[916] ^ layer_6[896]); 
    assign out[892] = ~(layer_6[764] | layer_6[777]); 
    wire [1:0] far_7_8033_0;    relay_conn far_7_8033_0_a(.in(layer_6[599]), .out(far_7_8033_0[0]));    relay_conn far_7_8033_0_b(.in(layer_6[681]), .out(far_7_8033_0[1]));
    wire [1:0] far_7_8033_1;    relay_conn far_7_8033_1_a(.in(far_7_8033_0[0]), .out(far_7_8033_1[0]));    relay_conn far_7_8033_1_b(.in(far_7_8033_0[1]), .out(far_7_8033_1[1]));
    assign out[893] = ~far_7_8033_1[1]; 
    wire [1:0] far_7_8034_0;    relay_conn far_7_8034_0_a(.in(layer_6[835]), .out(far_7_8034_0[0]));    relay_conn far_7_8034_0_b(.in(layer_6[931]), .out(far_7_8034_0[1]));
    wire [1:0] far_7_8034_1;    relay_conn far_7_8034_1_a(.in(far_7_8034_0[0]), .out(far_7_8034_1[0]));    relay_conn far_7_8034_1_b(.in(far_7_8034_0[1]), .out(far_7_8034_1[1]));
    wire [1:0] far_7_8034_2;    relay_conn far_7_8034_2_a(.in(far_7_8034_1[0]), .out(far_7_8034_2[0]));    relay_conn far_7_8034_2_b(.in(far_7_8034_1[1]), .out(far_7_8034_2[1]));
    assign out[894] = far_7_8034_2[0]; 
    wire [1:0] far_7_8035_0;    relay_conn far_7_8035_0_a(.in(layer_6[702]), .out(far_7_8035_0[0]));    relay_conn far_7_8035_0_b(.in(layer_6[743]), .out(far_7_8035_0[1]));
    assign out[895] = far_7_8035_0[0] & ~far_7_8035_0[1]; 
    assign out[896] = ~(layer_6[312] | layer_6[297]); 
    wire [1:0] far_7_8037_0;    relay_conn far_7_8037_0_a(.in(layer_6[732]), .out(far_7_8037_0[0]));    relay_conn far_7_8037_0_b(.in(layer_6[678]), .out(far_7_8037_0[1]));
    assign out[897] = ~far_7_8037_0[1]; 
    wire [1:0] far_7_8038_0;    relay_conn far_7_8038_0_a(.in(layer_6[923]), .out(far_7_8038_0[0]));    relay_conn far_7_8038_0_b(.in(layer_6[989]), .out(far_7_8038_0[1]));
    wire [1:0] far_7_8038_1;    relay_conn far_7_8038_1_a(.in(far_7_8038_0[0]), .out(far_7_8038_1[0]));    relay_conn far_7_8038_1_b(.in(far_7_8038_0[1]), .out(far_7_8038_1[1]));
    assign out[898] = far_7_8038_1[1]; 
    wire [1:0] far_7_8039_0;    relay_conn far_7_8039_0_a(.in(layer_6[320]), .out(far_7_8039_0[0]));    relay_conn far_7_8039_0_b(.in(layer_6[392]), .out(far_7_8039_0[1]));
    wire [1:0] far_7_8039_1;    relay_conn far_7_8039_1_a(.in(far_7_8039_0[0]), .out(far_7_8039_1[0]));    relay_conn far_7_8039_1_b(.in(far_7_8039_0[1]), .out(far_7_8039_1[1]));
    assign out[899] = ~(far_7_8039_1[0] | far_7_8039_1[1]); 
    wire [1:0] far_7_8040_0;    relay_conn far_7_8040_0_a(.in(layer_6[387]), .out(far_7_8040_0[0]));    relay_conn far_7_8040_0_b(.in(layer_6[449]), .out(far_7_8040_0[1]));
    assign out[900] = far_7_8040_0[0] & ~far_7_8040_0[1]; 
    wire [1:0] far_7_8041_0;    relay_conn far_7_8041_0_a(.in(layer_6[350]), .out(far_7_8041_0[0]));    relay_conn far_7_8041_0_b(.in(layer_6[425]), .out(far_7_8041_0[1]));
    wire [1:0] far_7_8041_1;    relay_conn far_7_8041_1_a(.in(far_7_8041_0[0]), .out(far_7_8041_1[0]));    relay_conn far_7_8041_1_b(.in(far_7_8041_0[1]), .out(far_7_8041_1[1]));
    assign out[901] = far_7_8041_1[0] & far_7_8041_1[1]; 
    wire [1:0] far_7_8042_0;    relay_conn far_7_8042_0_a(.in(layer_6[60]), .out(far_7_8042_0[0]));    relay_conn far_7_8042_0_b(.in(layer_6[151]), .out(far_7_8042_0[1]));
    wire [1:0] far_7_8042_1;    relay_conn far_7_8042_1_a(.in(far_7_8042_0[0]), .out(far_7_8042_1[0]));    relay_conn far_7_8042_1_b(.in(far_7_8042_0[1]), .out(far_7_8042_1[1]));
    assign out[902] = far_7_8042_1[0] & far_7_8042_1[1]; 
    assign out[903] = layer_6[372] & ~layer_6[381]; 
    wire [1:0] far_7_8044_0;    relay_conn far_7_8044_0_a(.in(layer_6[910]), .out(far_7_8044_0[0]));    relay_conn far_7_8044_0_b(.in(layer_6[819]), .out(far_7_8044_0[1]));
    wire [1:0] far_7_8044_1;    relay_conn far_7_8044_1_a(.in(far_7_8044_0[0]), .out(far_7_8044_1[0]));    relay_conn far_7_8044_1_b(.in(far_7_8044_0[1]), .out(far_7_8044_1[1]));
    assign out[904] = far_7_8044_1[1] & ~far_7_8044_1[0]; 
    wire [1:0] far_7_8045_0;    relay_conn far_7_8045_0_a(.in(layer_6[470]), .out(far_7_8045_0[0]));    relay_conn far_7_8045_0_b(.in(layer_6[582]), .out(far_7_8045_0[1]));
    wire [1:0] far_7_8045_1;    relay_conn far_7_8045_1_a(.in(far_7_8045_0[0]), .out(far_7_8045_1[0]));    relay_conn far_7_8045_1_b(.in(far_7_8045_0[1]), .out(far_7_8045_1[1]));
    wire [1:0] far_7_8045_2;    relay_conn far_7_8045_2_a(.in(far_7_8045_1[0]), .out(far_7_8045_2[0]));    relay_conn far_7_8045_2_b(.in(far_7_8045_1[1]), .out(far_7_8045_2[1]));
    assign out[905] = far_7_8045_2[0] & ~far_7_8045_2[1]; 
    wire [1:0] far_7_8046_0;    relay_conn far_7_8046_0_a(.in(layer_6[510]), .out(far_7_8046_0[0]));    relay_conn far_7_8046_0_b(.in(layer_6[478]), .out(far_7_8046_0[1]));
    assign out[906] = far_7_8046_0[1] & ~far_7_8046_0[0]; 
    assign out[907] = ~layer_6[35]; 
    assign out[908] = layer_6[151]; 
    wire [1:0] far_7_8049_0;    relay_conn far_7_8049_0_a(.in(layer_6[605]), .out(far_7_8049_0[0]));    relay_conn far_7_8049_0_b(.in(layer_6[651]), .out(far_7_8049_0[1]));
    assign out[909] = ~far_7_8049_0[1] | (far_7_8049_0[0] & far_7_8049_0[1]); 
    wire [1:0] far_7_8050_0;    relay_conn far_7_8050_0_a(.in(layer_6[629]), .out(far_7_8050_0[0]));    relay_conn far_7_8050_0_b(.in(layer_6[512]), .out(far_7_8050_0[1]));
    wire [1:0] far_7_8050_1;    relay_conn far_7_8050_1_a(.in(far_7_8050_0[0]), .out(far_7_8050_1[0]));    relay_conn far_7_8050_1_b(.in(far_7_8050_0[1]), .out(far_7_8050_1[1]));
    wire [1:0] far_7_8050_2;    relay_conn far_7_8050_2_a(.in(far_7_8050_1[0]), .out(far_7_8050_2[0]));    relay_conn far_7_8050_2_b(.in(far_7_8050_1[1]), .out(far_7_8050_2[1]));
    assign out[910] = ~(far_7_8050_2[0] | far_7_8050_2[1]); 
    wire [1:0] far_7_8051_0;    relay_conn far_7_8051_0_a(.in(layer_6[665]), .out(far_7_8051_0[0]));    relay_conn far_7_8051_0_b(.in(layer_6[700]), .out(far_7_8051_0[1]));
    assign out[911] = far_7_8051_0[1]; 
    wire [1:0] far_7_8052_0;    relay_conn far_7_8052_0_a(.in(layer_6[165]), .out(far_7_8052_0[0]));    relay_conn far_7_8052_0_b(.in(layer_6[219]), .out(far_7_8052_0[1]));
    assign out[912] = ~(far_7_8052_0[0] | far_7_8052_0[1]); 
    wire [1:0] far_7_8053_0;    relay_conn far_7_8053_0_a(.in(layer_6[359]), .out(far_7_8053_0[0]));    relay_conn far_7_8053_0_b(.in(layer_6[451]), .out(far_7_8053_0[1]));
    wire [1:0] far_7_8053_1;    relay_conn far_7_8053_1_a(.in(far_7_8053_0[0]), .out(far_7_8053_1[0]));    relay_conn far_7_8053_1_b(.in(far_7_8053_0[1]), .out(far_7_8053_1[1]));
    assign out[913] = ~far_7_8053_1[0]; 
    assign out[914] = layer_6[524]; 
    wire [1:0] far_7_8055_0;    relay_conn far_7_8055_0_a(.in(layer_6[873]), .out(far_7_8055_0[0]));    relay_conn far_7_8055_0_b(.in(layer_6[792]), .out(far_7_8055_0[1]));
    wire [1:0] far_7_8055_1;    relay_conn far_7_8055_1_a(.in(far_7_8055_0[0]), .out(far_7_8055_1[0]));    relay_conn far_7_8055_1_b(.in(far_7_8055_0[1]), .out(far_7_8055_1[1]));
    assign out[915] = far_7_8055_1[0] & ~far_7_8055_1[1]; 
    wire [1:0] far_7_8056_0;    relay_conn far_7_8056_0_a(.in(layer_6[597]), .out(far_7_8056_0[0]));    relay_conn far_7_8056_0_b(.in(layer_6[688]), .out(far_7_8056_0[1]));
    wire [1:0] far_7_8056_1;    relay_conn far_7_8056_1_a(.in(far_7_8056_0[0]), .out(far_7_8056_1[0]));    relay_conn far_7_8056_1_b(.in(far_7_8056_0[1]), .out(far_7_8056_1[1]));
    assign out[916] = far_7_8056_1[1]; 
    assign out[917] = layer_6[917]; 
    wire [1:0] far_7_8058_0;    relay_conn far_7_8058_0_a(.in(layer_6[526]), .out(far_7_8058_0[0]));    relay_conn far_7_8058_0_b(.in(layer_6[596]), .out(far_7_8058_0[1]));
    wire [1:0] far_7_8058_1;    relay_conn far_7_8058_1_a(.in(far_7_8058_0[0]), .out(far_7_8058_1[0]));    relay_conn far_7_8058_1_b(.in(far_7_8058_0[1]), .out(far_7_8058_1[1]));
    assign out[918] = ~far_7_8058_1[1]; 
    wire [1:0] far_7_8059_0;    relay_conn far_7_8059_0_a(.in(layer_6[944]), .out(far_7_8059_0[0]));    relay_conn far_7_8059_0_b(.in(layer_6[1018]), .out(far_7_8059_0[1]));
    wire [1:0] far_7_8059_1;    relay_conn far_7_8059_1_a(.in(far_7_8059_0[0]), .out(far_7_8059_1[0]));    relay_conn far_7_8059_1_b(.in(far_7_8059_0[1]), .out(far_7_8059_1[1]));
    assign out[919] = far_7_8059_1[1]; 
    wire [1:0] far_7_8060_0;    relay_conn far_7_8060_0_a(.in(layer_6[659]), .out(far_7_8060_0[0]));    relay_conn far_7_8060_0_b(.in(layer_6[539]), .out(far_7_8060_0[1]));
    wire [1:0] far_7_8060_1;    relay_conn far_7_8060_1_a(.in(far_7_8060_0[0]), .out(far_7_8060_1[0]));    relay_conn far_7_8060_1_b(.in(far_7_8060_0[1]), .out(far_7_8060_1[1]));
    wire [1:0] far_7_8060_2;    relay_conn far_7_8060_2_a(.in(far_7_8060_1[0]), .out(far_7_8060_2[0]));    relay_conn far_7_8060_2_b(.in(far_7_8060_1[1]), .out(far_7_8060_2[1]));
    assign out[920] = ~far_7_8060_2[0]; 
    assign out[921] = layer_6[765] & ~layer_6[769]; 
    assign out[922] = ~layer_6[859]; 
    assign out[923] = ~(layer_6[118] | layer_6[94]); 
    wire [1:0] far_7_8064_0;    relay_conn far_7_8064_0_a(.in(layer_6[71]), .out(far_7_8064_0[0]));    relay_conn far_7_8064_0_b(.in(layer_6[19]), .out(far_7_8064_0[1]));
    assign out[924] = ~far_7_8064_0[1]; 
    wire [1:0] far_7_8065_0;    relay_conn far_7_8065_0_a(.in(layer_6[210]), .out(far_7_8065_0[0]));    relay_conn far_7_8065_0_b(.in(layer_6[141]), .out(far_7_8065_0[1]));
    wire [1:0] far_7_8065_1;    relay_conn far_7_8065_1_a(.in(far_7_8065_0[0]), .out(far_7_8065_1[0]));    relay_conn far_7_8065_1_b(.in(far_7_8065_0[1]), .out(far_7_8065_1[1]));
    assign out[925] = far_7_8065_1[0] ^ far_7_8065_1[1]; 
    wire [1:0] far_7_8066_0;    relay_conn far_7_8066_0_a(.in(layer_6[634]), .out(far_7_8066_0[0]));    relay_conn far_7_8066_0_b(.in(layer_6[720]), .out(far_7_8066_0[1]));
    wire [1:0] far_7_8066_1;    relay_conn far_7_8066_1_a(.in(far_7_8066_0[0]), .out(far_7_8066_1[0]));    relay_conn far_7_8066_1_b(.in(far_7_8066_0[1]), .out(far_7_8066_1[1]));
    assign out[926] = far_7_8066_1[0] & far_7_8066_1[1]; 
    wire [1:0] far_7_8067_0;    relay_conn far_7_8067_0_a(.in(layer_6[229]), .out(far_7_8067_0[0]));    relay_conn far_7_8067_0_b(.in(layer_6[163]), .out(far_7_8067_0[1]));
    wire [1:0] far_7_8067_1;    relay_conn far_7_8067_1_a(.in(far_7_8067_0[0]), .out(far_7_8067_1[0]));    relay_conn far_7_8067_1_b(.in(far_7_8067_0[1]), .out(far_7_8067_1[1]));
    assign out[927] = far_7_8067_1[0] & far_7_8067_1[1]; 
    wire [1:0] far_7_8068_0;    relay_conn far_7_8068_0_a(.in(layer_6[995]), .out(far_7_8068_0[0]));    relay_conn far_7_8068_0_b(.in(layer_6[895]), .out(far_7_8068_0[1]));
    wire [1:0] far_7_8068_1;    relay_conn far_7_8068_1_a(.in(far_7_8068_0[0]), .out(far_7_8068_1[0]));    relay_conn far_7_8068_1_b(.in(far_7_8068_0[1]), .out(far_7_8068_1[1]));
    wire [1:0] far_7_8068_2;    relay_conn far_7_8068_2_a(.in(far_7_8068_1[0]), .out(far_7_8068_2[0]));    relay_conn far_7_8068_2_b(.in(far_7_8068_1[1]), .out(far_7_8068_2[1]));
    assign out[928] = ~far_7_8068_2[0]; 
    assign out[929] = layer_6[320]; 
    wire [1:0] far_7_8070_0;    relay_conn far_7_8070_0_a(.in(layer_6[479]), .out(far_7_8070_0[0]));    relay_conn far_7_8070_0_b(.in(layer_6[513]), .out(far_7_8070_0[1]));
    assign out[930] = far_7_8070_0[0] & far_7_8070_0[1]; 
    assign out[931] = layer_6[48] & layer_6[74]; 
    wire [1:0] far_7_8072_0;    relay_conn far_7_8072_0_a(.in(layer_6[845]), .out(far_7_8072_0[0]));    relay_conn far_7_8072_0_b(.in(layer_6[971]), .out(far_7_8072_0[1]));
    wire [1:0] far_7_8072_1;    relay_conn far_7_8072_1_a(.in(far_7_8072_0[0]), .out(far_7_8072_1[0]));    relay_conn far_7_8072_1_b(.in(far_7_8072_0[1]), .out(far_7_8072_1[1]));
    wire [1:0] far_7_8072_2;    relay_conn far_7_8072_2_a(.in(far_7_8072_1[0]), .out(far_7_8072_2[0]));    relay_conn far_7_8072_2_b(.in(far_7_8072_1[1]), .out(far_7_8072_2[1]));
    assign out[932] = far_7_8072_2[0] & far_7_8072_2[1]; 
    wire [1:0] far_7_8073_0;    relay_conn far_7_8073_0_a(.in(layer_6[456]), .out(far_7_8073_0[0]));    relay_conn far_7_8073_0_b(.in(layer_6[388]), .out(far_7_8073_0[1]));
    wire [1:0] far_7_8073_1;    relay_conn far_7_8073_1_a(.in(far_7_8073_0[0]), .out(far_7_8073_1[0]));    relay_conn far_7_8073_1_b(.in(far_7_8073_0[1]), .out(far_7_8073_1[1]));
    assign out[933] = ~(far_7_8073_1[0] | far_7_8073_1[1]); 
    wire [1:0] far_7_8074_0;    relay_conn far_7_8074_0_a(.in(layer_6[198]), .out(far_7_8074_0[0]));    relay_conn far_7_8074_0_b(.in(layer_6[267]), .out(far_7_8074_0[1]));
    wire [1:0] far_7_8074_1;    relay_conn far_7_8074_1_a(.in(far_7_8074_0[0]), .out(far_7_8074_1[0]));    relay_conn far_7_8074_1_b(.in(far_7_8074_0[1]), .out(far_7_8074_1[1]));
    assign out[934] = far_7_8074_1[0] & ~far_7_8074_1[1]; 
    wire [1:0] far_7_8075_0;    relay_conn far_7_8075_0_a(.in(layer_6[819]), .out(far_7_8075_0[0]));    relay_conn far_7_8075_0_b(.in(layer_6[746]), .out(far_7_8075_0[1]));
    wire [1:0] far_7_8075_1;    relay_conn far_7_8075_1_a(.in(far_7_8075_0[0]), .out(far_7_8075_1[0]));    relay_conn far_7_8075_1_b(.in(far_7_8075_0[1]), .out(far_7_8075_1[1]));
    assign out[935] = ~far_7_8075_1[1]; 
    wire [1:0] far_7_8076_0;    relay_conn far_7_8076_0_a(.in(layer_6[119]), .out(far_7_8076_0[0]));    relay_conn far_7_8076_0_b(.in(layer_6[190]), .out(far_7_8076_0[1]));
    wire [1:0] far_7_8076_1;    relay_conn far_7_8076_1_a(.in(far_7_8076_0[0]), .out(far_7_8076_1[0]));    relay_conn far_7_8076_1_b(.in(far_7_8076_0[1]), .out(far_7_8076_1[1]));
    assign out[936] = ~(far_7_8076_1[0] | far_7_8076_1[1]); 
    assign out[937] = ~layer_6[345]; 
    wire [1:0] far_7_8078_0;    relay_conn far_7_8078_0_a(.in(layer_6[605]), .out(far_7_8078_0[0]));    relay_conn far_7_8078_0_b(.in(layer_6[663]), .out(far_7_8078_0[1]));
    assign out[938] = ~(far_7_8078_0[0] | far_7_8078_0[1]); 
    assign out[939] = ~(layer_6[149] | layer_6[140]); 
    wire [1:0] far_7_8080_0;    relay_conn far_7_8080_0_a(.in(layer_6[26]), .out(far_7_8080_0[0]));    relay_conn far_7_8080_0_b(.in(layer_6[128]), .out(far_7_8080_0[1]));
    wire [1:0] far_7_8080_1;    relay_conn far_7_8080_1_a(.in(far_7_8080_0[0]), .out(far_7_8080_1[0]));    relay_conn far_7_8080_1_b(.in(far_7_8080_0[1]), .out(far_7_8080_1[1]));
    wire [1:0] far_7_8080_2;    relay_conn far_7_8080_2_a(.in(far_7_8080_1[0]), .out(far_7_8080_2[0]));    relay_conn far_7_8080_2_b(.in(far_7_8080_1[1]), .out(far_7_8080_2[1]));
    assign out[940] = far_7_8080_2[0] & far_7_8080_2[1]; 
    wire [1:0] far_7_8081_0;    relay_conn far_7_8081_0_a(.in(layer_6[920]), .out(far_7_8081_0[0]));    relay_conn far_7_8081_0_b(.in(layer_6[845]), .out(far_7_8081_0[1]));
    wire [1:0] far_7_8081_1;    relay_conn far_7_8081_1_a(.in(far_7_8081_0[0]), .out(far_7_8081_1[0]));    relay_conn far_7_8081_1_b(.in(far_7_8081_0[1]), .out(far_7_8081_1[1]));
    assign out[941] = far_7_8081_1[1]; 
    assign out[942] = layer_6[970] & layer_6[956]; 
    wire [1:0] far_7_8083_0;    relay_conn far_7_8083_0_a(.in(layer_6[966]), .out(far_7_8083_0[0]));    relay_conn far_7_8083_0_b(.in(layer_6[930]), .out(far_7_8083_0[1]));
    assign out[943] = far_7_8083_0[0] & far_7_8083_0[1]; 
    wire [1:0] far_7_8084_0;    relay_conn far_7_8084_0_a(.in(layer_6[412]), .out(far_7_8084_0[0]));    relay_conn far_7_8084_0_b(.in(layer_6[511]), .out(far_7_8084_0[1]));
    wire [1:0] far_7_8084_1;    relay_conn far_7_8084_1_a(.in(far_7_8084_0[0]), .out(far_7_8084_1[0]));    relay_conn far_7_8084_1_b(.in(far_7_8084_0[1]), .out(far_7_8084_1[1]));
    wire [1:0] far_7_8084_2;    relay_conn far_7_8084_2_a(.in(far_7_8084_1[0]), .out(far_7_8084_2[0]));    relay_conn far_7_8084_2_b(.in(far_7_8084_1[1]), .out(far_7_8084_2[1]));
    assign out[944] = far_7_8084_2[0] & far_7_8084_2[1]; 
    wire [1:0] far_7_8085_0;    relay_conn far_7_8085_0_a(.in(layer_6[659]), .out(far_7_8085_0[0]));    relay_conn far_7_8085_0_b(.in(layer_6[550]), .out(far_7_8085_0[1]));
    wire [1:0] far_7_8085_1;    relay_conn far_7_8085_1_a(.in(far_7_8085_0[0]), .out(far_7_8085_1[0]));    relay_conn far_7_8085_1_b(.in(far_7_8085_0[1]), .out(far_7_8085_1[1]));
    wire [1:0] far_7_8085_2;    relay_conn far_7_8085_2_a(.in(far_7_8085_1[0]), .out(far_7_8085_2[0]));    relay_conn far_7_8085_2_b(.in(far_7_8085_1[1]), .out(far_7_8085_2[1]));
    assign out[945] = ~(far_7_8085_2[0] | far_7_8085_2[1]); 
    wire [1:0] far_7_8086_0;    relay_conn far_7_8086_0_a(.in(layer_6[331]), .out(far_7_8086_0[0]));    relay_conn far_7_8086_0_b(.in(layer_6[216]), .out(far_7_8086_0[1]));
    wire [1:0] far_7_8086_1;    relay_conn far_7_8086_1_a(.in(far_7_8086_0[0]), .out(far_7_8086_1[0]));    relay_conn far_7_8086_1_b(.in(far_7_8086_0[1]), .out(far_7_8086_1[1]));
    wire [1:0] far_7_8086_2;    relay_conn far_7_8086_2_a(.in(far_7_8086_1[0]), .out(far_7_8086_2[0]));    relay_conn far_7_8086_2_b(.in(far_7_8086_1[1]), .out(far_7_8086_2[1]));
    assign out[946] = ~far_7_8086_2[1]; 
    wire [1:0] far_7_8087_0;    relay_conn far_7_8087_0_a(.in(layer_6[253]), .out(far_7_8087_0[0]));    relay_conn far_7_8087_0_b(.in(layer_6[204]), .out(far_7_8087_0[1]));
    assign out[947] = far_7_8087_0[0] & ~far_7_8087_0[1]; 
    wire [1:0] far_7_8088_0;    relay_conn far_7_8088_0_a(.in(layer_6[469]), .out(far_7_8088_0[0]));    relay_conn far_7_8088_0_b(.in(layer_6[435]), .out(far_7_8088_0[1]));
    assign out[948] = ~far_7_8088_0[0]; 
    wire [1:0] far_7_8089_0;    relay_conn far_7_8089_0_a(.in(layer_6[982]), .out(far_7_8089_0[0]));    relay_conn far_7_8089_0_b(.in(layer_6[859]), .out(far_7_8089_0[1]));
    wire [1:0] far_7_8089_1;    relay_conn far_7_8089_1_a(.in(far_7_8089_0[0]), .out(far_7_8089_1[0]));    relay_conn far_7_8089_1_b(.in(far_7_8089_0[1]), .out(far_7_8089_1[1]));
    wire [1:0] far_7_8089_2;    relay_conn far_7_8089_2_a(.in(far_7_8089_1[0]), .out(far_7_8089_2[0]));    relay_conn far_7_8089_2_b(.in(far_7_8089_1[1]), .out(far_7_8089_2[1]));
    assign out[949] = ~far_7_8089_2[1]; 
    wire [1:0] far_7_8090_0;    relay_conn far_7_8090_0_a(.in(layer_6[191]), .out(far_7_8090_0[0]));    relay_conn far_7_8090_0_b(.in(layer_6[128]), .out(far_7_8090_0[1]));
    assign out[950] = far_7_8090_0[0] & far_7_8090_0[1]; 
    assign out[951] = layer_6[422]; 
    wire [1:0] far_7_8092_0;    relay_conn far_7_8092_0_a(.in(layer_6[1019]), .out(far_7_8092_0[0]));    relay_conn far_7_8092_0_b(.in(layer_6[971]), .out(far_7_8092_0[1]));
    assign out[952] = far_7_8092_0[0] & ~far_7_8092_0[1]; 
    wire [1:0] far_7_8093_0;    relay_conn far_7_8093_0_a(.in(layer_6[109]), .out(far_7_8093_0[0]));    relay_conn far_7_8093_0_b(.in(layer_6[170]), .out(far_7_8093_0[1]));
    assign out[953] = far_7_8093_0[0]; 
    wire [1:0] far_7_8094_0;    relay_conn far_7_8094_0_a(.in(layer_6[706]), .out(far_7_8094_0[0]));    relay_conn far_7_8094_0_b(.in(layer_6[601]), .out(far_7_8094_0[1]));
    wire [1:0] far_7_8094_1;    relay_conn far_7_8094_1_a(.in(far_7_8094_0[0]), .out(far_7_8094_1[0]));    relay_conn far_7_8094_1_b(.in(far_7_8094_0[1]), .out(far_7_8094_1[1]));
    wire [1:0] far_7_8094_2;    relay_conn far_7_8094_2_a(.in(far_7_8094_1[0]), .out(far_7_8094_2[0]));    relay_conn far_7_8094_2_b(.in(far_7_8094_1[1]), .out(far_7_8094_2[1]));
    assign out[954] = far_7_8094_2[0] & far_7_8094_2[1]; 
    wire [1:0] far_7_8095_0;    relay_conn far_7_8095_0_a(.in(layer_6[321]), .out(far_7_8095_0[0]));    relay_conn far_7_8095_0_b(.in(layer_6[449]), .out(far_7_8095_0[1]));
    wire [1:0] far_7_8095_1;    relay_conn far_7_8095_1_a(.in(far_7_8095_0[0]), .out(far_7_8095_1[0]));    relay_conn far_7_8095_1_b(.in(far_7_8095_0[1]), .out(far_7_8095_1[1]));
    wire [1:0] far_7_8095_2;    relay_conn far_7_8095_2_a(.in(far_7_8095_1[0]), .out(far_7_8095_2[0]));    relay_conn far_7_8095_2_b(.in(far_7_8095_1[1]), .out(far_7_8095_2[1]));
    wire [1:0] far_7_8095_3;    relay_conn far_7_8095_3_a(.in(far_7_8095_2[0]), .out(far_7_8095_3[0]));    relay_conn far_7_8095_3_b(.in(far_7_8095_2[1]), .out(far_7_8095_3[1]));
    assign out[955] = ~(far_7_8095_3[0] | far_7_8095_3[1]); 
    wire [1:0] far_7_8096_0;    relay_conn far_7_8096_0_a(.in(layer_6[565]), .out(far_7_8096_0[0]));    relay_conn far_7_8096_0_b(.in(layer_6[442]), .out(far_7_8096_0[1]));
    wire [1:0] far_7_8096_1;    relay_conn far_7_8096_1_a(.in(far_7_8096_0[0]), .out(far_7_8096_1[0]));    relay_conn far_7_8096_1_b(.in(far_7_8096_0[1]), .out(far_7_8096_1[1]));
    wire [1:0] far_7_8096_2;    relay_conn far_7_8096_2_a(.in(far_7_8096_1[0]), .out(far_7_8096_2[0]));    relay_conn far_7_8096_2_b(.in(far_7_8096_1[1]), .out(far_7_8096_2[1]));
    assign out[956] = far_7_8096_2[1] & ~far_7_8096_2[0]; 
    wire [1:0] far_7_8097_0;    relay_conn far_7_8097_0_a(.in(layer_6[730]), .out(far_7_8097_0[0]));    relay_conn far_7_8097_0_b(.in(layer_6[803]), .out(far_7_8097_0[1]));
    wire [1:0] far_7_8097_1;    relay_conn far_7_8097_1_a(.in(far_7_8097_0[0]), .out(far_7_8097_1[0]));    relay_conn far_7_8097_1_b(.in(far_7_8097_0[1]), .out(far_7_8097_1[1]));
    assign out[957] = far_7_8097_1[0]; 
    wire [1:0] far_7_8098_0;    relay_conn far_7_8098_0_a(.in(layer_6[284]), .out(far_7_8098_0[0]));    relay_conn far_7_8098_0_b(.in(layer_6[350]), .out(far_7_8098_0[1]));
    wire [1:0] far_7_8098_1;    relay_conn far_7_8098_1_a(.in(far_7_8098_0[0]), .out(far_7_8098_1[0]));    relay_conn far_7_8098_1_b(.in(far_7_8098_0[1]), .out(far_7_8098_1[1]));
    assign out[958] = far_7_8098_1[1] & ~far_7_8098_1[0]; 
    wire [1:0] far_7_8099_0;    relay_conn far_7_8099_0_a(.in(layer_6[415]), .out(far_7_8099_0[0]));    relay_conn far_7_8099_0_b(.in(layer_6[334]), .out(far_7_8099_0[1]));
    wire [1:0] far_7_8099_1;    relay_conn far_7_8099_1_a(.in(far_7_8099_0[0]), .out(far_7_8099_1[0]));    relay_conn far_7_8099_1_b(.in(far_7_8099_0[1]), .out(far_7_8099_1[1]));
    assign out[959] = ~(far_7_8099_1[0] | far_7_8099_1[1]); 
    assign out[960] = ~(layer_6[468] | layer_6[449]); 
    wire [1:0] far_7_8101_0;    relay_conn far_7_8101_0_a(.in(layer_6[733]), .out(far_7_8101_0[0]));    relay_conn far_7_8101_0_b(.in(layer_6[811]), .out(far_7_8101_0[1]));
    wire [1:0] far_7_8101_1;    relay_conn far_7_8101_1_a(.in(far_7_8101_0[0]), .out(far_7_8101_1[0]));    relay_conn far_7_8101_1_b(.in(far_7_8101_0[1]), .out(far_7_8101_1[1]));
    assign out[961] = far_7_8101_1[0]; 
    wire [1:0] far_7_8102_0;    relay_conn far_7_8102_0_a(.in(layer_6[794]), .out(far_7_8102_0[0]));    relay_conn far_7_8102_0_b(.in(layer_6[889]), .out(far_7_8102_0[1]));
    wire [1:0] far_7_8102_1;    relay_conn far_7_8102_1_a(.in(far_7_8102_0[0]), .out(far_7_8102_1[0]));    relay_conn far_7_8102_1_b(.in(far_7_8102_0[1]), .out(far_7_8102_1[1]));
    assign out[962] = ~(far_7_8102_1[0] ^ far_7_8102_1[1]); 
    assign out[963] = layer_6[72] & ~layer_6[56]; 
    wire [1:0] far_7_8104_0;    relay_conn far_7_8104_0_a(.in(layer_6[821]), .out(far_7_8104_0[0]));    relay_conn far_7_8104_0_b(.in(layer_6[789]), .out(far_7_8104_0[1]));
    assign out[964] = far_7_8104_0[0] & far_7_8104_0[1]; 
    assign out[965] = ~(layer_6[92] | layer_6[94]); 
    wire [1:0] far_7_8106_0;    relay_conn far_7_8106_0_a(.in(layer_6[845]), .out(far_7_8106_0[0]));    relay_conn far_7_8106_0_b(.in(layer_6[766]), .out(far_7_8106_0[1]));
    wire [1:0] far_7_8106_1;    relay_conn far_7_8106_1_a(.in(far_7_8106_0[0]), .out(far_7_8106_1[0]));    relay_conn far_7_8106_1_b(.in(far_7_8106_0[1]), .out(far_7_8106_1[1]));
    assign out[966] = far_7_8106_1[0]; 
    wire [1:0] far_7_8107_0;    relay_conn far_7_8107_0_a(.in(layer_6[925]), .out(far_7_8107_0[0]));    relay_conn far_7_8107_0_b(.in(layer_6[984]), .out(far_7_8107_0[1]));
    assign out[967] = far_7_8107_0[0]; 
    wire [1:0] far_7_8108_0;    relay_conn far_7_8108_0_a(.in(layer_6[54]), .out(far_7_8108_0[0]));    relay_conn far_7_8108_0_b(.in(layer_6[129]), .out(far_7_8108_0[1]));
    wire [1:0] far_7_8108_1;    relay_conn far_7_8108_1_a(.in(far_7_8108_0[0]), .out(far_7_8108_1[0]));    relay_conn far_7_8108_1_b(.in(far_7_8108_0[1]), .out(far_7_8108_1[1]));
    assign out[968] = ~(far_7_8108_1[0] & far_7_8108_1[1]); 
    wire [1:0] far_7_8109_0;    relay_conn far_7_8109_0_a(.in(layer_6[226]), .out(far_7_8109_0[0]));    relay_conn far_7_8109_0_b(.in(layer_6[305]), .out(far_7_8109_0[1]));
    wire [1:0] far_7_8109_1;    relay_conn far_7_8109_1_a(.in(far_7_8109_0[0]), .out(far_7_8109_1[0]));    relay_conn far_7_8109_1_b(.in(far_7_8109_0[1]), .out(far_7_8109_1[1]));
    assign out[969] = ~(far_7_8109_1[0] | far_7_8109_1[1]); 
    wire [1:0] far_7_8110_0;    relay_conn far_7_8110_0_a(.in(layer_6[194]), .out(far_7_8110_0[0]));    relay_conn far_7_8110_0_b(.in(layer_6[257]), .out(far_7_8110_0[1]));
    assign out[970] = far_7_8110_0[1] & ~far_7_8110_0[0]; 
    wire [1:0] far_7_8111_0;    relay_conn far_7_8111_0_a(.in(layer_6[908]), .out(far_7_8111_0[0]));    relay_conn far_7_8111_0_b(.in(layer_6[822]), .out(far_7_8111_0[1]));
    wire [1:0] far_7_8111_1;    relay_conn far_7_8111_1_a(.in(far_7_8111_0[0]), .out(far_7_8111_1[0]));    relay_conn far_7_8111_1_b(.in(far_7_8111_0[1]), .out(far_7_8111_1[1]));
    assign out[971] = far_7_8111_1[1]; 
    wire [1:0] far_7_8112_0;    relay_conn far_7_8112_0_a(.in(layer_6[524]), .out(far_7_8112_0[0]));    relay_conn far_7_8112_0_b(.in(layer_6[456]), .out(far_7_8112_0[1]));
    wire [1:0] far_7_8112_1;    relay_conn far_7_8112_1_a(.in(far_7_8112_0[0]), .out(far_7_8112_1[0]));    relay_conn far_7_8112_1_b(.in(far_7_8112_0[1]), .out(far_7_8112_1[1]));
    assign out[972] = ~far_7_8112_1[0]; 
    wire [1:0] far_7_8113_0;    relay_conn far_7_8113_0_a(.in(layer_6[897]), .out(far_7_8113_0[0]));    relay_conn far_7_8113_0_b(.in(layer_6[802]), .out(far_7_8113_0[1]));
    wire [1:0] far_7_8113_1;    relay_conn far_7_8113_1_a(.in(far_7_8113_0[0]), .out(far_7_8113_1[0]));    relay_conn far_7_8113_1_b(.in(far_7_8113_0[1]), .out(far_7_8113_1[1]));
    assign out[973] = far_7_8113_1[0] & ~far_7_8113_1[1]; 
    wire [1:0] far_7_8114_0;    relay_conn far_7_8114_0_a(.in(layer_6[570]), .out(far_7_8114_0[0]));    relay_conn far_7_8114_0_b(.in(layer_6[650]), .out(far_7_8114_0[1]));
    wire [1:0] far_7_8114_1;    relay_conn far_7_8114_1_a(.in(far_7_8114_0[0]), .out(far_7_8114_1[0]));    relay_conn far_7_8114_1_b(.in(far_7_8114_0[1]), .out(far_7_8114_1[1]));
    assign out[974] = far_7_8114_1[1]; 
    wire [1:0] far_7_8115_0;    relay_conn far_7_8115_0_a(.in(layer_6[854]), .out(far_7_8115_0[0]));    relay_conn far_7_8115_0_b(.in(layer_6[972]), .out(far_7_8115_0[1]));
    wire [1:0] far_7_8115_1;    relay_conn far_7_8115_1_a(.in(far_7_8115_0[0]), .out(far_7_8115_1[0]));    relay_conn far_7_8115_1_b(.in(far_7_8115_0[1]), .out(far_7_8115_1[1]));
    wire [1:0] far_7_8115_2;    relay_conn far_7_8115_2_a(.in(far_7_8115_1[0]), .out(far_7_8115_2[0]));    relay_conn far_7_8115_2_b(.in(far_7_8115_1[1]), .out(far_7_8115_2[1]));
    assign out[975] = ~(far_7_8115_2[0] ^ far_7_8115_2[1]); 
    wire [1:0] far_7_8116_0;    relay_conn far_7_8116_0_a(.in(layer_6[652]), .out(far_7_8116_0[0]));    relay_conn far_7_8116_0_b(.in(layer_6[575]), .out(far_7_8116_0[1]));
    wire [1:0] far_7_8116_1;    relay_conn far_7_8116_1_a(.in(far_7_8116_0[0]), .out(far_7_8116_1[0]));    relay_conn far_7_8116_1_b(.in(far_7_8116_0[1]), .out(far_7_8116_1[1]));
    assign out[976] = far_7_8116_1[1] & ~far_7_8116_1[0]; 
    assign out[977] = ~layer_6[416]; 
    wire [1:0] far_7_8118_0;    relay_conn far_7_8118_0_a(.in(layer_6[229]), .out(far_7_8118_0[0]));    relay_conn far_7_8118_0_b(.in(layer_6[119]), .out(far_7_8118_0[1]));
    wire [1:0] far_7_8118_1;    relay_conn far_7_8118_1_a(.in(far_7_8118_0[0]), .out(far_7_8118_1[0]));    relay_conn far_7_8118_1_b(.in(far_7_8118_0[1]), .out(far_7_8118_1[1]));
    wire [1:0] far_7_8118_2;    relay_conn far_7_8118_2_a(.in(far_7_8118_1[0]), .out(far_7_8118_2[0]));    relay_conn far_7_8118_2_b(.in(far_7_8118_1[1]), .out(far_7_8118_2[1]));
    assign out[978] = far_7_8118_2[0] & ~far_7_8118_2[1]; 
    assign out[979] = layer_6[685]; 
    assign out[980] = layer_6[289] & ~layer_6[293]; 
    assign out[981] = ~layer_6[923]; 
    wire [1:0] far_7_8122_0;    relay_conn far_7_8122_0_a(.in(layer_6[293]), .out(far_7_8122_0[0]));    relay_conn far_7_8122_0_b(.in(layer_6[197]), .out(far_7_8122_0[1]));
    wire [1:0] far_7_8122_1;    relay_conn far_7_8122_1_a(.in(far_7_8122_0[0]), .out(far_7_8122_1[0]));    relay_conn far_7_8122_1_b(.in(far_7_8122_0[1]), .out(far_7_8122_1[1]));
    wire [1:0] far_7_8122_2;    relay_conn far_7_8122_2_a(.in(far_7_8122_1[0]), .out(far_7_8122_2[0]));    relay_conn far_7_8122_2_b(.in(far_7_8122_1[1]), .out(far_7_8122_2[1]));
    assign out[982] = ~far_7_8122_2[0] | (far_7_8122_2[0] & far_7_8122_2[1]); 
    assign out[983] = ~layer_6[416]; 
    wire [1:0] far_7_8124_0;    relay_conn far_7_8124_0_a(.in(layer_6[739]), .out(far_7_8124_0[0]));    relay_conn far_7_8124_0_b(.in(layer_6[781]), .out(far_7_8124_0[1]));
    assign out[984] = far_7_8124_0[0] & ~far_7_8124_0[1]; 
    wire [1:0] far_7_8125_0;    relay_conn far_7_8125_0_a(.in(layer_6[404]), .out(far_7_8125_0[0]));    relay_conn far_7_8125_0_b(.in(layer_6[472]), .out(far_7_8125_0[1]));
    wire [1:0] far_7_8125_1;    relay_conn far_7_8125_1_a(.in(far_7_8125_0[0]), .out(far_7_8125_1[0]));    relay_conn far_7_8125_1_b(.in(far_7_8125_0[1]), .out(far_7_8125_1[1]));
    assign out[985] = ~far_7_8125_1[1]; 
    wire [1:0] far_7_8126_0;    relay_conn far_7_8126_0_a(.in(layer_6[211]), .out(far_7_8126_0[0]));    relay_conn far_7_8126_0_b(.in(layer_6[130]), .out(far_7_8126_0[1]));
    wire [1:0] far_7_8126_1;    relay_conn far_7_8126_1_a(.in(far_7_8126_0[0]), .out(far_7_8126_1[0]));    relay_conn far_7_8126_1_b(.in(far_7_8126_0[1]), .out(far_7_8126_1[1]));
    assign out[986] = far_7_8126_1[0] ^ far_7_8126_1[1]; 
    wire [1:0] far_7_8127_0;    relay_conn far_7_8127_0_a(.in(layer_6[150]), .out(far_7_8127_0[0]));    relay_conn far_7_8127_0_b(.in(layer_6[47]), .out(far_7_8127_0[1]));
    wire [1:0] far_7_8127_1;    relay_conn far_7_8127_1_a(.in(far_7_8127_0[0]), .out(far_7_8127_1[0]));    relay_conn far_7_8127_1_b(.in(far_7_8127_0[1]), .out(far_7_8127_1[1]));
    wire [1:0] far_7_8127_2;    relay_conn far_7_8127_2_a(.in(far_7_8127_1[0]), .out(far_7_8127_2[0]));    relay_conn far_7_8127_2_b(.in(far_7_8127_1[1]), .out(far_7_8127_2[1]));
    assign out[987] = far_7_8127_2[1] & ~far_7_8127_2[0]; 
    assign out[988] = ~(layer_6[150] | layer_6[119]); 
    wire [1:0] far_7_8129_0;    relay_conn far_7_8129_0_a(.in(layer_6[324]), .out(far_7_8129_0[0]));    relay_conn far_7_8129_0_b(.in(layer_6[397]), .out(far_7_8129_0[1]));
    wire [1:0] far_7_8129_1;    relay_conn far_7_8129_1_a(.in(far_7_8129_0[0]), .out(far_7_8129_1[0]));    relay_conn far_7_8129_1_b(.in(far_7_8129_0[1]), .out(far_7_8129_1[1]));
    assign out[989] = ~far_7_8129_1[0]; 
    wire [1:0] far_7_8130_0;    relay_conn far_7_8130_0_a(.in(layer_6[153]), .out(far_7_8130_0[0]));    relay_conn far_7_8130_0_b(.in(layer_6[56]), .out(far_7_8130_0[1]));
    wire [1:0] far_7_8130_1;    relay_conn far_7_8130_1_a(.in(far_7_8130_0[0]), .out(far_7_8130_1[0]));    relay_conn far_7_8130_1_b(.in(far_7_8130_0[1]), .out(far_7_8130_1[1]));
    wire [1:0] far_7_8130_2;    relay_conn far_7_8130_2_a(.in(far_7_8130_1[0]), .out(far_7_8130_2[0]));    relay_conn far_7_8130_2_b(.in(far_7_8130_1[1]), .out(far_7_8130_2[1]));
    assign out[990] = far_7_8130_2[0] & ~far_7_8130_2[1]; 
    wire [1:0] far_7_8131_0;    relay_conn far_7_8131_0_a(.in(layer_6[778]), .out(far_7_8131_0[0]));    relay_conn far_7_8131_0_b(.in(layer_6[896]), .out(far_7_8131_0[1]));
    wire [1:0] far_7_8131_1;    relay_conn far_7_8131_1_a(.in(far_7_8131_0[0]), .out(far_7_8131_1[0]));    relay_conn far_7_8131_1_b(.in(far_7_8131_0[1]), .out(far_7_8131_1[1]));
    wire [1:0] far_7_8131_2;    relay_conn far_7_8131_2_a(.in(far_7_8131_1[0]), .out(far_7_8131_2[0]));    relay_conn far_7_8131_2_b(.in(far_7_8131_1[1]), .out(far_7_8131_2[1]));
    assign out[991] = far_7_8131_2[0]; 
    wire [1:0] far_7_8132_0;    relay_conn far_7_8132_0_a(.in(layer_6[1009]), .out(far_7_8132_0[0]));    relay_conn far_7_8132_0_b(.in(layer_6[916]), .out(far_7_8132_0[1]));
    wire [1:0] far_7_8132_1;    relay_conn far_7_8132_1_a(.in(far_7_8132_0[0]), .out(far_7_8132_1[0]));    relay_conn far_7_8132_1_b(.in(far_7_8132_0[1]), .out(far_7_8132_1[1]));
    assign out[992] = far_7_8132_1[0] ^ far_7_8132_1[1]; 
    wire [1:0] far_7_8133_0;    relay_conn far_7_8133_0_a(.in(layer_6[141]), .out(far_7_8133_0[0]));    relay_conn far_7_8133_0_b(.in(layer_6[267]), .out(far_7_8133_0[1]));
    wire [1:0] far_7_8133_1;    relay_conn far_7_8133_1_a(.in(far_7_8133_0[0]), .out(far_7_8133_1[0]));    relay_conn far_7_8133_1_b(.in(far_7_8133_0[1]), .out(far_7_8133_1[1]));
    wire [1:0] far_7_8133_2;    relay_conn far_7_8133_2_a(.in(far_7_8133_1[0]), .out(far_7_8133_2[0]));    relay_conn far_7_8133_2_b(.in(far_7_8133_1[1]), .out(far_7_8133_2[1]));
    assign out[993] = far_7_8133_2[1] & ~far_7_8133_2[0]; 
    wire [1:0] far_7_8134_0;    relay_conn far_7_8134_0_a(.in(layer_6[666]), .out(far_7_8134_0[0]));    relay_conn far_7_8134_0_b(.in(layer_6[711]), .out(far_7_8134_0[1]));
    assign out[994] = ~(far_7_8134_0[0] | far_7_8134_0[1]); 
    wire [1:0] far_7_8135_0;    relay_conn far_7_8135_0_a(.in(layer_6[848]), .out(far_7_8135_0[0]));    relay_conn far_7_8135_0_b(.in(layer_6[783]), .out(far_7_8135_0[1]));
    wire [1:0] far_7_8135_1;    relay_conn far_7_8135_1_a(.in(far_7_8135_0[0]), .out(far_7_8135_1[0]));    relay_conn far_7_8135_1_b(.in(far_7_8135_0[1]), .out(far_7_8135_1[1]));
    assign out[995] = far_7_8135_1[0] ^ far_7_8135_1[1]; 
    wire [1:0] far_7_8136_0;    relay_conn far_7_8136_0_a(.in(layer_6[511]), .out(far_7_8136_0[0]));    relay_conn far_7_8136_0_b(.in(layer_6[392]), .out(far_7_8136_0[1]));
    wire [1:0] far_7_8136_1;    relay_conn far_7_8136_1_a(.in(far_7_8136_0[0]), .out(far_7_8136_1[0]));    relay_conn far_7_8136_1_b(.in(far_7_8136_0[1]), .out(far_7_8136_1[1]));
    wire [1:0] far_7_8136_2;    relay_conn far_7_8136_2_a(.in(far_7_8136_1[0]), .out(far_7_8136_2[0]));    relay_conn far_7_8136_2_b(.in(far_7_8136_1[1]), .out(far_7_8136_2[1]));
    assign out[996] = far_7_8136_2[0]; 
    wire [1:0] far_7_8137_0;    relay_conn far_7_8137_0_a(.in(layer_6[623]), .out(far_7_8137_0[0]));    relay_conn far_7_8137_0_b(.in(layer_6[685]), .out(far_7_8137_0[1]));
    assign out[997] = far_7_8137_0[1]; 
    wire [1:0] far_7_8138_0;    relay_conn far_7_8138_0_a(.in(layer_6[478]), .out(far_7_8138_0[0]));    relay_conn far_7_8138_0_b(.in(layer_6[392]), .out(far_7_8138_0[1]));
    wire [1:0] far_7_8138_1;    relay_conn far_7_8138_1_a(.in(far_7_8138_0[0]), .out(far_7_8138_1[0]));    relay_conn far_7_8138_1_b(.in(far_7_8138_0[1]), .out(far_7_8138_1[1]));
    assign out[998] = ~far_7_8138_1[0]; 
    wire [1:0] far_7_8139_0;    relay_conn far_7_8139_0_a(.in(layer_6[908]), .out(far_7_8139_0[0]));    relay_conn far_7_8139_0_b(.in(layer_6[845]), .out(far_7_8139_0[1]));
    assign out[999] = far_7_8139_0[1]; 
    wire [1:0] far_7_8140_0;    relay_conn far_7_8140_0_a(.in(layer_6[611]), .out(far_7_8140_0[0]));    relay_conn far_7_8140_0_b(.in(layer_6[648]), .out(far_7_8140_0[1]));
    assign out[1000] = far_7_8140_0[0] & ~far_7_8140_0[1]; 
    wire [1:0] far_7_8141_0;    relay_conn far_7_8141_0_a(.in(layer_6[392]), .out(far_7_8141_0[0]));    relay_conn far_7_8141_0_b(.in(layer_6[504]), .out(far_7_8141_0[1]));
    wire [1:0] far_7_8141_1;    relay_conn far_7_8141_1_a(.in(far_7_8141_0[0]), .out(far_7_8141_1[0]));    relay_conn far_7_8141_1_b(.in(far_7_8141_0[1]), .out(far_7_8141_1[1]));
    wire [1:0] far_7_8141_2;    relay_conn far_7_8141_2_a(.in(far_7_8141_1[0]), .out(far_7_8141_2[0]));    relay_conn far_7_8141_2_b(.in(far_7_8141_1[1]), .out(far_7_8141_2[1]));
    assign out[1001] = far_7_8141_2[1]; 
    assign out[1002] = layer_6[492] & ~layer_6[474]; 
    wire [1:0] far_7_8143_0;    relay_conn far_7_8143_0_a(.in(layer_6[718]), .out(far_7_8143_0[0]));    relay_conn far_7_8143_0_b(.in(layer_6[682]), .out(far_7_8143_0[1]));
    assign out[1003] = ~far_7_8143_0[1]; 
    assign out[1004] = layer_6[651] & ~layer_6[645]; 
    wire [1:0] far_7_8145_0;    relay_conn far_7_8145_0_a(.in(layer_6[740]), .out(far_7_8145_0[0]));    relay_conn far_7_8145_0_b(.in(layer_6[802]), .out(far_7_8145_0[1]));
    assign out[1005] = ~(far_7_8145_0[0] | far_7_8145_0[1]); 
    assign out[1006] = ~layer_6[324]; 
    wire [1:0] far_7_8147_0;    relay_conn far_7_8147_0_a(.in(layer_6[178]), .out(far_7_8147_0[0]));    relay_conn far_7_8147_0_b(.in(layer_6[141]), .out(far_7_8147_0[1]));
    assign out[1007] = ~(far_7_8147_0[0] | far_7_8147_0[1]); 
    wire [1:0] far_7_8148_0;    relay_conn far_7_8148_0_a(.in(layer_6[625]), .out(far_7_8148_0[0]));    relay_conn far_7_8148_0_b(.in(layer_6[497]), .out(far_7_8148_0[1]));
    wire [1:0] far_7_8148_1;    relay_conn far_7_8148_1_a(.in(far_7_8148_0[0]), .out(far_7_8148_1[0]));    relay_conn far_7_8148_1_b(.in(far_7_8148_0[1]), .out(far_7_8148_1[1]));
    wire [1:0] far_7_8148_2;    relay_conn far_7_8148_2_a(.in(far_7_8148_1[0]), .out(far_7_8148_2[0]));    relay_conn far_7_8148_2_b(.in(far_7_8148_1[1]), .out(far_7_8148_2[1]));
    wire [1:0] far_7_8148_3;    relay_conn far_7_8148_3_a(.in(far_7_8148_2[0]), .out(far_7_8148_3[0]));    relay_conn far_7_8148_3_b(.in(far_7_8148_2[1]), .out(far_7_8148_3[1]));
    assign out[1008] = far_7_8148_3[1] & ~far_7_8148_3[0]; 
    assign out[1009] = layer_6[431] & ~layer_6[449]; 
    assign out[1010] = layer_6[624] & ~layer_6[635]; 
    wire [1:0] far_7_8151_0;    relay_conn far_7_8151_0_a(.in(layer_6[403]), .out(far_7_8151_0[0]));    relay_conn far_7_8151_0_b(.in(layer_6[364]), .out(far_7_8151_0[1]));
    assign out[1011] = ~far_7_8151_0[1] | (far_7_8151_0[0] & far_7_8151_0[1]); 
    assign out[1012] = layer_6[458] & ~layer_6[480]; 
    wire [1:0] far_7_8153_0;    relay_conn far_7_8153_0_a(.in(layer_6[692]), .out(far_7_8153_0[0]));    relay_conn far_7_8153_0_b(.in(layer_6[812]), .out(far_7_8153_0[1]));
    wire [1:0] far_7_8153_1;    relay_conn far_7_8153_1_a(.in(far_7_8153_0[0]), .out(far_7_8153_1[0]));    relay_conn far_7_8153_1_b(.in(far_7_8153_0[1]), .out(far_7_8153_1[1]));
    wire [1:0] far_7_8153_2;    relay_conn far_7_8153_2_a(.in(far_7_8153_1[0]), .out(far_7_8153_2[0]));    relay_conn far_7_8153_2_b(.in(far_7_8153_1[1]), .out(far_7_8153_2[1]));
    assign out[1013] = far_7_8153_2[0]; 
    assign out[1014] = layer_6[71] & ~layer_6[97]; 
    wire [1:0] far_7_8155_0;    relay_conn far_7_8155_0_a(.in(layer_6[636]), .out(far_7_8155_0[0]));    relay_conn far_7_8155_0_b(.in(layer_6[511]), .out(far_7_8155_0[1]));
    wire [1:0] far_7_8155_1;    relay_conn far_7_8155_1_a(.in(far_7_8155_0[0]), .out(far_7_8155_1[0]));    relay_conn far_7_8155_1_b(.in(far_7_8155_0[1]), .out(far_7_8155_1[1]));
    wire [1:0] far_7_8155_2;    relay_conn far_7_8155_2_a(.in(far_7_8155_1[0]), .out(far_7_8155_2[0]));    relay_conn far_7_8155_2_b(.in(far_7_8155_1[1]), .out(far_7_8155_2[1]));
    assign out[1015] = far_7_8155_2[1]; 
    wire [1:0] far_7_8156_0;    relay_conn far_7_8156_0_a(.in(layer_6[60]), .out(far_7_8156_0[0]));    relay_conn far_7_8156_0_b(.in(layer_6[163]), .out(far_7_8156_0[1]));
    wire [1:0] far_7_8156_1;    relay_conn far_7_8156_1_a(.in(far_7_8156_0[0]), .out(far_7_8156_1[0]));    relay_conn far_7_8156_1_b(.in(far_7_8156_0[1]), .out(far_7_8156_1[1]));
    wire [1:0] far_7_8156_2;    relay_conn far_7_8156_2_a(.in(far_7_8156_1[0]), .out(far_7_8156_2[0]));    relay_conn far_7_8156_2_b(.in(far_7_8156_1[1]), .out(far_7_8156_2[1]));
    assign out[1016] = far_7_8156_2[0] & far_7_8156_2[1]; 
    wire [1:0] far_7_8157_0;    relay_conn far_7_8157_0_a(.in(layer_6[720]), .out(far_7_8157_0[0]));    relay_conn far_7_8157_0_b(.in(layer_6[670]), .out(far_7_8157_0[1]));
    assign out[1017] = far_7_8157_0[0] & ~far_7_8157_0[1]; 
    wire [1:0] far_7_8158_0;    relay_conn far_7_8158_0_a(.in(layer_6[71]), .out(far_7_8158_0[0]));    relay_conn far_7_8158_0_b(.in(layer_6[31]), .out(far_7_8158_0[1]));
    assign out[1018] = far_7_8158_0[0] & far_7_8158_0[1]; 
    assign out[1019] = ~layer_6[416]; 

endmodule
