// Generated from: binarized_20250122-110005_acc9041_seed876599_epochs300_3x1300_b256_lrm10-1with_dataset.npz

module net (
    input  wire [254:0] in,
    output wire [1299:0] out,
    output wire [2549:0] categories
);
    wire [1300:0] layer_0;
    wire [1300:0] layer_1;

    // Layer 0 ============================================================
    assign layer_0[0] = in[75] | in[92]; 
    assign layer_0[1] = in[89] | in[214]; 
    assign layer_0[2] = in[131] | in[133]; 
    assign layer_0[3] = in[252] | in[101]; 
    assign layer_0[4] = in[100] | in[92]; 
    assign layer_0[5] = in[246] | in[116]; 
    assign layer_0[6] = in[139] | in[163]; 
    assign layer_0[7] = in[124] | in[117]; 
    assign layer_0[8] = in[90]; 
    assign layer_0[9] = in[116] | in[229]; 
    assign layer_0[10] = ~in[40]; 
    assign layer_0[11] = in[85] & ~in[188]; 
    assign layer_0[12] = in[115] | in[101]; 
    assign layer_0[13] = in[116] | in[75]; 
    assign layer_0[14] = in[101] | in[108]; 
    assign layer_0[15] = in[75]; 
    assign layer_0[16] = in[146] | in[116]; 
    assign layer_0[17] = in[27] | in[101]; 
    assign layer_0[18] = in[116] | in[117]; 
    assign layer_0[19] = in[108] | in[116]; 
    assign layer_0[20] = in[108] | in[248]; 
    assign layer_0[21] = in[92] | in[74]; 
    assign layer_0[22] = in[77] | in[90]; 
    assign layer_0[23] = in[132]; 
    assign layer_0[24] = in[91]; 
    assign layer_0[25] = in[132]; 
    assign layer_0[26] = in[132] | in[124]; 
    assign layer_0[27] = in[230] | in[100]; 
    assign layer_0[28] = ~in[40]; 
    assign layer_0[29] = in[101] | in[115]; 
    assign layer_0[30] = in[232] | in[75]; 
    assign layer_0[31] = in[246] | in[74]; 
    assign layer_0[32] = in[100] | in[246]; 
    assign layer_0[33] = in[235] | in[86]; 
    assign layer_0[34] = in[90] | in[92]; 
    assign layer_0[35] = ~in[151]; 
    assign layer_0[36] = in[101]; 
    assign layer_0[37] = in[101] | in[116]; 
    assign layer_0[38] = ~in[182]; 
    assign layer_0[39] = in[107] | in[115]; 
    assign layer_0[40] = in[92] | in[90]; 
    assign layer_0[41] = in[117] | in[115]; 
    assign layer_0[42] = in[235] | in[91]; 
    assign layer_0[43] = in[52] | in[91]; 
    assign layer_0[44] = in[91] | in[92]; 
    assign layer_0[45] = in[232] | in[230]; 
    assign layer_0[46] = in[132]; 
    assign layer_0[47] = in[117] ^ in[172]; 
    assign layer_0[48] = in[118] & ~in[22]; 
    assign layer_0[49] = in[115] | in[90]; 
    assign layer_0[50] = in[117] | in[100]; 
    assign layer_0[51] = in[90] | in[171]; 
    assign layer_0[52] = in[72] & ~in[61]; 
    assign layer_0[53] = in[131] | in[117]; 
    assign layer_0[54] = ~(in[121] | in[231]); 
    assign layer_0[55] = in[247] ^ in[233]; 
    assign layer_0[56] = in[115] | in[132]; 
    assign layer_0[57] = in[232] | in[90]; 
    assign layer_0[58] = in[132] | in[108]; 
    assign layer_0[59] = ~in[151]; 
    assign layer_0[60] = in[108] | in[116]; 
    assign layer_0[61] = in[100] | in[247]; 
    assign layer_0[62] = in[101] | in[83]; 
    assign layer_0[63] = in[231] | in[233]; 
    assign layer_0[64] = ~in[150]; 
    assign layer_0[65] = in[102] | in[117]; 
    assign layer_0[66] = in[115] | in[117]; 
    assign layer_0[67] = ~in[40]; 
    assign layer_0[68] = in[74]; 
    assign layer_0[69] = in[85] | in[194]; 
    assign layer_0[70] = in[117] | in[116]; 
    assign layer_0[71] = ~in[40]; 
    assign layer_0[72] = in[234] | in[91]; 
    assign layer_0[73] = in[216] | in[229]; 
    assign layer_0[74] = in[101] | in[182]; 
    assign layer_0[75] = in[84] | in[91]; 
    assign layer_0[76] = in[92] | in[232]; 
    assign layer_0[77] = in[76] | in[85]; 
    assign layer_0[78] = in[100] | in[247]; 
    assign layer_0[79] = in[91] | in[116]; 
    assign layer_0[80] = in[248] | in[116]; 
    assign layer_0[81] = in[248] | in[101]; 
    assign layer_0[82] = in[138] & ~in[197]; 
    assign layer_0[83] = in[132] | in[246]; 
    assign layer_0[84] = in[101]; 
    assign layer_0[85] = in[132] | in[132]; 
    assign layer_0[86] = in[91]; 
    assign layer_0[87] = in[108] | in[234]; 
    assign layer_0[88] = in[101]; 
    assign layer_0[89] = in[101] | in[116]; 
    assign layer_0[90] = in[155] ^ in[102]; 
    assign layer_0[91] = in[90]; 
    assign layer_0[92] = in[83] | in[116]; 
    assign layer_0[93] = in[116] | in[108]; 
    assign layer_0[94] = in[90]; 
    assign layer_0[95] = in[59] | in[90]; 
    assign layer_0[96] = ~in[41] | (in[41] & in[99]); 
    assign layer_0[97] = in[117]; 
    assign layer_0[98] = ~in[40]; 
    assign layer_0[99] = ~(in[151] | in[150]); 
    assign layer_0[100] = in[85] | in[101]; 
    assign layer_0[101] = in[232] | in[90]; 
    assign layer_0[102] = ~in[135]; 
    assign layer_0[103] = in[90]; 
    assign layer_0[104] = in[185] | in[117]; 
    assign layer_0[105] = in[187] ^ in[101]; 
    assign layer_0[106] = in[84] ^ in[147]; 
    assign layer_0[107] = in[92] | in[90]; 
    assign layer_0[108] = in[90] | in[249]; 
    assign layer_0[109] = in[100] | in[91]; 
    assign layer_0[110] = in[33] | in[90]; 
    assign layer_0[111] = in[101] | in[115]; 
    assign layer_0[112] = in[92] | in[116]; 
    assign layer_0[113] = in[123] | in[139]; 
    assign layer_0[114] = ~in[216] | (in[216] & in[245]); 
    assign layer_0[115] = in[74]; 
    assign layer_0[116] = in[101]; 
    assign layer_0[117] = in[100] | in[101]; 
    assign layer_0[118] = in[90]; 
    assign layer_0[119] = in[116] | in[229]; 
    assign layer_0[120] = in[85]; 
    assign layer_0[121] = in[116] | in[99]; 
    assign layer_0[122] = ~in[135] | (in[247] & in[135]); 
    assign layer_0[123] = in[139]; 
    assign layer_0[124] = ~in[39]; 
    assign layer_0[125] = in[123]; 
    assign layer_0[126] = ~in[165] | (in[147] & in[165]); 
    assign layer_0[127] = in[90]; 
    assign layer_0[128] = in[99] | in[90]; 
    assign layer_0[129] = in[86] | in[147]; 
    assign layer_0[130] = in[86]; 
    assign layer_0[131] = in[246] ^ in[116]; 
    assign layer_0[132] = in[249] | in[107]; 
    assign layer_0[133] = in[164] ^ in[123]; 
    assign layer_0[134] = in[116] | in[116]; 
    assign layer_0[135] = in[141] | in[116]; 
    assign layer_0[136] = in[85]; 
    assign layer_0[137] = in[108] | in[90]; 
    assign layer_0[138] = in[132] | in[248]; 
    assign layer_0[139] = in[101] | in[99]; 
    assign layer_0[140] = in[26] | in[138]; 
    assign layer_0[141] = in[54] | in[170]; 
    assign layer_0[142] = in[100] | in[101]; 
    assign layer_0[143] = in[3] ^ in[75]; 
    assign layer_0[144] = in[139] | in[247]; 
    assign layer_0[145] = in[245] | in[132]; 
    assign layer_0[146] = in[101] & ~in[23]; 
    assign layer_0[147] = in[99] | in[101]; 
    assign layer_0[148] = in[93] | in[100]; 
    assign layer_0[149] = in[91] | in[92]; 
    assign layer_0[150] = in[157] ^ in[100]; 
    assign layer_0[151] = in[101] | in[92]; 
    assign layer_0[152] = in[131] | in[232]; 
    assign layer_0[153] = ~in[136] | (in[232] & in[136]); 
    assign layer_0[154] = in[91] & ~in[195]; 
    assign layer_0[155] = in[90] | in[247]; 
    assign layer_0[156] = in[90] | in[100]; 
    assign layer_0[157] = in[101] | in[115]; 
    assign layer_0[158] = in[101] | in[108]; 
    assign layer_0[159] = in[101] | in[125]; 
    assign layer_0[160] = in[90]; 
    assign layer_0[161] = in[99] | in[91]; 
    assign layer_0[162] = ~in[40]; 
    assign layer_0[163] = in[101]; 
    assign layer_0[164] = in[100] | in[75]; 
    assign layer_0[165] = in[91] | in[249]; 
    assign layer_0[166] = in[90] | in[93]; 
    assign layer_0[167] = in[247] | in[116]; 
    assign layer_0[168] = in[108] | in[106]; 
    assign layer_0[169] = in[90]; 
    assign layer_0[170] = in[108] | in[115]; 
    assign layer_0[171] = in[100] | in[117]; 
    assign layer_0[172] = in[91]; 
    assign layer_0[173] = in[91]; 
    assign layer_0[174] = in[90]; 
    assign layer_0[175] = in[22] | in[116]; 
    assign layer_0[176] = in[230] | in[90]; 
    assign layer_0[177] = in[69] | in[106]; 
    assign layer_0[178] = in[116]; 
    assign layer_0[179] = in[93] | in[85]; 
    assign layer_0[180] = in[100] ^ in[245]; 
    assign layer_0[181] = in[116] | in[117]; 
    assign layer_0[182] = in[229] | in[90]; 
    assign layer_0[183] = in[74] | in[147]; 
    assign layer_0[184] = in[116]; 
    assign layer_0[185] = in[91]; 
    assign layer_0[186] = in[76] | in[91]; 
    assign layer_0[187] = in[117] | in[116]; 
    assign layer_0[188] = in[116] | in[246]; 
    assign layer_0[189] = in[132] | in[228]; 
    assign layer_0[190] = in[75] | in[92]; 
    assign layer_0[191] = in[91]; 
    assign layer_0[192] = in[74] & ~in[40]; 
    assign layer_0[193] = in[116] | in[246]; 
    assign layer_0[194] = in[116] | in[117]; 
    assign layer_0[195] = in[107] & ~in[41]; 
    assign layer_0[196] = in[248] | in[132]; 
    assign layer_0[197] = in[91] | in[226]; 
    assign layer_0[198] = in[246] | in[116]; 
    assign layer_0[199] = ~in[182]; 
    assign layer_0[200] = in[245] | in[83]; 
    assign layer_0[201] = in[244] ^ in[116]; 
    assign layer_0[202] = in[149] | in[91]; 
    assign layer_0[203] = in[116] ^ in[248]; 
    assign layer_0[204] = in[100]; 
    assign layer_0[205] = in[116] | in[230]; 
    assign layer_0[206] = in[67] | in[91]; 
    assign layer_0[207] = ~in[119]; 
    assign layer_0[208] = ~(in[40] | in[42]); 
    assign layer_0[209] = in[101] | in[100]; 
    assign layer_0[210] = in[99]; 
    assign layer_0[211] = in[131] | in[101]; 
    assign layer_0[212] = in[246] | in[116]; 
    assign layer_0[213] = in[108]; 
    assign layer_0[214] = in[233] | in[91]; 
    assign layer_0[215] = in[116]; 
    assign layer_0[216] = in[117] | in[100]; 
    assign layer_0[217] = in[247] | in[132]; 
    assign layer_0[218] = in[91] | in[90]; 
    assign layer_0[219] = in[123] & ~in[38]; 
    assign layer_0[220] = in[133] ^ in[172]; 
    assign layer_0[221] = in[107]; 
    assign layer_0[222] = in[231] | in[116]; 
    assign layer_0[223] = in[101] ^ in[188]; 
    assign layer_0[224] = in[100]; 
    assign layer_0[225] = in[85] | in[93]; 
    assign layer_0[226] = in[90]; 
    assign layer_0[227] = in[75] | in[232]; 
    assign layer_0[228] = in[116] | in[108]; 
    assign layer_0[229] = in[106] & ~in[41]; 
    assign layer_0[230] = in[249] | in[230]; 
    assign layer_0[231] = in[138]; 
    assign layer_0[232] = in[91] | in[75]; 
    assign layer_0[233] = in[74] | in[233]; 
    assign layer_0[234] = in[230] | in[116]; 
    assign layer_0[235] = in[155] ^ in[133]; 
    assign layer_0[236] = in[27] | in[117]; 
    assign layer_0[237] = in[75]; 
    assign layer_0[238] = in[247] | in[132]; 
    assign layer_0[239] = in[187] ^ in[86]; 
    assign layer_0[240] = in[227] | in[154]; 
    assign layer_0[241] = in[90]; 
    assign layer_0[242] = in[117] ^ in[203]; 
    assign layer_0[243] = in[52] | in[116]; 
    assign layer_0[244] = ~in[152] | (in[152] & in[247]); 
    assign layer_0[245] = in[247] ^ in[148]; 
    assign layer_0[246] = in[132] | in[132]; 
    assign layer_0[247] = in[242] ^ in[116]; 
    assign layer_0[248] = in[172] ^ in[154]; 
    assign layer_0[249] = in[132] | in[247]; 
    assign layer_0[250] = ~(in[151] | in[152]); 
    assign layer_0[251] = in[247] | in[101]; 
    assign layer_0[252] = in[247] | in[116]; 
    assign layer_0[253] = in[85]; 
    assign layer_0[254] = in[231] | in[232]; 
    assign layer_0[255] = ~in[41] | (in[41] & in[108]); 
    assign layer_0[256] = in[109] | in[90]; 
    assign layer_0[257] = in[91] | in[74]; 
    assign layer_0[258] = in[233] | in[231]; 
    assign layer_0[259] = in[247] | in[90]; 
    assign layer_0[260] = in[86] | in[101]; 
    assign layer_0[261] = in[116] | in[247]; 
    assign layer_0[262] = in[247] | in[99]; 
    assign layer_0[263] = in[132] | in[92]; 
    assign layer_0[264] = in[99] | in[91]; 
    assign layer_0[265] = in[132] | in[246]; 
    assign layer_0[266] = in[248] | in[132]; 
    assign layer_0[267] = in[229] | in[248]; 
    assign layer_0[268] = in[85] ^ in[173]; 
    assign layer_0[269] = in[90] | in[231]; 
    assign layer_0[270] = in[75]; 
    assign layer_0[271] = ~in[40]; 
    assign layer_0[272] = in[117] | in[124]; 
    assign layer_0[273] = in[248] | in[117]; 
    assign layer_0[274] = in[100] | in[84]; 
    assign layer_0[275] = ~in[40]; 
    assign layer_0[276] = in[101] | in[116]; 
    assign layer_0[277] = in[75] | in[66]; 
    assign layer_0[278] = in[69] ^ in[154]; 
    assign layer_0[279] = in[91]; 
    assign layer_0[280] = in[230] | in[116]; 
    assign layer_0[281] = in[133] | in[132]; 
    assign layer_0[282] = in[91] | in[100]; 
    assign layer_0[283] = in[102] & ~in[51]; 
    assign layer_0[284] = in[52] | in[117]; 
    assign layer_0[285] = in[248] | in[100]; 
    assign layer_0[286] = in[67] | in[132]; 
    assign layer_0[287] = in[247] | in[116]; 
    assign layer_0[288] = in[90] | in[234]; 
    assign layer_0[289] = in[116] | in[246]; 
    assign layer_0[290] = in[74]; 
    assign layer_0[291] = in[116]; 
    assign layer_0[292] = in[248] ^ in[108]; 
    assign layer_0[293] = in[94] ^ in[138]; 
    assign layer_0[294] = in[90] | in[93]; 
    assign layer_0[295] = in[90]; 
    assign layer_0[296] = in[116] | in[132]; 
    assign layer_0[297] = in[230] | in[100]; 
    assign layer_0[298] = in[108] | in[108]; 
    assign layer_0[299] = in[101] ^ in[25]; 
    assign layer_0[300] = in[116] | in[116]; 
    assign layer_0[301] = ~(in[38] | in[119]); 
    assign layer_0[302] = in[246] | in[100]; 
    assign layer_0[303] = in[87] & ~in[39]; 
    assign layer_0[304] = in[138]; 
    assign layer_0[305] = in[100]; 
    assign layer_0[306] = in[132] | in[108]; 
    assign layer_0[307] = in[90]; 
    assign layer_0[308] = in[250] | in[108]; 
    assign layer_0[309] = in[85] | in[244]; 
    assign layer_0[310] = in[226] | in[101]; 
    assign layer_0[311] = in[101] | in[244]; 
    assign layer_0[312] = in[101] | in[116]; 
    assign layer_0[313] = in[116] | in[229]; 
    assign layer_0[314] = ~(in[186] | in[134]); 
    assign layer_0[315] = in[231] | in[116]; 
    assign layer_0[316] = in[133] | in[115]; 
    assign layer_0[317] = in[100] | in[93]; 
    assign layer_0[318] = ~(in[43] | in[41]); 
    assign layer_0[319] = in[90]; 
    assign layer_0[320] = ~in[150]; 
    assign layer_0[321] = in[156] ^ in[132]; 
    assign layer_0[322] = in[91] & ~in[24]; 
    assign layer_0[323] = in[116]; 
    assign layer_0[324] = in[91] | in[100]; 
    assign layer_0[325] = in[115] | in[75]; 
    assign layer_0[326] = in[217] | in[93]; 
    assign layer_0[327] = in[116] & ~in[79]; 
    assign layer_0[328] = in[90]; 
    assign layer_0[329] = in[116] | in[247]; 
    assign layer_0[330] = in[92] | in[74]; 
    assign layer_0[331] = in[100]; 
    assign layer_0[332] = in[116] | in[116]; 
    assign layer_0[333] = in[100] ^ in[93]; 
    assign layer_0[334] = in[91] | in[99]; 
    assign layer_0[335] = in[108] | in[101]; 
    assign layer_0[336] = in[100] | in[247]; 
    assign layer_0[337] = in[116] | in[91]; 
    assign layer_0[338] = in[108] ^ in[74]; 
    assign layer_0[339] = in[101]; 
    assign layer_0[340] = in[132]; 
    assign layer_0[341] = in[100] | in[92]; 
    assign layer_0[342] = ~in[135] | (in[135] & in[115]); 
    assign layer_0[343] = in[108] | in[116]; 
    assign layer_0[344] = ~in[167] | (in[167] & in[100]); 
    assign layer_0[345] = in[93] | in[76]; 
    assign layer_0[346] = in[91] | in[99]; 
    assign layer_0[347] = in[148] ^ in[247]; 
    assign layer_0[348] = in[132] | in[247]; 
    assign layer_0[349] = in[232] | in[108]; 
    assign layer_0[350] = in[132] | in[245]; 
    assign layer_0[351] = in[101]; 
    assign layer_0[352] = in[101] | in[116]; 
    assign layer_0[353] = in[138]; 
    assign layer_0[354] = ~in[119]; 
    assign layer_0[355] = in[74] ^ in[11]; 
    assign layer_0[356] = in[116] | in[115]; 
    assign layer_0[357] = in[101] | in[248]; 
    assign layer_0[358] = in[123] | in[25]; 
    assign layer_0[359] = in[90] | in[230]; 
    assign layer_0[360] = in[90]; 
    assign layer_0[361] = in[91]; 
    assign layer_0[362] = in[93] | in[116]; 
    assign layer_0[363] = in[90]; 
    assign layer_0[364] = in[132] | in[117]; 
    assign layer_0[365] = in[109] ^ in[107]; 
    assign layer_0[366] = in[100]; 
    assign layer_0[367] = in[100] | in[91]; 
    assign layer_0[368] = in[68] | in[124]; 
    assign layer_0[369] = in[116] | in[247]; 
    assign layer_0[370] = in[100] | in[91]; 
    assign layer_0[371] = in[227] | in[132]; 
    assign layer_0[372] = in[108] | in[101]; 
    assign layer_0[373] = in[100] | in[86]; 
    assign layer_0[374] = in[116] | in[91]; 
    assign layer_0[375] = in[67] | in[246]; 
    assign layer_0[376] = in[90]; 
    assign layer_0[377] = in[92]; 
    assign layer_0[378] = in[248] ^ in[116]; 
    assign layer_0[379] = in[116]; 
    assign layer_0[380] = in[229] | in[232]; 
    assign layer_0[381] = in[132] | in[26]; 
    assign layer_0[382] = ~in[151]; 
    assign layer_0[383] = ~in[40]; 
    assign layer_0[384] = in[91] | in[74]; 
    assign layer_0[385] = in[107] & ~in[42]; 
    assign layer_0[386] = in[100] | in[108]; 
    assign layer_0[387] = in[132] | in[246]; 
    assign layer_0[388] = ~in[167]; 
    assign layer_0[389] = in[148] ^ in[246]; 
    assign layer_0[390] = in[86]; 
    assign layer_0[391] = ~in[40]; 
    assign layer_0[392] = in[99] | in[108]; 
    assign layer_0[393] = in[131] | in[91]; 
    assign layer_0[394] = in[132] | in[229]; 
    assign layer_0[395] = in[91] | in[83]; 
    assign layer_0[396] = in[67] | in[90]; 
    assign layer_0[397] = in[231]; 
    assign layer_0[398] = in[69] & ~in[202]; 
    assign layer_0[399] = in[185] | in[187]; 
    assign layer_0[400] = in[92] | in[100]; 
    assign layer_0[401] = in[100] | in[108]; 
    assign layer_0[402] = in[101] | in[116]; 
    assign layer_0[403] = in[117]; 
    assign layer_0[404] = in[232] | in[91]; 
    assign layer_0[405] = in[108] | in[74]; 
    assign layer_0[406] = in[138] & ~in[150]; 
    assign layer_0[407] = in[101]; 
    assign layer_0[408] = in[69] ^ in[132]; 
    assign layer_0[409] = in[246] | in[116]; 
    assign layer_0[410] = in[90] | in[92]; 
    assign layer_0[411] = in[90]; 
    assign layer_0[412] = in[246] | in[116]; 
    assign layer_0[413] = in[100]; 
    assign layer_0[414] = in[90] & ~in[166]; 
    assign layer_0[415] = ~in[135]; 
    assign layer_0[416] = in[248] | in[91]; 
    assign layer_0[417] = in[75]; 
    assign layer_0[418] = in[90] | in[92]; 
    assign layer_0[419] = in[106] ^ in[109]; 
    assign layer_0[420] = in[246] | in[132]; 
    assign layer_0[421] = in[74] | in[94]; 
    assign layer_0[422] = in[116] | in[230]; 
    assign layer_0[423] = in[132] | in[92]; 
    assign layer_0[424] = in[172] ^ in[86]; 
    assign layer_0[425] = in[69] | in[116]; 
    assign layer_0[426] = in[86]; 
    assign layer_0[427] = ~in[166]; 
    assign layer_0[428] = in[108] | in[101]; 
    assign layer_0[429] = in[90]; 
    assign layer_0[430] = in[248] | in[230]; 
    assign layer_0[431] = in[75]; 
    assign layer_0[432] = in[91]; 
    assign layer_0[433] = in[155] | in[117]; 
    assign layer_0[434] = in[246] | in[131]; 
    assign layer_0[435] = in[91] | in[2]; 
    assign layer_0[436] = in[99] | in[91]; 
    assign layer_0[437] = in[116] | in[101]; 
    assign layer_0[438] = in[133] | in[92]; 
    assign layer_0[439] = in[231] | in[90]; 
    assign layer_0[440] = in[90]; 
    assign layer_0[441] = in[92] | in[90]; 
    assign layer_0[442] = in[213] | in[90]; 
    assign layer_0[443] = in[235] | in[234]; 
    assign layer_0[444] = ~in[136] | (in[136] & in[246]); 
    assign layer_0[445] = in[91]; 
    assign layer_0[446] = in[100] | in[109]; 
    assign layer_0[447] = in[84]; 
    assign layer_0[448] = ~in[39]; 
    assign layer_0[449] = in[90] | in[247]; 
    assign layer_0[450] = in[101] | in[115]; 
    assign layer_0[451] = in[74]; 
    assign layer_0[452] = in[116] | in[92]; 
    assign layer_0[453] = in[92] | in[91]; 
    assign layer_0[454] = in[245] | in[100]; 
    assign layer_0[455] = in[85] ^ in[172]; 
    assign layer_0[456] = in[232] | in[230]; 
    assign layer_0[457] = in[154] | in[53]; 
    assign layer_0[458] = in[246] | in[132]; 
    assign layer_0[459] = in[100] | in[230]; 
    assign layer_0[460] = in[106]; 
    assign layer_0[461] = in[116]; 
    assign layer_0[462] = in[247] | in[74]; 
    assign layer_0[463] = in[74] | in[83]; 
    assign layer_0[464] = in[232] | in[100]; 
    assign layer_0[465] = in[101] | in[116]; 
    assign layer_0[466] = in[75] | in[248]; 
    assign layer_0[467] = ~in[41]; 
    assign layer_0[468] = in[91] | in[116]; 
    assign layer_0[469] = in[116] | in[115]; 
    assign layer_0[470] = in[229] | in[248]; 
    assign layer_0[471] = in[75]; 
    assign layer_0[472] = in[248] | in[99]; 
    assign layer_0[473] = in[233] | in[90]; 
    assign layer_0[474] = in[116] | in[91]; 
    assign layer_0[475] = ~in[135] | (in[248] & in[135]); 
    assign layer_0[476] = in[91] | in[99]; 
    assign layer_0[477] = in[90]; 
    assign layer_0[478] = in[116] | in[101]; 
    assign layer_0[479] = in[100] & ~in[189]; 
    assign layer_0[480] = in[115] | in[91]; 
    assign layer_0[481] = in[86] & ~in[39]; 
    assign layer_0[482] = in[230] | in[232]; 
    assign layer_0[483] = in[116] | in[247]; 
    assign layer_0[484] = in[76] | in[91]; 
    assign layer_0[485] = in[138] & ~in[179]; 
    assign layer_0[486] = in[90] | in[231]; 
    assign layer_0[487] = in[116]; 
    assign layer_0[488] = in[100]; 
    assign layer_0[489] = in[90] ^ in[192]; 
    assign layer_0[490] = in[108] | in[132]; 
    assign layer_0[491] = in[91] | in[92]; 
    assign layer_0[492] = in[100]; 
    assign layer_0[493] = in[91] | in[165]; 
    assign layer_0[494] = ~in[40]; 
    assign layer_0[495] = in[94] ^ in[106]; 
    assign layer_0[496] = in[90]; 
    assign layer_0[497] = in[115] | in[91]; 
    assign layer_0[498] = in[101] | in[99]; 
    assign layer_0[499] = ~in[88] | (in[88] & in[108]); 
    assign layer_0[500] = in[247] ^ in[83]; 
    assign layer_0[501] = in[116] | in[116]; 
    assign layer_0[502] = in[102]; 
    assign layer_0[503] = in[75]; 
    assign layer_0[504] = in[115] | in[91]; 
    assign layer_0[505] = in[124] | in[101]; 
    assign layer_0[506] = in[179] | in[155]; 
    assign layer_0[507] = in[247] | in[116]; 
    assign layer_0[508] = in[91] & ~in[37]; 
    assign layer_0[509] = in[100] | in[108]; 
    assign layer_0[510] = in[116] | in[101]; 
    assign layer_0[511] = in[154]; 
    assign layer_0[512] = in[100] | in[116]; 
    assign layer_0[513] = in[108] | in[70]; 
    assign layer_0[514] = ~in[150] | (in[150] & in[116]); 
    assign layer_0[515] = in[132] | in[246]; 
    assign layer_0[516] = in[100] ^ in[230]; 
    assign layer_0[517] = in[246] | in[132]; 
    assign layer_0[518] = in[219] | in[68]; 
    assign layer_0[519] = in[115] | in[116]; 
    assign layer_0[520] = in[117] ^ in[156]; 
    assign layer_0[521] = in[247] | in[74]; 
    assign layer_0[522] = in[116] | in[100]; 
    assign layer_0[523] = ~in[119] | (in[116] & in[119]); 
    assign layer_0[524] = in[116] | in[245]; 
    assign layer_0[525] = in[22] ^ in[116]; 
    assign layer_0[526] = ~in[135] | (in[135] & in[115]); 
    assign layer_0[527] = in[117]; 
    assign layer_0[528] = in[154] | in[70]; 
    assign layer_0[529] = ~in[41]; 
    assign layer_0[530] = in[100] | in[101]; 
    assign layer_0[531] = in[158] ^ in[85]; 
    assign layer_0[532] = in[149] | in[85]; 
    assign layer_0[533] = ~in[136]; 
    assign layer_0[534] = ~in[135] | (in[135] & in[101]); 
    assign layer_0[535] = in[100] & ~in[128]; 
    assign layer_0[536] = in[83] | in[101]; 
    assign layer_0[537] = in[75] | in[74]; 
    assign layer_0[538] = in[230] | in[233]; 
    assign layer_0[539] = in[98] | in[101]; 
    assign layer_0[540] = in[109] | in[116]; 
    assign layer_0[541] = ~in[150] | (in[150] & in[250]); 
    assign layer_0[542] = in[222] | in[101]; 
    assign layer_0[543] = in[107]; 
    assign layer_0[544] = ~in[166] | (in[166] & in[92]); 
    assign layer_0[545] = ~in[41]; 
    assign layer_0[546] = in[117] | in[186]; 
    assign layer_0[547] = in[91] & ~in[38]; 
    assign layer_0[548] = in[247] | in[116]; 
    assign layer_0[549] = in[92]; 
    assign layer_0[550] = in[75] | in[100]; 
    assign layer_0[551] = in[92] | in[247]; 
    assign layer_0[552] = in[124] | in[117]; 
    assign layer_0[553] = in[91]; 
    assign layer_0[554] = ~in[135]; 
    assign layer_0[555] = ~in[165] | (in[165] & in[94]); 
    assign layer_0[556] = in[101] | in[101]; 
    assign layer_0[557] = in[116] | in[116]; 
    assign layer_0[558] = in[91]; 
    assign layer_0[559] = in[90] | in[93]; 
    assign layer_0[560] = in[117] | in[116]; 
    assign layer_0[561] = in[74] | in[249]; 
    assign layer_0[562] = in[116] | in[245]; 
    assign layer_0[563] = in[115] | in[91]; 
    assign layer_0[564] = in[101]; 
    assign layer_0[565] = in[102]; 
    assign layer_0[566] = in[147] | in[247]; 
    assign layer_0[567] = ~(in[233] | in[136]); 
    assign layer_0[568] = in[74]; 
    assign layer_0[569] = in[91]; 
    assign layer_0[570] = ~in[40]; 
    assign layer_0[571] = in[228] | in[247]; 
    assign layer_0[572] = in[91] & ~in[180]; 
    assign layer_0[573] = ~in[168] | (in[212] & in[168]); 
    assign layer_0[574] = in[117] | in[116]; 
    assign layer_0[575] = in[75] | in[67]; 
    assign layer_0[576] = in[99] | in[116]; 
    assign layer_0[577] = in[102] | in[123]; 
    assign layer_0[578] = in[88]; 
    assign layer_0[579] = in[84] | in[100]; 
    assign layer_0[580] = in[84] ^ in[107]; 
    assign layer_0[581] = ~in[103] | (in[173] & in[103]); 
    assign layer_0[582] = ~in[39]; 
    assign layer_0[583] = in[116] | in[68]; 
    assign layer_0[584] = in[230] | in[116]; 
    assign layer_0[585] = in[115] | in[116]; 
    assign layer_0[586] = in[91] | in[232]; 
    assign layer_0[587] = in[108] | in[116]; 
    assign layer_0[588] = in[99] ^ in[92]; 
    assign layer_0[589] = ~in[135] | (in[135] & in[97]); 
    assign layer_0[590] = in[248] | in[116]; 
    assign layer_0[591] = in[92] | in[100]; 
    assign layer_0[592] = in[91] | in[231]; 
    assign layer_0[593] = in[131] | in[230]; 
    assign layer_0[594] = in[100] | in[92]; 
    assign layer_0[595] = in[116] | in[101]; 
    assign layer_0[596] = ~in[150]; 
    assign layer_0[597] = in[73] & ~in[43]; 
    assign layer_0[598] = in[90] | in[109]; 
    assign layer_0[599] = in[93] | in[90]; 
    assign layer_0[600] = in[116]; 
    assign layer_0[601] = in[92] | in[100]; 
    assign layer_0[602] = in[84] | in[74]; 
    assign layer_0[603] = in[101] | in[101]; 
    assign layer_0[604] = in[231] | in[115]; 
    assign layer_0[605] = ~in[166] | (in[166] & in[230]); 
    assign layer_0[606] = ~in[40]; 
    assign layer_0[607] = in[132] | in[117]; 
    assign layer_0[608] = in[116] | in[117]; 
    assign layer_0[609] = in[230] | in[83]; 
    assign layer_0[610] = ~in[39] | (in[39] & in[246]); 
    assign layer_0[611] = in[101] | in[99]; 
    assign layer_0[612] = in[91] | in[147]; 
    assign layer_0[613] = in[91]; 
    assign layer_0[614] = in[132] | in[147]; 
    assign layer_0[615] = in[90] | in[30]; 
    assign layer_0[616] = in[131] | in[101]; 
    assign layer_0[617] = in[102]; 
    assign layer_0[618] = in[91] | in[232]; 
    assign layer_0[619] = in[246] | in[132]; 
    assign layer_0[620] = in[85] & ~in[40]; 
    assign layer_0[621] = in[131] | in[82]; 
    assign layer_0[622] = in[84] | in[229]; 
    assign layer_0[623] = ~in[40]; 
    assign layer_0[624] = in[90]; 
    assign layer_0[625] = in[116] | in[116]; 
    assign layer_0[626] = in[74] | in[74]; 
    assign layer_0[627] = in[132] | in[124]; 
    assign layer_0[628] = in[100]; 
    assign layer_0[629] = in[244] | in[117]; 
    assign layer_0[630] = ~in[39]; 
    assign layer_0[631] = in[101] | in[84]; 
    assign layer_0[632] = in[116] | in[108]; 
    assign layer_0[633] = in[232] | in[116]; 
    assign layer_0[634] = ~in[151] | (in[247] & in[151]); 
    assign layer_0[635] = in[248] | in[101]; 
    assign layer_0[636] = in[246] | in[115]; 
    assign layer_0[637] = in[187] ^ in[86]; 
    assign layer_0[638] = in[116] | in[127]; 
    assign layer_0[639] = in[84] & ~in[197]; 
    assign layer_0[640] = in[132] | in[247]; 
    assign layer_0[641] = in[52] | in[116]; 
    assign layer_0[642] = in[99] | in[230]; 
    assign layer_0[643] = in[90]; 
    assign layer_0[644] = in[101]; 
    assign layer_0[645] = in[139] | in[101]; 
    assign layer_0[646] = in[116] | in[116]; 
    assign layer_0[647] = in[132] ^ in[246]; 
    assign layer_0[648] = in[247] | in[250]; 
    assign layer_0[649] = in[85]; 
    assign layer_0[650] = in[116] | in[244]; 
    assign layer_0[651] = ~in[135]; 
    assign layer_0[652] = in[115] | in[101]; 
    assign layer_0[653] = in[100] | in[230]; 
    assign layer_0[654] = in[116] | in[83]; 
    assign layer_0[655] = in[116] ^ in[246]; 
    assign layer_0[656] = in[116] | in[102]; 
    assign layer_0[657] = in[106] | in[99]; 
    assign layer_0[658] = in[92] | in[90]; 
    assign layer_0[659] = in[83] | in[91]; 
    assign layer_0[660] = in[100] | in[92]; 
    assign layer_0[661] = in[108] | in[100]; 
    assign layer_0[662] = in[90]; 
    assign layer_0[663] = in[86]; 
    assign layer_0[664] = in[132] | in[101]; 
    assign layer_0[665] = in[117] | in[115]; 
    assign layer_0[666] = in[101] | in[108]; 
    assign layer_0[667] = in[132]; 
    assign layer_0[668] = in[108] | in[116]; 
    assign layer_0[669] = in[115] | in[101]; 
    assign layer_0[670] = in[246] | in[91]; 
    assign layer_0[671] = in[90]; 
    assign layer_0[672] = in[172] ^ in[139]; 
    assign layer_0[673] = in[117] | in[100]; 
    assign layer_0[674] = in[116] | in[108]; 
    assign layer_0[675] = in[69] & ~in[203]; 
    assign layer_0[676] = in[101] | in[115]; 
    assign layer_0[677] = in[131] | in[246]; 
    assign layer_0[678] = in[91] | in[100]; 
    assign layer_0[679] = in[116]; 
    assign layer_0[680] = in[246] | in[85]; 
    assign layer_0[681] = ~(in[151] | in[235]); 
    assign layer_0[682] = in[90] | in[92]; 
    assign layer_0[683] = in[109] | in[100]; 
    assign layer_0[684] = ~in[166]; 
    assign layer_0[685] = in[69]; 
    assign layer_0[686] = in[68] | in[116]; 
    assign layer_0[687] = in[102] & ~in[39]; 
    assign layer_0[688] = in[101] | in[67]; 
    assign layer_0[689] = in[124] | in[100]; 
    assign layer_0[690] = in[230] | in[70]; 
    assign layer_0[691] = in[90] | in[92]; 
    assign layer_0[692] = in[91] | in[234]; 
    assign layer_0[693] = in[247] | in[116]; 
    assign layer_0[694] = in[91]; 
    assign layer_0[695] = in[116] | in[248]; 
    assign layer_0[696] = in[231] | in[90]; 
    assign layer_0[697] = in[116] | in[69]; 
    assign layer_0[698] = in[131] | in[101]; 
    assign layer_0[699] = in[74]; 
    assign layer_0[700] = in[90] ^ in[93]; 
    assign layer_0[701] = in[91]; 
    assign layer_0[702] = in[149] ^ in[107]; 
    assign layer_0[703] = in[100] | in[116]; 
    assign layer_0[704] = in[86] | in[95]; 
    assign layer_0[705] = in[100] | in[230]; 
    assign layer_0[706] = ~(in[57] ^ in[71]); 
    assign layer_0[707] = in[90] | in[52]; 
    assign layer_0[708] = in[116] ^ in[25]; 
    assign layer_0[709] = in[169]; 
    assign layer_0[710] = ~in[182]; 
    assign layer_0[711] = in[100] | in[248]; 
    assign layer_0[712] = ~in[135]; 
    assign layer_0[713] = in[116] | in[101]; 
    assign layer_0[714] = in[102] | in[94]; 
    assign layer_0[715] = in[90] | in[76]; 
    assign layer_0[716] = in[75]; 
    assign layer_0[717] = in[132] | in[247]; 
    assign layer_0[718] = in[132] | in[124]; 
    assign layer_0[719] = ~in[151]; 
    assign layer_0[720] = in[101]; 
    assign layer_0[721] = in[93] | in[90]; 
    assign layer_0[722] = in[90] | in[75]; 
    assign layer_0[723] = in[84] | in[92]; 
    assign layer_0[724] = ~in[40]; 
    assign layer_0[725] = ~in[151]; 
    assign layer_0[726] = in[107]; 
    assign layer_0[727] = in[101]; 
    assign layer_0[728] = in[231] | in[147]; 
    assign layer_0[729] = in[116] | in[99]; 
    assign layer_0[730] = in[92] | in[132]; 
    assign layer_0[731] = in[117] | in[115]; 
    assign layer_0[732] = in[132] | in[132]; 
    assign layer_0[733] = in[101] | in[100]; 
    assign layer_0[734] = in[245] | in[132]; 
    assign layer_0[735] = in[170] | in[108]; 
    assign layer_0[736] = in[92] | in[90]; 
    assign layer_0[737] = in[99] | in[91]; 
    assign layer_0[738] = ~in[119] | (in[247] & in[119]); 
    assign layer_0[739] = in[92] ^ in[90]; 
    assign layer_0[740] = in[229] | in[248]; 
    assign layer_0[741] = in[116] | in[108]; 
    assign layer_0[742] = in[101] | in[247]; 
    assign layer_0[743] = ~in[39]; 
    assign layer_0[744] = in[91]; 
    assign layer_0[745] = in[116] | in[245]; 
    assign layer_0[746] = in[91] | in[132]; 
    assign layer_0[747] = ~in[150] | (in[115] & in[150]); 
    assign layer_0[748] = in[83]; 
    assign layer_0[749] = in[132]; 
    assign layer_0[750] = in[100] | in[58]; 
    assign layer_0[751] = in[187] ^ in[117]; 
    assign layer_0[752] = in[90] | in[93]; 
    assign layer_0[753] = in[84] | in[91]; 
    assign layer_0[754] = in[99] | in[117]; 
    assign layer_0[755] = in[109] ^ in[232]; 
    assign layer_0[756] = ~in[182]; 
    assign layer_0[757] = in[247] | in[117]; 
    assign layer_0[758] = in[123]; 
    assign layer_0[759] = in[246] | in[132]; 
    assign layer_0[760] = in[75] & ~in[242]; 
    assign layer_0[761] = in[156] ^ in[117]; 
    assign layer_0[762] = in[247] | in[100]; 
    assign layer_0[763] = in[132] | in[107]; 
    assign layer_0[764] = in[245] | in[116]; 
    assign layer_0[765] = ~in[182]; 
    assign layer_0[766] = in[91] | in[115]; 
    assign layer_0[767] = in[101] | in[100]; 
    assign layer_0[768] = ~(in[135] | in[166]); 
    assign layer_0[769] = in[91]; 
    assign layer_0[770] = ~in[167] | (in[167] & in[75]); 
    assign layer_0[771] = in[91]; 
    assign layer_0[772] = in[74] | in[75]; 
    assign layer_0[773] = in[101]; 
    assign layer_0[774] = in[90]; 
    assign layer_0[775] = in[117] | in[109]; 
    assign layer_0[776] = ~in[182]; 
    assign layer_0[777] = in[246] | in[132]; 
    assign layer_0[778] = in[91] | in[232]; 
    assign layer_0[779] = ~in[40]; 
    assign layer_0[780] = ~in[150] | (in[150] & in[247]); 
    assign layer_0[781] = in[117] & ~in[52]; 
    assign layer_0[782] = in[83]; 
    assign layer_0[783] = in[108] | in[101]; 
    assign layer_0[784] = in[101] ^ in[128]; 
    assign layer_0[785] = in[100] | in[108]; 
    assign layer_0[786] = in[86]; 
    assign layer_0[787] = in[116]; 
    assign layer_0[788] = in[172] ^ in[117]; 
    assign layer_0[789] = in[90]; 
    assign layer_0[790] = in[100] | in[92]; 
    assign layer_0[791] = in[91] | in[99]; 
    assign layer_0[792] = ~in[151] | (in[249] & in[151]); 
    assign layer_0[793] = ~in[135]; 
    assign layer_0[794] = in[230] | in[100]; 
    assign layer_0[795] = in[92] | in[116]; 
    assign layer_0[796] = in[248] ^ in[108]; 
    assign layer_0[797] = in[116] | in[100]; 
    assign layer_0[798] = in[100] | in[68]; 
    assign layer_0[799] = ~in[41]; 
    assign layer_0[800] = in[91] | in[68]; 
    assign layer_0[801] = in[99] | in[101]; 
    assign layer_0[802] = in[100] | in[230]; 
    assign layer_0[803] = in[156] ^ in[116]; 
    assign layer_0[804] = in[70] | in[78]; 
    assign layer_0[805] = in[116] | in[116]; 
    assign layer_0[806] = in[117] & ~in[187]; 
    assign layer_0[807] = in[171] | in[117]; 
    assign layer_0[808] = in[147] | in[117]; 
    assign layer_0[809] = in[100]; 
    assign layer_0[810] = in[90] | in[92]; 
    assign layer_0[811] = in[116]; 
    assign layer_0[812] = in[117] | in[70]; 
    assign layer_0[813] = in[116] | in[245]; 
    assign layer_0[814] = in[116] | in[70]; 
    assign layer_0[815] = in[90]; 
    assign layer_0[816] = ~in[39]; 
    assign layer_0[817] = in[116]; 
    assign layer_0[818] = in[115] | in[102]; 
    assign layer_0[819] = in[52] | in[155]; 
    assign layer_0[820] = ~(in[167] & in[166]); 
    assign layer_0[821] = in[91] | in[92]; 
    assign layer_0[822] = in[116]; 
    assign layer_0[823] = ~in[119]; 
    assign layer_0[824] = in[154]; 
    assign layer_0[825] = in[132] | in[76]; 
    assign layer_0[826] = in[52] | in[91]; 
    assign layer_0[827] = in[101] | in[115]; 
    assign layer_0[828] = in[100]; 
    assign layer_0[829] = in[116] | in[108]; 
    assign layer_0[830] = in[229] | in[116]; 
    assign layer_0[831] = in[101] | in[52]; 
    assign layer_0[832] = in[90]; 
    assign layer_0[833] = in[91] | in[77]; 
    assign layer_0[834] = in[132] | in[246]; 
    assign layer_0[835] = in[133]; 
    assign layer_0[836] = in[84] | in[108]; 
    assign layer_0[837] = in[91]; 
    assign layer_0[838] = in[107] | in[115]; 
    assign layer_0[839] = in[101]; 
    assign layer_0[840] = in[115] | in[230]; 
    assign layer_0[841] = in[116] | in[92]; 
    assign layer_0[842] = in[91]; 
    assign layer_0[843] = in[74] | in[68]; 
    assign layer_0[844] = in[90] | in[75]; 
    assign layer_0[845] = in[233] | in[75]; 
    assign layer_0[846] = in[117] | in[116]; 
    assign layer_0[847] = in[115] | in[91]; 
    assign layer_0[848] = in[132] | in[124]; 
    assign layer_0[849] = in[90] & ~in[23]; 
    assign layer_0[850] = in[247] | in[116]; 
    assign layer_0[851] = in[154] ^ in[241]; 
    assign layer_0[852] = in[138]; 
    assign layer_0[853] = in[75] | in[90]; 
    assign layer_0[854] = in[45] ^ in[91]; 
    assign layer_0[855] = in[115] | in[117]; 
    assign layer_0[856] = in[74] | in[248]; 
    assign layer_0[857] = ~in[151]; 
    assign layer_0[858] = in[115] | in[117]; 
    assign layer_0[859] = in[117] ^ in[171]; 
    assign layer_0[860] = in[90] | in[93]; 
    assign layer_0[861] = ~(in[136] | in[235]); 
    assign layer_0[862] = in[248] | in[132]; 
    assign layer_0[863] = in[132] | in[248]; 
    assign layer_0[864] = in[248] | in[132]; 
    assign layer_0[865] = in[91]; 
    assign layer_0[866] = ~in[120] | (in[120] & in[132]); 
    assign layer_0[867] = in[247] | in[132]; 
    assign layer_0[868] = in[92] | in[54]; 
    assign layer_0[869] = in[74] | in[123]; 
    assign layer_0[870] = ~in[166] | (in[166] & in[247]); 
    assign layer_0[871] = in[92] | in[90]; 
    assign layer_0[872] = in[116] | in[247]; 
    assign layer_0[873] = ~(in[151] | in[208]); 
    assign layer_0[874] = in[132] | in[163]; 
    assign layer_0[875] = in[101]; 
    assign layer_0[876] = in[84] | in[132]; 
    assign layer_0[877] = in[76] | in[218]; 
    assign layer_0[878] = in[101] | in[100]; 
    assign layer_0[879] = in[116]; 
    assign layer_0[880] = in[91]; 
    assign layer_0[881] = in[74] | in[75]; 
    assign layer_0[882] = in[117] ^ in[187]; 
    assign layer_0[883] = in[91] | in[92]; 
    assign layer_0[884] = ~in[135] | (in[247] & in[135]); 
    assign layer_0[885] = in[248] | in[91]; 
    assign layer_0[886] = in[90]; 
    assign layer_0[887] = in[213] | in[232]; 
    assign layer_0[888] = in[101] | in[109]; 
    assign layer_0[889] = in[133] | in[148]; 
    assign layer_0[890] = in[101] | in[164]; 
    assign layer_0[891] = in[90]; 
    assign layer_0[892] = in[247] | in[234]; 
    assign layer_0[893] = in[9] | in[90]; 
    assign layer_0[894] = in[62] | in[86]; 
    assign layer_0[895] = in[101]; 
    assign layer_0[896] = in[156] ^ in[123]; 
    assign layer_0[897] = in[83] | in[68]; 
    assign layer_0[898] = in[169] & ~in[181]; 
    assign layer_0[899] = in[84]; 
    assign layer_0[900] = in[123] & ~in[141]; 
    assign layer_0[901] = in[116] | in[90]; 
    assign layer_0[902] = in[116]; 
    assign layer_0[903] = in[116] | in[147]; 
    assign layer_0[904] = in[164] | in[116]; 
    assign layer_0[905] = in[116] | in[117]; 
    assign layer_0[906] = in[154] | in[139]; 
    assign layer_0[907] = in[101] | in[101]; 
    assign layer_0[908] = in[246] | in[100]; 
    assign layer_0[909] = in[246] | in[75]; 
    assign layer_0[910] = ~in[40] | (in[40] & in[125]); 
    assign layer_0[911] = in[116] | in[108]; 
    assign layer_0[912] = in[246]; 
    assign layer_0[913] = in[132] | in[92]; 
    assign layer_0[914] = in[85]; 
    assign layer_0[915] = in[107] & ~in[44]; 
    assign layer_0[916] = in[101]; 
    assign layer_0[917] = in[115] | in[230]; 
    assign layer_0[918] = in[86]; 
    assign layer_0[919] = in[117]; 
    assign layer_0[920] = in[91] | in[108]; 
    assign layer_0[921] = in[132] | in[108]; 
    assign layer_0[922] = in[116] | in[98]; 
    assign layer_0[923] = in[106] | in[246]; 
    assign layer_0[924] = in[90] | in[248]; 
    assign layer_0[925] = in[117]; 
    assign layer_0[926] = in[116]; 
    assign layer_0[927] = ~(in[41] | in[42]); 
    assign layer_0[928] = in[74] | in[75]; 
    assign layer_0[929] = in[245] | in[116]; 
    assign layer_0[930] = in[92] | in[90]; 
    assign layer_0[931] = in[101]; 
    assign layer_0[932] = in[91]; 
    assign layer_0[933] = in[123] | in[248]; 
    assign layer_0[934] = in[101] | in[100]; 
    assign layer_0[935] = in[91] | in[90]; 
    assign layer_0[936] = in[132] | in[101]; 
    assign layer_0[937] = in[116]; 
    assign layer_0[938] = in[233] | in[92]; 
    assign layer_0[939] = in[100] ^ in[117]; 
    assign layer_0[940] = in[91]; 
    assign layer_0[941] = in[92] | in[247]; 
    assign layer_0[942] = in[84] | in[75]; 
    assign layer_0[943] = in[100] | in[99]; 
    assign layer_0[944] = in[231] | in[108]; 
    assign layer_0[945] = ~in[121]; 
    assign layer_0[946] = ~(in[151] | in[234]); 
    assign layer_0[947] = in[232] | in[90]; 
    assign layer_0[948] = in[154]; 
    assign layer_0[949] = in[92] | in[91]; 
    assign layer_0[950] = in[85] & ~in[25]; 
    assign layer_0[951] = in[90]; 
    assign layer_0[952] = in[230] | in[116]; 
    assign layer_0[953] = in[90] & ~in[39]; 
    assign layer_0[954] = in[116]; 
    assign layer_0[955] = in[38] ^ in[86]; 
    assign layer_0[956] = in[123] | in[156]; 
    assign layer_0[957] = in[83] | in[245]; 
    assign layer_0[958] = in[132]; 
    assign layer_0[959] = in[213] | in[74]; 
    assign layer_0[960] = in[86] | in[26]; 
    assign layer_0[961] = in[92]; 
    assign layer_0[962] = in[88] & ~in[188]; 
    assign layer_0[963] = in[75] | in[94]; 
    assign layer_0[964] = in[247] | in[132]; 
    assign layer_0[965] = in[90]; 
    assign layer_0[966] = in[101] | in[204]; 
    assign layer_0[967] = in[74]; 
    assign layer_0[968] = in[100] | in[248]; 
    assign layer_0[969] = in[248] ^ in[132]; 
    assign layer_0[970] = ~in[166] | (in[166] & in[233]); 
    assign layer_0[971] = ~in[151]; 
    assign layer_0[972] = in[229] | in[116]; 
    assign layer_0[973] = in[90]; 
    assign layer_0[974] = in[91]; 
    assign layer_0[975] = in[116]; 
    assign layer_0[976] = in[99] | in[232]; 
    assign layer_0[977] = in[90]; 
    assign layer_0[978] = in[117] | in[124]; 
    assign layer_0[979] = in[101]; 
    assign layer_0[980] = in[148] | in[123]; 
    assign layer_0[981] = in[232] ^ in[229]; 
    assign layer_0[982] = ~in[135]; 
    assign layer_0[983] = in[154]; 
    assign layer_0[984] = in[117] | in[116]; 
    assign layer_0[985] = in[247] | in[116]; 
    assign layer_0[986] = in[132] | in[247]; 
    assign layer_0[987] = in[90] | in[91]; 
    assign layer_0[988] = in[74]; 
    assign layer_0[989] = in[248] | in[92]; 
    assign layer_0[990] = in[154] ^ in[53]; 
    assign layer_0[991] = in[68] | in[117]; 
    assign layer_0[992] = in[101]; 
    assign layer_0[993] = in[231] | in[99]; 
    assign layer_0[994] = in[101]; 
    assign layer_0[995] = ~in[182] | (in[92] & in[182]); 
    assign layer_0[996] = in[92] ^ in[89]; 
    assign layer_0[997] = in[117] & ~in[94]; 
    assign layer_0[998] = in[237] | in[91]; 
    assign layer_0[999] = in[116] | in[246]; 
    assign layer_0[1000] = in[132]; 
    assign layer_0[1001] = in[90]; 
    assign layer_0[1002] = in[132] | in[115]; 
    assign layer_0[1003] = in[117] | in[67]; 
    assign layer_0[1004] = in[84]; 
    assign layer_0[1005] = in[100]; 
    assign layer_0[1006] = in[116] | in[115]; 
    assign layer_0[1007] = in[86] & ~in[173]; 
    assign layer_0[1008] = ~in[40] | (in[92] & in[40]); 
    assign layer_0[1009] = in[116] | in[101]; 
    assign layer_0[1010] = in[247] | in[100]; 
    assign layer_0[1011] = in[102] | in[115]; 
    assign layer_0[1012] = in[101]; 
    assign layer_0[1013] = in[90]; 
    assign layer_0[1014] = in[116]; 
    assign layer_0[1015] = in[89] & ~in[41]; 
    assign layer_0[1016] = in[247] | in[116]; 
    assign layer_0[1017] = in[108] | in[101]; 
    assign layer_0[1018] = ~in[40]; 
    assign layer_0[1019] = in[90]; 
    assign layer_0[1020] = in[91]; 
    assign layer_0[1021] = ~in[135]; 
    assign layer_0[1022] = in[92] ^ in[45]; 
    assign layer_0[1023] = ~in[135]; 
    assign layer_0[1024] = in[86]; 
    assign layer_0[1025] = in[91]; 
    assign layer_0[1026] = in[74] | in[76]; 
    assign layer_0[1027] = ~in[40]; 
    assign layer_0[1028] = in[99] | in[75]; 
    assign layer_0[1029] = ~(in[39] | in[42]); 
    assign layer_0[1030] = in[116]; 
    assign layer_0[1031] = in[247] | in[101]; 
    assign layer_0[1032] = in[84] | in[101]; 
    assign layer_0[1033] = in[101] | in[124]; 
    assign layer_0[1034] = in[84] | in[229]; 
    assign layer_0[1035] = in[101] | in[109]; 
    assign layer_0[1036] = in[101]; 
    assign layer_0[1037] = ~in[166]; 
    assign layer_0[1038] = in[90]; 
    assign layer_0[1039] = in[131] | in[101]; 
    assign layer_0[1040] = in[90]; 
    assign layer_0[1041] = in[91] | in[249]; 
    assign layer_0[1042] = in[246] | in[84]; 
    assign layer_0[1043] = in[70]; 
    assign layer_0[1044] = in[116] | in[247]; 
    assign layer_0[1045] = in[149] | in[148]; 
    assign layer_0[1046] = ~in[105] | (in[77] & in[105]); 
    assign layer_0[1047] = in[116] | in[246]; 
    assign layer_0[1048] = in[106] | in[109]; 
    assign layer_0[1049] = in[100] | in[70]; 
    assign layer_0[1050] = in[131] ^ in[248]; 
    assign layer_0[1051] = in[101] | in[92]; 
    assign layer_0[1052] = in[91] | in[77]; 
    assign layer_0[1053] = in[90] | in[115]; 
    assign layer_0[1054] = in[234] | in[132]; 
    assign layer_0[1055] = in[85]; 
    assign layer_0[1056] = in[90] | in[91]; 
    assign layer_0[1057] = in[116] | in[247]; 
    assign layer_0[1058] = in[116]; 
    assign layer_0[1059] = in[154] ^ in[156]; 
    assign layer_0[1060] = in[92] | in[101]; 
    assign layer_0[1061] = in[67] | in[108]; 
    assign layer_0[1062] = in[75]; 
    assign layer_0[1063] = in[92] | in[106]; 
    assign layer_0[1064] = in[139]; 
    assign layer_0[1065] = in[71] | in[132]; 
    assign layer_0[1066] = in[132] | in[230]; 
    assign layer_0[1067] = in[89] ^ in[76]; 
    assign layer_0[1068] = in[124] | in[116]; 
    assign layer_0[1069] = in[85]; 
    assign layer_0[1070] = in[124] | in[116]; 
    assign layer_0[1071] = in[248] | in[116]; 
    assign layer_0[1072] = in[116] | in[247]; 
    assign layer_0[1073] = in[132] | in[154]; 
    assign layer_0[1074] = in[90]; 
    assign layer_0[1075] = in[101]; 
    assign layer_0[1076] = in[90] | in[116]; 
    assign layer_0[1077] = in[230] | in[132]; 
    assign layer_0[1078] = in[99] | in[101]; 
    assign layer_0[1079] = in[185] | in[71]; 
    assign layer_0[1080] = in[132] | in[132]; 
    assign layer_0[1081] = in[101] | in[99]; 
    assign layer_0[1082] = in[75] & ~in[41]; 
    assign layer_0[1083] = in[76] | in[74]; 
    assign layer_0[1084] = in[117] & ~in[23]; 
    assign layer_0[1085] = in[75]; 
    assign layer_0[1086] = in[247] | in[74]; 
    assign layer_0[1087] = in[100] | in[86]; 
    assign layer_0[1088] = in[93] ^ in[90]; 
    assign layer_0[1089] = in[132] | in[247]; 
    assign layer_0[1090] = in[90]; 
    assign layer_0[1091] = in[74] | in[75]; 
    assign layer_0[1092] = in[171] ^ in[101]; 
    assign layer_0[1093] = in[108] | in[116]; 
    assign layer_0[1094] = in[115] | in[20]; 
    assign layer_0[1095] = in[248] | in[246]; 
    assign layer_0[1096] = in[245] | in[132]; 
    assign layer_0[1097] = in[91] | in[100]; 
    assign layer_0[1098] = ~in[40]; 
    assign layer_0[1099] = in[156] ^ in[101]; 
    assign layer_0[1100] = in[116] ^ in[143]; 
    assign layer_0[1101] = in[245] | in[132]; 
    assign layer_0[1102] = in[116] | in[247]; 
    assign layer_0[1103] = in[232] | in[91]; 
    assign layer_0[1104] = in[117] ^ in[172]; 
    assign layer_0[1105] = in[107]; 
    assign layer_0[1106] = in[90] | in[92]; 
    assign layer_0[1107] = ~in[40]; 
    assign layer_0[1108] = in[69] | in[139]; 
    assign layer_0[1109] = in[90]; 
    assign layer_0[1110] = in[109] | in[91]; 
    assign layer_0[1111] = in[84] | in[76]; 
    assign layer_0[1112] = in[231] | in[228]; 
    assign layer_0[1113] = in[246] | in[249]; 
    assign layer_0[1114] = in[123]; 
    assign layer_0[1115] = in[230] | in[132]; 
    assign layer_0[1116] = in[132] | in[132]; 
    assign layer_0[1117] = ~in[105] | (in[234] & in[105]); 
    assign layer_0[1118] = in[156] ^ in[117]; 
    assign layer_0[1119] = in[91] | in[115]; 
    assign layer_0[1120] = in[92] | in[116]; 
    assign layer_0[1121] = in[51] | in[91]; 
    assign layer_0[1122] = in[230] | in[233]; 
    assign layer_0[1123] = in[92] | in[91]; 
    assign layer_0[1124] = in[109] | in[91]; 
    assign layer_0[1125] = in[108] | in[100]; 
    assign layer_0[1126] = in[156] ^ in[154]; 
    assign layer_0[1127] = in[108] | in[133]; 
    assign layer_0[1128] = in[230] | in[131]; 
    assign layer_0[1129] = in[147] | in[90]; 
    assign layer_0[1130] = in[116]; 
    assign layer_0[1131] = ~(in[233] | in[137]); 
    assign layer_0[1132] = in[90] ^ in[52]; 
    assign layer_0[1133] = in[101]; 
    assign layer_0[1134] = ~in[120] | (in[120] & in[61]); 
    assign layer_0[1135] = in[91] | in[233]; 
    assign layer_0[1136] = in[92] | in[100]; 
    assign layer_0[1137] = in[90]; 
    assign layer_0[1138] = in[93] | in[90]; 
    assign layer_0[1139] = in[75] | in[58]; 
    assign layer_0[1140] = in[90] | in[249]; 
    assign layer_0[1141] = in[115] | in[101]; 
    assign layer_0[1142] = in[101] & ~in[172]; 
    assign layer_0[1143] = in[101] | in[100]; 
    assign layer_0[1144] = in[91] | in[92]; 
    assign layer_0[1145] = in[74]; 
    assign layer_0[1146] = in[117] | in[85]; 
    assign layer_0[1147] = in[116] | in[76]; 
    assign layer_0[1148] = in[133] | in[133]; 
    assign layer_0[1149] = in[116] | in[247]; 
    assign layer_0[1150] = in[247] | in[116]; 
    assign layer_0[1151] = in[116]; 
    assign layer_0[1152] = in[90]; 
    assign layer_0[1153] = in[91]; 
    assign layer_0[1154] = in[215] & ~in[156]; 
    assign layer_0[1155] = in[156] ^ in[101]; 
    assign layer_0[1156] = in[247] | in[115]; 
    assign layer_0[1157] = in[108] | in[116]; 
    assign layer_0[1158] = in[230] | in[232]; 
    assign layer_0[1159] = in[132] | in[116]; 
    assign layer_0[1160] = in[24] | in[26]; 
    assign layer_0[1161] = ~(in[120] | in[152]); 
    assign layer_0[1162] = in[116] & ~in[22]; 
    assign layer_0[1163] = in[100] | in[75]; 
    assign layer_0[1164] = in[74] | in[75]; 
    assign layer_0[1165] = ~in[40]; 
    assign layer_0[1166] = in[248] | in[74]; 
    assign layer_0[1167] = in[92] | in[83]; 
    assign layer_0[1168] = in[100] | in[91]; 
    assign layer_0[1169] = in[116] | in[244]; 
    assign layer_0[1170] = in[53] ^ in[101]; 
    assign layer_0[1171] = ~in[182] | (in[182] & in[53]); 
    assign layer_0[1172] = in[197] & ~in[62]; 
    assign layer_0[1173] = in[116] | in[229]; 
    assign layer_0[1174] = in[108] | in[248]; 
    assign layer_0[1175] = in[116] | in[108]; 
    assign layer_0[1176] = in[101]; 
    assign layer_0[1177] = ~in[151]; 
    assign layer_0[1178] = in[116] | in[100]; 
    assign layer_0[1179] = ~in[40]; 
    assign layer_0[1180] = in[132]; 
    assign layer_0[1181] = in[74] | in[91]; 
    assign layer_0[1182] = in[117]; 
    assign layer_0[1183] = in[91] | in[68]; 
    assign layer_0[1184] = in[116]; 
    assign layer_0[1185] = in[156] ^ in[117]; 
    assign layer_0[1186] = in[92]; 
    assign layer_0[1187] = in[156] | in[218]; 
    assign layer_0[1188] = in[248] | in[116]; 
    assign layer_0[1189] = in[117] | in[83]; 
    assign layer_0[1190] = in[90] | in[92]; 
    assign layer_0[1191] = ~in[40]; 
    assign layer_0[1192] = in[90]; 
    assign layer_0[1193] = in[139] | in[26]; 
    assign layer_0[1194] = in[125] | in[108]; 
    assign layer_0[1195] = in[92] | in[101]; 
    assign layer_0[1196] = in[116]; 
    assign layer_0[1197] = in[116] | in[246]; 
    assign layer_0[1198] = in[116] | in[248]; 
    assign layer_0[1199] = in[102]; 
    assign layer_0[1200] = in[122] & ~in[156]; 
    assign layer_0[1201] = in[83] | in[90]; 
    assign layer_0[1202] = in[132] | in[92]; 
    assign layer_0[1203] = in[90]; 
    assign layer_0[1204] = in[68] ^ in[117]; 
    assign layer_0[1205] = in[116]; 
    assign layer_0[1206] = in[102]; 
    assign layer_0[1207] = in[132]; 
    assign layer_0[1208] = in[247] | in[148]; 
    assign layer_0[1209] = in[132]; 
    assign layer_0[1210] = in[90] | in[75]; 
    assign layer_0[1211] = in[92] | in[100]; 
    assign layer_0[1212] = in[90] & ~in[25]; 
    assign layer_0[1213] = in[246] | in[116]; 
    assign layer_0[1214] = in[108] | in[116]; 
    assign layer_0[1215] = in[99] & ~in[37]; 
    assign layer_0[1216] = in[230] | in[228]; 
    assign layer_0[1217] = in[117]; 
    assign layer_0[1218] = in[53] | in[163]; 
    assign layer_0[1219] = in[101]; 
    assign layer_0[1220] = in[51] | in[91]; 
    assign layer_0[1221] = in[84] ^ in[62]; 
    assign layer_0[1222] = in[91] | in[85]; 
    assign layer_0[1223] = ~in[135] | (in[135] & in[116]); 
    assign layer_0[1224] = in[132] | in[91]; 
    assign layer_0[1225] = in[107]; 
    assign layer_0[1226] = in[90] & ~in[166]; 
    assign layer_0[1227] = in[108] | in[116]; 
    assign layer_0[1228] = in[116] | in[109]; 
    assign layer_0[1229] = ~(in[166] | in[40]); 
    assign layer_0[1230] = in[68] & ~in[203]; 
    assign layer_0[1231] = ~in[41] | (in[41] & in[116]); 
    assign layer_0[1232] = in[100]; 
    assign layer_0[1233] = in[124] | in[116]; 
    assign layer_0[1234] = in[147] | in[116]; 
    assign layer_0[1235] = in[117]; 
    assign layer_0[1236] = in[246] | in[101]; 
    assign layer_0[1237] = in[123]; 
    assign layer_0[1238] = in[170] ^ in[203]; 
    assign layer_0[1239] = in[109] | in[101]; 
    assign layer_0[1240] = in[248] | in[85]; 
    assign layer_0[1241] = in[101] | in[124]; 
    assign layer_0[1242] = in[117] | in[172]; 
    assign layer_0[1243] = in[91]; 
    assign layer_0[1244] = in[131] | in[184]; 
    assign layer_0[1245] = in[91]; 
    assign layer_0[1246] = in[101] | in[247]; 
    assign layer_0[1247] = in[91]; 
    assign layer_0[1248] = in[26] | in[132]; 
    assign layer_0[1249] = in[84]; 
    assign layer_0[1250] = in[83] | in[91]; 
    assign layer_0[1251] = in[99] | in[117]; 
    assign layer_0[1252] = in[108] | in[116]; 
    assign layer_0[1253] = in[247] | in[132]; 
    assign layer_0[1254] = in[248] | in[132]; 
    assign layer_0[1255] = in[101]; 
    assign layer_0[1256] = in[132] | in[247]; 
    assign layer_0[1257] = in[91] | in[52]; 
    assign layer_0[1258] = in[90] | in[75]; 
    assign layer_0[1259] = ~in[134]; 
    assign layer_0[1260] = in[91] | in[116]; 
    assign layer_0[1261] = in[116] | in[100]; 
    assign layer_0[1262] = in[91] | in[100]; 
    assign layer_0[1263] = in[92] | in[100]; 
    assign layer_0[1264] = in[230] | in[132]; 
    assign layer_0[1265] = in[108]; 
    assign layer_0[1266] = in[247] | in[116]; 
    assign layer_0[1267] = in[61] | in[147]; 
    assign layer_0[1268] = in[92] | in[91]; 
    assign layer_0[1269] = ~in[39]; 
    assign layer_0[1270] = in[132] ^ in[245]; 
    assign layer_0[1271] = in[74] | in[91]; 
    assign layer_0[1272] = in[75] | in[100]; 
    assign layer_0[1273] = in[170] ^ in[86]; 
    assign layer_0[1274] = ~in[40]; 
    assign layer_0[1275] = in[163] | in[155]; 
    assign layer_0[1276] = ~in[151]; 
    assign layer_0[1277] = in[132] ^ in[67]; 
    assign layer_0[1278] = in[133] | in[132]; 
    assign layer_0[1279] = in[100] | in[248]; 
    assign layer_0[1280] = in[231] | in[86]; 
    assign layer_0[1281] = in[91]; 
    assign layer_0[1282] = in[116] | in[248]; 
    assign layer_0[1283] = in[109] | in[107]; 
    assign layer_0[1284] = in[73] | in[132]; 
    assign layer_0[1285] = ~in[40]; 
    assign layer_0[1286] = in[231] | in[99]; 
    assign layer_0[1287] = in[233] ^ in[230]; 
    assign layer_0[1288] = in[106]; 
    assign layer_0[1289] = in[100] | in[91]; 
    assign layer_0[1290] = ~in[166] | (in[166] & in[148]); 
    assign layer_0[1291] = in[101]; 
    assign layer_0[1292] = in[88] & ~in[180]; 
    assign layer_0[1293] = in[116]; 
    assign layer_0[1294] = in[246] | in[116]; 
    assign layer_0[1295] = in[108] | in[154]; 
    assign layer_0[1296] = in[90]; 
    assign layer_0[1297] = in[93] ^ in[90]; 
    assign layer_0[1298] = in[90] | in[93]; 
    assign layer_0[1299] = in[246] | in[115]; 
    // Layer 1 ============================================================
    assign layer_1[0] = ~layer_0[1081]; 
    assign layer_1[1] = ~layer_0[874]; 
    assign layer_1[2] = ~(layer_0[1007] & layer_0[606]); 
    assign layer_1[3] = ~layer_0[835]; 
    assign layer_1[4] = ~(layer_0[2] | layer_0[2]); 
    assign layer_1[5] = ~layer_0[785]; 
    assign layer_1[6] = ~layer_0[168]; 
    assign layer_1[7] = ~layer_0[606]; 
    assign layer_1[8] = ~layer_0[606]; 
    assign layer_1[9] = ~(layer_0[657] | layer_0[168]); 
    assign layer_1[10] = ~layer_0[1275]; 
    assign layer_1[11] = ~layer_0[731]; 
    assign layer_1[12] = ~layer_0[1172]; 
    assign layer_1[13] = ~layer_0[657]; 
    assign layer_1[14] = ~layer_0[994]; 
    assign layer_1[15] = ~layer_0[371]; 
    assign layer_1[16] = ~layer_0[939]; 
    assign layer_1[17] = ~layer_0[1084]; 
    assign layer_1[18] = ~layer_0[470]; 
    assign layer_1[19] = ~layer_0[139]; 
    assign layer_1[20] = ~layer_0[54]; 
    assign layer_1[21] = ~layer_0[1045]; 
    assign layer_1[22] = ~(layer_0[933] & layer_0[597]); 
    assign layer_1[23] = ~layer_0[855]; 
    assign layer_1[24] = ~layer_0[246]; 
    assign layer_1[25] = ~(layer_0[1046] | layer_0[326]); 
    assign layer_1[26] = ~(layer_0[0] | layer_0[1190]); 
    assign layer_1[27] = ~layer_0[52]; 
    assign layer_1[28] = ~layer_0[312]; 
    assign layer_1[29] = ~(layer_0[365] & layer_0[736]); 
    assign layer_1[30] = ~layer_0[504]; 
    assign layer_1[31] = ~layer_0[555]; 
    assign layer_1[32] = ~layer_0[630]; 
    assign layer_1[33] = ~layer_0[1084]; 
    assign layer_1[34] = ~layer_0[951]; 
    assign layer_1[35] = ~layer_0[420]; 
    assign layer_1[36] = ~layer_0[1217]; 
    assign layer_1[37] = ~layer_0[114]; 
    assign layer_1[38] = ~layer_0[1230]; 
    assign layer_1[39] = ~layer_0[943]; 
    assign layer_1[40] = ~layer_0[1062]; 
    assign layer_1[41] = ~layer_0[1154]; 
    assign layer_1[42] = ~layer_0[1149]; 
    assign layer_1[43] = ~layer_0[52]; 
    assign layer_1[44] = ~layer_0[1142]; 
    assign layer_1[45] = ~layer_0[581]; 
    assign layer_1[46] = ~layer_0[532]; 
    assign layer_1[47] = ~layer_0[283]; 
    assign layer_1[48] = ~layer_0[934]; 
    assign layer_1[49] = ~layer_0[524]; 
    assign layer_1[50] = ~(layer_0[52] & layer_0[750]); 
    assign layer_1[51] = ~layer_0[76]; 
    assign layer_1[52] = ~layer_0[470]; 
    assign layer_1[53] = ~layer_0[996]; 
    assign layer_1[54] = ~layer_0[139]; 
    assign layer_1[55] = ~layer_0[167]; 
    assign layer_1[56] = ~layer_0[691]; 
    assign layer_1[57] = ~layer_0[90]; 
    assign layer_1[58] = layer_0[1200] & ~layer_0[457]; 
    assign layer_1[59] = ~layer_0[1194]; 
    assign layer_1[60] = ~layer_0[493]; 
    assign layer_1[61] = ~layer_0[1054]; 
    assign layer_1[62] = ~layer_0[1292]; 
    assign layer_1[63] = ~layer_0[1011]; 
    assign layer_1[64] = ~(layer_0[904] | layer_0[818]); 
    assign layer_1[65] = ~layer_0[644]; 
    assign layer_1[66] = ~layer_0[1299]; 
    assign layer_1[67] = ~layer_0[1222]; 
    assign layer_1[68] = ~(layer_0[1183] | layer_0[691]); 
    assign layer_1[69] = ~layer_0[1085]; 
    assign layer_1[70] = ~layer_0[807]; 
    assign layer_1[71] = ~layer_0[943]; 
    assign layer_1[72] = ~layer_0[1134]; 
    assign layer_1[73] = ~layer_0[371]; 
    assign layer_1[74] = ~layer_0[111]; 
    assign layer_1[75] = ~layer_0[589]; 
    assign layer_1[76] = ~(layer_0[1037] | layer_0[99]); 
    assign layer_1[77] = ~layer_0[1065]; 
    assign layer_1[78] = ~layer_0[1065]; 
    assign layer_1[79] = ~layer_0[236]; 
    assign layer_1[80] = ~layer_0[652]; 
    assign layer_1[81] = ~(layer_0[114] | layer_0[444]); 
    assign layer_1[82] = ~layer_0[1007]; 
    assign layer_1[83] = ~layer_0[244]; 
    assign layer_1[84] = ~layer_0[470]; 
    assign layer_1[85] = ~(layer_0[700] & layer_0[1018]); 
    assign layer_1[86] = ~layer_0[54]; 
    assign layer_1[87] = ~layer_0[999]; 
    assign layer_1[88] = ~layer_0[1292]; 
    assign layer_1[89] = ~layer_0[581]; 
    assign layer_1[90] = ~layer_0[1143]; 
    assign layer_1[91] = ~layer_0[380]; 
    assign layer_1[92] = ~layer_0[804]; 
    assign layer_1[93] = ~layer_0[606]; 
    assign layer_1[94] = ~layer_0[994]; 
    assign layer_1[95] = ~layer_0[581]; 
    assign layer_1[96] = ~layer_0[700]; 
    assign layer_1[97] = ~layer_0[1230]; 
    assign layer_1[98] = ~layer_0[425]; 
    assign layer_1[99] = ~layer_0[1067]; 
    assign layer_1[100] = ~layer_0[573]; 
    assign layer_1[101] = ~layer_0[162]; 
    assign layer_1[102] = ~layer_0[1015]; 
    assign layer_1[103] = ~layer_0[10]; 
    assign layer_1[104] = ~layer_0[82]; 
    assign layer_1[105] = ~layer_0[681]; 
    assign layer_1[106] = ~layer_0[308]; 
    assign layer_1[107] = ~layer_0[1190]; 
    assign layer_1[108] = ~layer_0[1160]; 
    assign layer_1[109] = ~layer_0[240]; 
    assign layer_1[110] = ~(layer_0[573] | layer_0[1046]); 
    assign layer_1[111] = ~layer_0[1299]; 
    assign layer_1[112] = ~layer_0[308]; 
    assign layer_1[113] = ~layer_0[244]; 
    assign layer_1[114] = ~layer_0[208]; 
    assign layer_1[115] = ~(layer_0[162] & layer_0[1202]); 
    assign layer_1[116] = ~layer_0[855]; 
    assign layer_1[117] = ~layer_0[799]; 
    assign layer_1[118] = ~layer_0[983]; 
    assign layer_1[119] = ~layer_0[66]; 
    assign layer_1[120] = ~layer_0[167]; 
    assign layer_1[121] = ~layer_0[208]; 
    assign layer_1[122] = ~layer_0[283]; 
    assign layer_1[123] = ~layer_0[1230]; 
    assign layer_1[124] = ~layer_0[962]; 
    assign layer_1[125] = ~layer_0[1292]; 
    assign layer_1[126] = ~layer_0[200]; 
    assign layer_1[127] = ~layer_0[38]; 
    assign layer_1[128] = ~layer_0[652]; 
    assign layer_1[129] = ~layer_0[1059]; 
    assign layer_1[130] = ~layer_0[861]; 
    assign layer_1[131] = ~layer_0[573]; 
    assign layer_1[132] = ~layer_0[392]; 
    assign layer_1[133] = ~layer_0[233]; 
    assign layer_1[134] = ~layer_0[308]; 
    assign layer_1[135] = ~layer_0[398]; 
    assign layer_1[136] = ~layer_0[1202]; 
    assign layer_1[137] = ~layer_0[457]; 
    assign layer_1[138] = ~layer_0[139]; 
    assign layer_1[139] = ~(layer_0[889] & layer_0[82]); 
    assign layer_1[140] = ~layer_0[493]; 
    assign layer_1[141] = ~layer_0[1067]; 
    assign layer_1[142] = ~layer_0[685]; 
    assign layer_1[143] = ~(layer_0[398] ^ layer_0[262]); 
    assign layer_1[144] = ~layer_0[1067]; 
    assign layer_1[145] = ~(layer_0[907] | layer_0[1299]); 
    assign layer_1[146] = ~layer_0[532]; 
    assign layer_1[147] = ~layer_0[126]; 
    assign layer_1[148] = ~layer_0[890]; 
    assign layer_1[149] = ~layer_0[1045]; 
    assign layer_1[150] = ~layer_0[1054]; 
    assign layer_1[151] = ~(layer_0[76] & layer_0[1131]); 
    assign layer_1[152] = ~layer_0[501]; 
    assign layer_1[153] = ~layer_0[890]; 
    assign layer_1[154] = ~layer_0[194]; 
    assign layer_1[155] = ~layer_0[1054]; 
    assign layer_1[156] = ~layer_0[452]; 
    assign layer_1[157] = ~layer_0[139]; 
    assign layer_1[158] = ~layer_0[1287]; 
    assign layer_1[159] = ~(layer_0[283] & layer_0[606]); 
    assign layer_1[160] = ~layer_0[1299]; 
    assign layer_1[161] = ~layer_0[652]; 
    assign layer_1[162] = ~layer_0[82]; 
    assign layer_1[163] = ~layer_0[890]; 
    assign layer_1[164] = ~layer_0[469]; 
    assign layer_1[165] = ~layer_0[1088]; 
    assign layer_1[166] = ~layer_0[573]; 
    assign layer_1[167] = ~layer_0[470]; 
    assign layer_1[168] = ~layer_0[1057]; 
    assign layer_1[169] = ~layer_0[792]; 
    assign layer_1[170] = ~(layer_0[1193] | layer_0[1022]); 
    assign layer_1[171] = ~(layer_0[199] & layer_0[52]); 
    assign layer_1[172] = ~layer_0[1081]; 
    assign layer_1[173] = ~layer_0[426]; 
    assign layer_1[174] = ~layer_0[524]; 
    assign layer_1[175] = ~layer_0[365]; 
    assign layer_1[176] = ~layer_0[652]; 
    assign layer_1[177] = ~layer_0[652]; 
    assign layer_1[178] = ~layer_0[1292]; 
    assign layer_1[179] = ~layer_0[446]; 
    assign layer_1[180] = ~layer_0[1084]; 
    assign layer_1[181] = ~layer_0[460]; 
    assign layer_1[182] = ~layer_0[731]; 
    assign layer_1[183] = ~layer_0[996]; 
    assign layer_1[184] = ~layer_0[806]; 
    assign layer_1[185] = ~layer_0[1081]; 
    assign layer_1[186] = ~layer_0[1117]; 
    assign layer_1[187] = ~layer_0[1149]; 
    assign layer_1[188] = ~layer_0[581]; 
    assign layer_1[189] = ~layer_0[1237]; 
    assign layer_1[190] = ~layer_0[406]; 
    assign layer_1[191] = ~layer_0[571]; 
    assign layer_1[192] = ~layer_0[236]; 
    assign layer_1[193] = ~layer_0[606]; 
    assign layer_1[194] = ~layer_0[115]; 
    assign layer_1[195] = ~layer_0[419]; 
    assign layer_1[196] = ~(layer_0[652] | layer_0[365]); 
    assign layer_1[197] = ~layer_0[10]; 
    assign layer_1[198] = ~(layer_0[1183] | layer_0[575]); 
    assign layer_1[199] = ~layer_0[82]; 
    assign layer_1[200] = ~layer_0[652]; 
    assign layer_1[201] = ~layer_0[433]; 
    assign layer_1[202] = ~layer_0[283]; 
    assign layer_1[203] = ~layer_0[76]; 
    assign layer_1[204] = ~layer_0[457]; 
    assign layer_1[205] = ~layer_0[702]; 
    assign layer_1[206] = ~layer_0[365]; 
    assign layer_1[207] = ~layer_0[395]; 
    assign layer_1[208] = ~(layer_0[1258] & layer_0[1161]); 
    assign layer_1[209] = ~layer_0[1063]; 
    assign layer_1[210] = ~layer_0[139]; 
    assign layer_1[211] = ~layer_0[807]; 
    assign layer_1[212] = ~(layer_0[0] | layer_0[388]); 
    assign layer_1[213] = ~layer_0[1065]; 
    assign layer_1[214] = ~layer_0[493]; 
    assign layer_1[215] = ~layer_0[996]; 
    assign layer_1[216] = ~layer_0[52]; 
    assign layer_1[217] = ~layer_0[577]; 
    assign layer_1[218] = ~layer_0[1081]; 
    assign layer_1[219] = ~(layer_0[1247] | layer_0[1193]); 
    assign layer_1[220] = ~layer_0[1054]; 
    assign layer_1[221] = ~layer_0[524]; 
    assign layer_1[222] = ~layer_0[861]; 
    assign layer_1[223] = ~layer_0[1054]; 
    assign layer_1[224] = ~layer_0[581]; 
    assign layer_1[225] = ~layer_0[1081]; 
    assign layer_1[226] = ~(layer_0[1160] | layer_0[168]); 
    assign layer_1[227] = ~layer_0[736]; 
    assign layer_1[228] = ~layer_0[1183]; 
    assign layer_1[229] = ~layer_0[82]; 
    assign layer_1[230] = ~layer_0[73]; 
    assign layer_1[231] = ~layer_0[1299]; 
    assign layer_1[232] = ~layer_0[994]; 
    assign layer_1[233] = ~layer_0[581]; 
    assign layer_1[234] = ~(layer_0[917] ^ layer_0[406]); 
    assign layer_1[235] = ~layer_0[136]; 
    assign layer_1[236] = ~layer_0[202]; 
    assign layer_1[237] = ~layer_0[819]; 
    assign layer_1[238] = ~layer_0[76]; 
    assign layer_1[239] = ~layer_0[606]; 
    assign layer_1[240] = ~layer_0[691]; 
    assign layer_1[241] = ~layer_0[785]; 
    assign layer_1[242] = ~layer_0[589]; 
    assign layer_1[243] = ~layer_0[35]; 
    assign layer_1[244] = ~layer_0[52]; 
    assign layer_1[245] = ~layer_0[41]; 
    assign layer_1[246] = ~layer_0[381]; 
    assign layer_1[247] = ~layer_0[167]; 
    assign layer_1[248] = ~layer_0[1236]; 
    assign layer_1[249] = ~(layer_0[597] & layer_0[513]); 
    assign layer_1[250] = ~layer_0[470]; 
    assign layer_1[251] = ~layer_0[1099]; 
    assign layer_1[252] = ~layer_0[532]; 
    assign layer_1[253] = ~layer_0[415]; 
    assign layer_1[254] = ~(layer_0[555] | layer_0[397]); 
    assign layer_1[255] = ~layer_0[671]; 
    assign layer_1[256] = ~layer_0[597]; 
    assign layer_1[257] = ~layer_0[652]; 
    assign layer_1[258] = ~layer_0[862]; 
    assign layer_1[259] = ~layer_0[1081]; 
    assign layer_1[260] = ~layer_0[168]; 
    assign layer_1[261] = ~layer_0[470]; 
    assign layer_1[262] = ~layer_0[1165]; 
    assign layer_1[263] = ~layer_0[781]; 
    assign layer_1[264] = ~(layer_0[1249] ^ layer_0[687]); 
    assign layer_1[265] = ~layer_0[1099]; 
    assign layer_1[266] = ~layer_0[236]; 
    assign layer_1[267] = ~layer_0[657]; 
    assign layer_1[268] = ~(layer_0[1172] & layer_0[2]); 
    assign layer_1[269] = ~layer_0[139]; 
    assign layer_1[270] = ~layer_0[1081]; 
    assign layer_1[271] = ~layer_0[805]; 
    assign layer_1[272] = ~layer_0[426]; 
    assign layer_1[273] = ~layer_0[1067]; 
    assign layer_1[274] = ~layer_0[1015]; 
    assign layer_1[275] = ~layer_0[768]; 
    assign layer_1[276] = ~(layer_0[358] | layer_0[869]); 
    assign layer_1[277] = ~layer_0[785]; 
    assign layer_1[278] = ~layer_0[293]; 
    assign layer_1[279] = ~layer_0[443]; 
    assign layer_1[280] = ~layer_0[1054]; 
    assign layer_1[281] = ~layer_0[630]; 
    assign layer_1[282] = ~layer_0[41]; 
    assign layer_1[283] = ~layer_0[855]; 
    assign layer_1[284] = ~layer_0[278]; 
    assign layer_1[285] = ~layer_0[581]; 
    assign layer_1[286] = ~layer_0[167]; 
    assign layer_1[287] = ~layer_0[252]; 
    assign layer_1[288] = ~layer_0[446]; 
    assign layer_1[289] = ~(layer_0[1099] & layer_0[52]); 
    assign layer_1[290] = ~layer_0[64]; 
    assign layer_1[291] = ~layer_0[502]; 
    assign layer_1[292] = ~layer_0[1054]; 
    assign layer_1[293] = ~layer_0[10]; 
    assign layer_1[294] = ~layer_0[1299]; 
    assign layer_1[295] = ~layer_0[51]; 
    assign layer_1[296] = ~layer_0[890]; 
    assign layer_1[297] = ~layer_0[768]; 
    assign layer_1[298] = ~(layer_0[388] | layer_0[1258]); 
    assign layer_1[299] = ~layer_0[470]; 
    assign layer_1[300] = ~layer_0[1247]; 
    assign layer_1[301] = ~(layer_0[939] | layer_0[780]); 
    assign layer_1[302] = ~layer_0[371]; 
    assign layer_1[303] = ~layer_0[652]; 
    assign layer_1[304] = ~layer_0[82]; 
    assign layer_1[305] = ~layer_0[1099]; 
    assign layer_1[306] = ~layer_0[294]; 
    assign layer_1[307] = ~layer_0[934]; 
    assign layer_1[308] = ~layer_0[1292]; 
    assign layer_1[309] = ~layer_0[1172]; 
    assign layer_1[310] = ~layer_0[481]; 
    assign layer_1[311] = ~layer_0[1238]; 
    assign layer_1[312] = ~layer_0[781]; 
    assign layer_1[313] = ~layer_0[1290]; 
    assign layer_1[314] = ~layer_0[76]; 
    assign layer_1[315] = ~layer_0[82]; 
    assign layer_1[316] = ~(layer_0[781] | layer_0[379]); 
    assign layer_1[317] = ~layer_0[731]; 
    assign layer_1[318] = ~(layer_0[957] & layer_0[481]); 
    assign layer_1[319] = ~layer_0[644]; 
    assign layer_1[320] = ~layer_0[195]; 
    assign layer_1[321] = ~layer_0[373]; 
    assign layer_1[322] = ~layer_0[738]; 
    assign layer_1[323] = ~layer_0[41]; 
    assign layer_1[324] = ~layer_0[168]; 
    assign layer_1[325] = ~(layer_0[597] | layer_0[481]); 
    assign layer_1[326] = ~layer_0[855]; 
    assign layer_1[327] = ~layer_0[568]; 
    assign layer_1[328] = ~layer_0[283]; 
    assign layer_1[329] = ~layer_0[371]; 
    assign layer_1[330] = ~layer_0[1081]; 
    assign layer_1[331] = ~layer_0[1241]; 
    assign layer_1[332] = ~layer_0[64]; 
    assign layer_1[333] = ~layer_0[1190]; 
    assign layer_1[334] = ~layer_0[1007]; 
    assign layer_1[335] = ~layer_0[1018]; 
    assign layer_1[336] = ~layer_0[10]; 
    assign layer_1[337] = ~layer_0[907]; 
    assign layer_1[338] = ~layer_0[82]; 
    assign layer_1[339] = ~layer_0[1085]; 
    assign layer_1[340] = ~layer_0[1044]; 
    assign layer_1[341] = ~layer_0[1072]; 
    assign layer_1[342] = ~layer_0[194]; 
    assign layer_1[343] = ~layer_0[996]; 
    assign layer_1[344] = ~layer_0[10]; 
    assign layer_1[345] = ~layer_0[82]; 
    assign layer_1[346] = ~layer_0[555]; 
    assign layer_1[347] = ~layer_0[606]; 
    assign layer_1[348] = ~layer_0[943]; 
    assign layer_1[349] = ~layer_0[1194]; 
    assign layer_1[350] = ~layer_0[806]; 
    assign layer_1[351] = ~layer_0[691]; 
    assign layer_1[352] = ~layer_0[398]; 
    assign layer_1[353] = ~(layer_0[69] | layer_0[1170]); 
    assign layer_1[354] = ~layer_0[283]; 
    assign layer_1[355] = ~layer_0[113]; 
    assign layer_1[356] = ~layer_0[581]; 
    assign layer_1[357] = ~layer_0[1087]; 
    assign layer_1[358] = ~layer_0[934]; 
    assign layer_1[359] = ~layer_0[1007]; 
    assign layer_1[360] = ~layer_0[819]; 
    assign layer_1[361] = ~layer_0[82]; 
    assign layer_1[362] = ~layer_0[920]; 
    assign layer_1[363] = ~layer_0[835]; 
    assign layer_1[364] = ~layer_0[581]; 
    assign layer_1[365] = ~layer_0[194]; 
    assign layer_1[366] = ~layer_0[934]; 
    assign layer_1[367] = ~layer_0[1247]; 
    assign layer_1[368] = ~layer_0[1067]; 
    assign layer_1[369] = ~layer_0[899]; 
    assign layer_1[370] = ~layer_0[382]; 
    assign layer_1[371] = ~layer_0[308]; 
    assign layer_1[372] = ~layer_0[768]; 
    assign layer_1[373] = ~layer_0[581]; 
    assign layer_1[374] = ~layer_0[623]; 
    assign layer_1[375] = ~layer_0[774]; 
    assign layer_1[376] = ~layer_0[589]; 
    assign layer_1[377] = ~layer_0[524]; 
    assign layer_1[378] = ~layer_0[862]; 
    assign layer_1[379] = ~layer_0[702]; 
    assign layer_1[380] = ~layer_0[589]; 
    assign layer_1[381] = ~layer_0[1084]; 
    assign layer_1[382] = ~layer_0[82]; 
    assign layer_1[383] = ~layer_0[64]; 
    assign layer_1[384] = ~layer_0[167]; 
    assign layer_1[385] = ~(layer_0[225] & layer_0[589]); 
    assign layer_1[386] = ~layer_0[308]; 
    assign layer_1[387] = ~layer_0[141]; 
    assign layer_1[388] = ~layer_0[1299]; 
    assign layer_1[389] = ~layer_0[1183]; 
    assign layer_1[390] = ~layer_0[41]; 
    assign layer_1[391] = ~layer_0[700]; 
    assign layer_1[392] = ~layer_0[51]; 
    assign layer_1[393] = ~layer_0[934]; 
    assign layer_1[394] = ~layer_0[38]; 
    assign layer_1[395] = ~layer_0[898]; 
    assign layer_1[396] = layer_0[518] & ~layer_0[452]; 
    assign layer_1[397] = ~layer_0[731]; 
    assign layer_1[398] = ~layer_0[806]; 
    assign layer_1[399] = ~layer_0[1190]; 
    assign layer_1[400] = ~layer_0[308]; 
    assign layer_1[401] = ~(layer_0[856] ^ layer_0[1249]); 
    assign layer_1[402] = ~layer_0[691]; 
    assign layer_1[403] = ~layer_0[524]; 
    assign layer_1[404] = ~layer_0[589]; 
    assign layer_1[405] = ~layer_0[785]; 
    assign layer_1[406] = ~(layer_0[819] | layer_0[702]); 
    assign layer_1[407] = ~layer_0[855]; 
    assign layer_1[408] = ~layer_0[283]; 
    assign layer_1[409] = ~(layer_0[2] & layer_0[139]); 
    assign layer_1[410] = ~(layer_0[528] | layer_0[141]); 
    assign layer_1[411] = ~(layer_0[316] | layer_0[708]); 
    assign layer_1[412] = ~layer_0[898]; 
    assign layer_1[413] = ~layer_0[1230]; 
    assign layer_1[414] = ~layer_0[443]; 
    assign layer_1[415] = ~layer_0[388]; 
    assign layer_1[416] = ~layer_0[373]; 
    assign layer_1[417] = ~layer_0[1014]; 
    assign layer_1[418] = ~layer_0[1081]; 
    assign layer_1[419] = ~layer_0[398]; 
    assign layer_1[420] = ~(layer_0[613] & layer_0[419]); 
    assign layer_1[421] = ~layer_0[1054]; 
    assign layer_1[422] = ~layer_0[706]; 
    assign layer_1[423] = ~layer_0[581]; 
    assign layer_1[424] = ~layer_0[775]; 
    assign layer_1[425] = ~(layer_0[0] | layer_0[1183]); 
    assign layer_1[426] = ~layer_0[304]; 
    assign layer_1[427] = ~layer_0[73]; 
    assign layer_1[428] = ~layer_0[818]; 
    assign layer_1[429] = ~layer_0[589]; 
    assign layer_1[430] = ~layer_0[1183]; 
    assign layer_1[431] = ~layer_0[735]; 
    assign layer_1[432] = ~layer_0[581]; 
    assign layer_1[433] = ~layer_0[304]; 
    assign layer_1[434] = ~layer_0[168]; 
    assign layer_1[435] = ~layer_0[786]; 
    assign layer_1[436] = ~(layer_0[943] & layer_0[848]); 
    assign layer_1[437] = ~layer_0[354]; 
    assign layer_1[438] = ~(layer_0[195] ^ layer_0[1230]); 
    assign layer_1[439] = ~layer_0[571]; 
    assign layer_1[440] = ~layer_0[1087]; 
    assign layer_1[441] = ~layer_0[1045]; 
    assign layer_1[442] = ~layer_0[890]; 
    assign layer_1[443] = ~layer_0[781]; 
    assign layer_1[444] = ~layer_0[652]; 
    assign layer_1[445] = ~layer_0[819]; 
    assign layer_1[446] = ~layer_0[1200]; 
    assign layer_1[447] = ~layer_0[1230]; 
    assign layer_1[448] = ~layer_0[1113]; 
    assign layer_1[449] = ~layer_0[1099]; 
    assign layer_1[450] = ~layer_0[208]; 
    assign layer_1[451] = ~layer_0[48]; 
    assign layer_1[452] = ~layer_0[1194]; 
    assign layer_1[453] = ~layer_0[1200]; 
    assign layer_1[454] = ~layer_0[581]; 
    assign layer_1[455] = ~layer_0[579]; 
    assign layer_1[456] = ~(layer_0[652] & layer_0[781]); 
    assign layer_1[457] = ~layer_0[495]; 
    assign layer_1[458] = ~layer_0[415]; 
    assign layer_1[459] = ~layer_0[652]; 
    assign layer_1[460] = layer_0[293]; 
    assign layer_1[461] = ~layer_0[406]; 
    assign layer_1[462] = ~layer_0[1161]; 
    assign layer_1[463] = ~layer_0[731]; 
    assign layer_1[464] = ~layer_0[983]; 
    assign layer_1[465] = ~layer_0[252]; 
    assign layer_1[466] = ~(layer_0[304] & layer_0[208]); 
    assign layer_1[467] = ~layer_0[470]; 
    assign layer_1[468] = ~layer_0[64]; 
    assign layer_1[469] = ~layer_0[371]; 
    assign layer_1[470] = ~layer_0[655]; 
    assign layer_1[471] = ~layer_0[481]; 
    assign layer_1[472] = ~layer_0[167]; 
    assign layer_1[473] = ~layer_0[524]; 
    assign layer_1[474] = ~layer_0[579]; 
    assign layer_1[475] = ~layer_0[310]; 
    assign layer_1[476] = ~(layer_0[1247] | layer_0[419]); 
    assign layer_1[477] = ~layer_0[111]; 
    assign layer_1[478] = ~layer_0[114]; 
    assign layer_1[479] = ~layer_0[785]; 
    assign layer_1[480] = ~layer_0[76]; 
    assign layer_1[481] = ~layer_0[199]; 
    assign layer_1[482] = ~(layer_0[955] | layer_0[236]); 
    assign layer_1[483] = ~layer_0[781]; 
    assign layer_1[484] = ~layer_0[806]; 
    assign layer_1[485] = ~layer_0[135]; 
    assign layer_1[486] = ~layer_0[1059]; 
    assign layer_1[487] = ~layer_0[855]; 
    assign layer_1[488] = ~layer_0[41]; 
    assign layer_1[489] = ~layer_0[1030]; 
    assign layer_1[490] = ~layer_0[251]; 
    assign layer_1[491] = ~layer_0[589]; 
    assign layer_1[492] = ~layer_0[52]; 
    assign layer_1[493] = ~layer_0[168]; 
    assign layer_1[494] = ~layer_0[495]; 
    assign layer_1[495] = ~layer_0[52]; 
    assign layer_1[496] = ~layer_0[863]; 
    assign layer_1[497] = ~layer_0[1292]; 
    assign layer_1[498] = ~layer_0[283]; 
    assign layer_1[499] = ~layer_0[114]; 
    assign layer_1[500] = ~layer_0[135]; 
    assign layer_1[501] = ~layer_0[283]; 
    assign layer_1[502] = ~(layer_0[691] & layer_0[168]); 
    assign layer_1[503] = ~layer_0[82]; 
    assign layer_1[504] = ~layer_0[1085]; 
    assign layer_1[505] = ~layer_0[644]; 
    assign layer_1[506] = ~layer_0[308]; 
    assign layer_1[507] = ~layer_0[1230]; 
    assign layer_1[508] = ~layer_0[524]; 
    assign layer_1[509] = ~layer_0[855]; 
    assign layer_1[510] = ~layer_0[946]; 
    assign layer_1[511] = ~layer_0[742]; 
    assign layer_1[512] = ~layer_0[206]; 
    assign layer_1[513] = ~layer_0[199]; 
    assign layer_1[514] = ~layer_0[2]; 
    assign layer_1[515] = ~layer_0[700]; 
    assign layer_1[516] = ~layer_0[581]; 
    assign layer_1[517] = ~layer_0[862]; 
    assign layer_1[518] = ~(layer_0[283] | layer_0[1030]); 
    assign layer_1[519] = ~layer_0[446]; 
    assign layer_1[520] = ~layer_0[781]; 
    assign layer_1[521] = ~layer_0[1202]; 
    assign layer_1[522] = ~layer_0[236]; 
    assign layer_1[523] = ~layer_0[167]; 
    assign layer_1[524] = ~layer_0[308]; 
    assign layer_1[525] = ~layer_0[1007]; 
    assign layer_1[526] = ~(layer_0[460] | layer_0[0]); 
    assign layer_1[527] = ~layer_0[524]; 
    assign layer_1[528] = ~layer_0[1004]; 
    assign layer_1[529] = ~layer_0[371]; 
    assign layer_1[530] = ~layer_0[1046]; 
    assign layer_1[531] = ~layer_0[1247]; 
    assign layer_1[532] = ~(layer_0[877] | layer_0[597]); 
    assign layer_1[533] = ~layer_0[371]; 
    assign layer_1[534] = ~layer_0[934]; 
    assign layer_1[535] = ~(layer_0[946] & layer_0[41]); 
    assign layer_1[536] = ~layer_0[606]; 
    assign layer_1[537] = ~layer_0[283]; 
    assign layer_1[538] = ~layer_0[245]; 
    assign layer_1[539] = ~(layer_0[657] & layer_0[1164]); 
    assign layer_1[540] = ~layer_0[508]; 
    assign layer_1[541] = ~layer_0[704]; 
    assign layer_1[542] = ~layer_0[1014]; 
    assign layer_1[543] = ~layer_0[581]; 
    assign layer_1[544] = ~layer_0[704]; 
    assign layer_1[545] = ~layer_0[371]; 
    assign layer_1[546] = ~(layer_0[1161] | layer_0[1161]); 
    assign layer_1[547] = ~(layer_0[970] | layer_0[597]); 
    assign layer_1[548] = ~layer_0[700]; 
    assign layer_1[549] = ~layer_0[371]; 
    assign layer_1[550] = ~(layer_0[783] | layer_0[825]); 
    assign layer_1[551] = ~layer_0[639]; 
    assign layer_1[552] = ~layer_0[1026]; 
    assign layer_1[553] = 1'b1; 
    assign layer_1[554] = ~layer_0[244]; 
    assign layer_1[555] = ~layer_0[546]; 
    assign layer_1[556] = ~layer_0[139]; 
    assign layer_1[557] = ~layer_0[457]; 
    assign layer_1[558] = ~layer_0[805]; 
    assign layer_1[559] = ~layer_0[657]; 
    assign layer_1[560] = ~layer_0[54]; 
    assign layer_1[561] = ~layer_0[76]; 
    assign layer_1[562] = ~layer_0[446]; 
    assign layer_1[563] = ~layer_0[82]; 
    assign layer_1[564] = ~layer_0[785]; 
    assign layer_1[565] = ~(layer_0[225] | layer_0[1111]); 
    assign layer_1[566] = ~layer_0[371]; 
    assign layer_1[567] = ~layer_0[798]; 
    assign layer_1[568] = ~layer_0[910]; 
    assign layer_1[569] = ~layer_0[572]; 
    assign layer_1[570] = ~layer_0[652]; 
    assign layer_1[571] = ~layer_0[354]; 
    assign layer_1[572] = ~layer_0[1275]; 
    assign layer_1[573] = ~layer_0[1067]; 
    assign layer_1[574] = ~layer_0[1085]; 
    assign layer_1[575] = ~layer_0[1183]; 
    assign layer_1[576] = ~layer_0[731]; 
    assign layer_1[577] = ~layer_0[371]; 
    assign layer_1[578] = ~layer_0[967]; 
    assign layer_1[579] = ~layer_0[934]; 
    assign layer_1[580] = ~layer_0[855]; 
    assign layer_1[581] = ~(layer_0[1187] | layer_0[882]); 
    assign layer_1[582] = ~layer_0[806]; 
    assign layer_1[583] = ~layer_0[581]; 
    assign layer_1[584] = ~layer_0[478]; 
    assign layer_1[585] = ~layer_0[528]; 
    assign layer_1[586] = ~(layer_0[190] | layer_0[722]); 
    assign layer_1[587] = ~layer_0[657]; 
    assign layer_1[588] = ~layer_0[446]; 
    assign layer_1[589] = ~layer_0[943]; 
    assign layer_1[590] = ~layer_0[1290]; 
    assign layer_1[591] = ~layer_0[597]; 
    assign layer_1[592] = ~layer_0[700]; 
    assign layer_1[593] = ~layer_0[200]; 
    assign layer_1[594] = ~layer_0[807]; 
    assign layer_1[595] = ~layer_0[231]; 
    assign layer_1[596] = ~layer_0[2]; 
    assign layer_1[597] = ~layer_0[731]; 
    assign layer_1[598] = ~(layer_0[52] & layer_0[731]); 
    assign layer_1[599] = ~layer_0[657]; 
    assign layer_1[600] = ~layer_0[1270]; 
    assign layer_1[601] = ~layer_0[371]; 
    assign layer_1[602] = ~(layer_0[227] | layer_0[1067]); 
    assign layer_1[603] = ~layer_0[502]; 
    assign layer_1[604] = ~layer_0[1081]; 
    assign layer_1[605] = ~layer_0[371]; 
    assign layer_1[606] = ~layer_0[308]; 
    assign layer_1[607] = ~layer_0[1247]; 
    assign layer_1[608] = ~layer_0[460]; 
    assign layer_1[609] = ~(layer_0[388] | layer_0[481]); 
    assign layer_1[610] = ~layer_0[861]; 
    assign layer_1[611] = ~layer_0[606]; 
    assign layer_1[612] = ~layer_0[630]; 
    assign layer_1[613] = ~layer_0[906]; 
    assign layer_1[614] = ~layer_0[606]; 
    assign layer_1[615] = ~layer_0[283]; 
    assign layer_1[616] = ~layer_0[890]; 
    assign layer_1[617] = ~layer_0[959]; 
    assign layer_1[618] = ~(layer_0[1007] | layer_0[225]); 
    assign layer_1[619] = ~layer_0[1007]; 
    assign layer_1[620] = ~layer_0[691]; 
    assign layer_1[621] = ~layer_0[606]; 
    assign layer_1[622] = ~layer_0[785]; 
    assign layer_1[623] = ~layer_0[606]; 
    assign layer_1[624] = ~layer_0[774]; 
    assign layer_1[625] = ~layer_0[832]; 
    assign layer_1[626] = ~layer_0[326]; 
    assign layer_1[627] = ~layer_0[200]; 
    assign layer_1[628] = ~layer_0[943]; 
    assign layer_1[629] = ~layer_0[1045]; 
    assign layer_1[630] = ~layer_0[774]; 
    assign layer_1[631] = ~layer_0[280]; 
    assign layer_1[632] = ~layer_0[818]; 
    assign layer_1[633] = ~layer_0[532]; 
    assign layer_1[634] = ~layer_0[704]; 
    assign layer_1[635] = ~layer_0[700]; 
    assign layer_1[636] = ~layer_0[375]; 
    assign layer_1[637] = ~layer_0[308]; 
    assign layer_1[638] = ~layer_0[1099]; 
    assign layer_1[639] = ~layer_0[855]; 
    assign layer_1[640] = ~layer_0[338]; 
    assign layer_1[641] = ~(layer_0[735] | layer_0[433]); 
    assign layer_1[642] = ~layer_0[54]; 
    assign layer_1[643] = ~layer_0[167]; 
    assign layer_1[644] = ~layer_0[781]; 
    assign layer_1[645] = ~layer_0[446]; 
    assign layer_1[646] = ~layer_0[1292]; 
    assign layer_1[647] = ~layer_0[6]; 
    assign layer_1[648] = ~(layer_0[1292] ^ layer_0[415]); 
    assign layer_1[649] = ~layer_0[501]; 
    assign layer_1[650] = ~layer_0[606]; 
    assign layer_1[651] = ~layer_0[861]; 
    assign layer_1[652] = ~layer_0[395]; 
    assign layer_1[653] = ~(layer_0[887] | layer_0[199]); 
    assign layer_1[654] = ~layer_0[113]; 
    assign layer_1[655] = ~(layer_0[202] | layer_0[1183]); 
    assign layer_1[656] = ~layer_0[581]; 
    assign layer_1[657] = ~layer_0[996]; 
    assign layer_1[658] = ~layer_0[524]; 
    assign layer_1[659] = ~layer_0[652]; 
    assign layer_1[660] = ~layer_0[652]; 
    assign layer_1[661] = ~layer_0[996]; 
    assign layer_1[662] = ~layer_0[861]; 
    assign layer_1[663] = ~layer_0[231]; 
    assign layer_1[664] = ~layer_0[1299]; 
    assign layer_1[665] = ~layer_0[443]; 
    assign layer_1[666] = ~layer_0[1247]; 
    assign layer_1[667] = ~layer_0[212]; 
    assign layer_1[668] = ~layer_0[446]; 
    assign layer_1[669] = ~layer_0[314]; 
    assign layer_1[670] = ~(layer_0[1297] & layer_0[168]); 
    assign layer_1[671] = ~layer_0[219]; 
    assign layer_1[672] = ~layer_0[589]; 
    assign layer_1[673] = ~layer_0[1099]; 
    assign layer_1[674] = ~layer_0[1190]; 
    assign layer_1[675] = ~layer_0[1113]; 
    assign layer_1[676] = ~layer_0[994]; 
    assign layer_1[677] = ~layer_0[700]; 
    assign layer_1[678] = ~layer_0[236]; 
    assign layer_1[679] = ~layer_0[64]; 
    assign layer_1[680] = ~layer_0[1190]; 
    assign layer_1[681] = ~layer_0[1099]; 
    assign layer_1[682] = ~layer_0[1194]; 
    assign layer_1[683] = ~layer_0[1292]; 
    assign layer_1[684] = ~layer_0[1125]; 
    assign layer_1[685] = ~(layer_0[168] & layer_0[881]); 
    assign layer_1[686] = ~layer_0[502]; 
    assign layer_1[687] = ~layer_0[1161]; 
    assign layer_1[688] = ~layer_0[1299]; 
    assign layer_1[689] = ~layer_0[1099]; 
    assign layer_1[690] = ~layer_0[381]; 
    assign layer_1[691] = ~layer_0[1067]; 
    assign layer_1[692] = ~layer_0[76]; 
    assign layer_1[693] = ~layer_0[457]; 
    assign layer_1[694] = ~layer_0[167]; 
    assign layer_1[695] = ~layer_0[111]; 
    assign layer_1[696] = ~layer_0[252]; 
    assign layer_1[697] = ~(layer_0[431] | layer_0[532]); 
    assign layer_1[698] = ~layer_0[541]; 
    assign layer_1[699] = ~layer_0[639]; 
    assign layer_1[700] = ~(layer_0[518] ^ layer_0[981]); 
    assign layer_1[701] = ~layer_0[657]; 
    assign layer_1[702] = ~layer_0[167]; 
    assign layer_1[703] = ~layer_0[555]; 
    assign layer_1[704] = ~layer_0[573]; 
    assign layer_1[705] = ~layer_0[283]; 
    assign layer_1[706] = ~layer_0[898]; 
    assign layer_1[707] = ~layer_0[691]; 
    assign layer_1[708] = ~(layer_0[818] & layer_0[338]); 
    assign layer_1[709] = ~layer_0[76]; 
    assign layer_1[710] = ~layer_0[962]; 
    assign layer_1[711] = ~(layer_0[760] | layer_0[1063]); 
    assign layer_1[712] = ~layer_0[785]; 
    assign layer_1[713] = ~layer_0[700]; 
    assign layer_1[714] = ~layer_0[996]; 
    assign layer_1[715] = ~layer_0[141]; 
    assign layer_1[716] = ~(layer_0[1171] | layer_0[1190]); 
    assign layer_1[717] = ~layer_0[371]; 
    assign layer_1[718] = ~(layer_0[1184] & layer_0[650]); 
    assign layer_1[719] = ~layer_0[589]; 
    assign layer_1[720] = ~layer_0[1087]; 
    assign layer_1[721] = ~(layer_0[154] | layer_0[1125]); 
    assign layer_1[722] = ~layer_0[178]; 
    assign layer_1[723] = ~layer_0[775]; 
    assign layer_1[724] = ~layer_0[1054]; 
    assign layer_1[725] = ~layer_0[76]; 
    assign layer_1[726] = ~layer_0[314]; 
    assign layer_1[727] = layer_0[330]; 
    assign layer_1[728] = ~layer_0[194]; 
    assign layer_1[729] = ~layer_0[354]; 
    assign layer_1[730] = ~layer_0[82]; 
    assign layer_1[731] = ~layer_0[446]; 
    assign layer_1[732] = ~layer_0[1059]; 
    assign layer_1[733] = ~layer_0[502]; 
    assign layer_1[734] = ~layer_0[433]; 
    assign layer_1[735] = ~layer_0[187]; 
    assign layer_1[736] = ~layer_0[819]; 
    assign layer_1[737] = ~layer_0[606]; 
    assign layer_1[738] = ~layer_0[111]; 
    assign layer_1[739] = ~layer_0[1063]; 
    assign layer_1[740] = ~layer_0[1195]; 
    assign layer_1[741] = ~layer_0[415]; 
    assign layer_1[742] = ~layer_0[768]; 
    assign layer_1[743] = ~layer_0[657]; 
    assign layer_1[744] = ~layer_0[76]; 
    assign layer_1[745] = ~layer_0[1287]; 
    assign layer_1[746] = ~layer_0[293]; 
    assign layer_1[747] = ~(layer_0[552] | layer_0[955]); 
    assign layer_1[748] = ~layer_0[863]; 
    assign layer_1[749] = ~layer_0[806]; 
    assign layer_1[750] = ~layer_0[381]; 
    assign layer_1[751] = ~layer_0[371]; 
    assign layer_1[752] = ~layer_0[76]; 
    assign layer_1[753] = ~layer_0[443]; 
    assign layer_1[754] = ~layer_0[855]; 
    assign layer_1[755] = ~layer_0[807]; 
    assign layer_1[756] = ~layer_0[959]; 
    assign layer_1[757] = ~layer_0[606]; 
    assign layer_1[758] = ~(layer_0[1275] | layer_0[870]); 
    assign layer_1[759] = ~layer_0[639]; 
    assign layer_1[760] = ~layer_0[785]; 
    assign layer_1[761] = ~(layer_0[682] & layer_0[956]); 
    assign layer_1[762] = ~layer_0[200]; 
    assign layer_1[763] = ~layer_0[657]; 
    assign layer_1[764] = ~layer_0[76]; 
    assign layer_1[765] = ~layer_0[1099]; 
    assign layer_1[766] = ~layer_0[236]; 
    assign layer_1[767] = ~layer_0[250]; 
    assign layer_1[768] = ~layer_0[1226]; 
    assign layer_1[769] = 1'b1; 
    assign layer_1[770] = ~layer_0[1244]; 
    assign layer_1[771] = ~layer_0[589]; 
    assign layer_1[772] = ~layer_0[1149]; 
    assign layer_1[773] = ~layer_0[308]; 
    assign layer_1[774] = ~layer_0[113]; 
    assign layer_1[775] = ~layer_0[1085]; 
    assign layer_1[776] = ~layer_0[244]; 
    assign layer_1[777] = ~layer_0[212]; 
    assign layer_1[778] = ~layer_0[573]; 
    assign layer_1[779] = ~(layer_0[657] | layer_0[1049]); 
    assign layer_1[780] = ~layer_0[777]; 
    assign layer_1[781] = ~layer_0[354]; 
    assign layer_1[782] = ~layer_0[656]; 
    assign layer_1[783] = ~layer_0[606]; 
    assign layer_1[784] = ~layer_0[731]; 
    assign layer_1[785] = ~(layer_0[890] | layer_0[652]); 
    assign layer_1[786] = ~layer_0[807]; 
    assign layer_1[787] = ~layer_0[240]; 
    assign layer_1[788] = ~layer_0[41]; 
    assign layer_1[789] = ~layer_0[783]; 
    assign layer_1[790] = ~(layer_0[644] | layer_0[630]); 
    assign layer_1[791] = ~layer_0[82]; 
    assign layer_1[792] = ~layer_0[167]; 
    assign layer_1[793] = layer_0[318] ^ layer_0[1190]; 
    assign layer_1[794] = ~layer_0[1046]; 
    assign layer_1[795] = ~layer_0[581]; 
    assign layer_1[796] = ~layer_0[1007]; 
    assign layer_1[797] = ~layer_0[589]; 
    assign layer_1[798] = ~(layer_0[1183] | layer_0[691]); 
    assign layer_1[799] = ~layer_0[236]; 
    assign layer_1[800] = ~layer_0[652]; 
    assign layer_1[801] = ~layer_0[82]; 
    assign layer_1[802] = ~(layer_0[139] & layer_0[972]); 
    assign layer_1[803] = ~layer_0[996]; 
    assign layer_1[804] = ~layer_0[652]; 
    assign layer_1[805] = ~layer_0[524]; 
    assign layer_1[806] = ~layer_0[691]; 
    assign layer_1[807] = ~layer_0[215]; 
    assign layer_1[808] = ~layer_0[740]; 
    assign layer_1[809] = ~layer_0[898]; 
    assign layer_1[810] = ~(layer_0[1044] & layer_0[690]); 
    assign layer_1[811] = ~layer_0[939]; 
    assign layer_1[812] = ~layer_0[1022]; 
    assign layer_1[813] = ~(layer_0[77] | layer_0[452]); 
    assign layer_1[814] = ~(layer_0[956] & layer_0[1110]); 
    assign layer_1[815] = ~layer_0[823]; 
    assign layer_1[816] = ~layer_0[1087]; 
    assign layer_1[817] = ~layer_0[345]; 
    assign layer_1[818] = ~layer_0[807]; 
    assign layer_1[819] = ~layer_0[948]; 
    assign layer_1[820] = ~layer_0[168]; 
    assign layer_1[821] = ~layer_0[1067]; 
    assign layer_1[822] = ~(layer_0[506] | layer_0[499]); 
    assign layer_1[823] = ~layer_0[365]; 
    assign layer_1[824] = ~layer_0[206]; 
    assign layer_1[825] = ~layer_0[644]; 
    assign layer_1[826] = ~layer_0[1054]; 
    assign layer_1[827] = ~layer_0[806]; 
    assign layer_1[828] = ~(layer_0[575] | layer_0[388]); 
    assign layer_1[829] = ~layer_0[644]; 
    assign layer_1[830] = ~(layer_0[597] | layer_0[1247]); 
    assign layer_1[831] = ~layer_0[874]; 
    assign layer_1[832] = ~layer_0[283]; 
    assign layer_1[833] = ~layer_0[579]; 
    assign layer_1[834] = ~layer_0[499]; 
    assign layer_1[835] = ~layer_0[1054]; 
    assign layer_1[836] = ~layer_0[630]; 
    assign layer_1[837] = ~(layer_0[10] & layer_0[898]); 
    assign layer_1[838] = ~layer_0[652]; 
    assign layer_1[839] = ~layer_0[1067]; 
    assign layer_1[840] = ~layer_0[1085]; 
    assign layer_1[841] = ~layer_0[6]; 
    assign layer_1[842] = ~layer_0[82]; 
    assign layer_1[843] = ~layer_0[1218]; 
    assign layer_1[844] = ~(layer_0[869] | layer_0[1284]); 
    assign layer_1[845] = ~layer_0[606]; 
    assign layer_1[846] = ~layer_0[606]; 
    assign layer_1[847] = ~(layer_0[1222] | layer_0[69]); 
    assign layer_1[848] = ~layer_0[1015]; 
    assign layer_1[849] = ~layer_0[194]; 
    assign layer_1[850] = ~layer_0[1247]; 
    assign layer_1[851] = ~layer_0[738]; 
    assign layer_1[852] = ~(layer_0[691] & layer_0[168]); 
    assign layer_1[853] = ~layer_0[700]; 
    assign layer_1[854] = ~layer_0[1108]; 
    assign layer_1[855] = ~layer_0[581]; 
    assign layer_1[856] = ~layer_0[1194]; 
    assign layer_1[857] = ~layer_0[1154]; 
    assign layer_1[858] = ~(layer_0[1267] | layer_0[1244]); 
    assign layer_1[859] = ~layer_0[606]; 
    assign layer_1[860] = ~layer_0[524]; 
    assign layer_1[861] = ~layer_0[835]; 
    assign layer_1[862] = ~layer_0[970]; 
    assign layer_1[863] = ~(layer_0[433] | layer_0[1267]); 
    assign layer_1[864] = ~layer_0[199]; 
    assign layer_1[865] = ~layer_0[1099]; 
    assign layer_1[866] = ~(layer_0[388] | layer_0[681]); 
    assign layer_1[867] = ~layer_0[252]; 
    assign layer_1[868] = ~layer_0[1299]; 
    assign layer_1[869] = ~layer_0[714]; 
    assign layer_1[870] = ~layer_0[202]; 
    assign layer_1[871] = ~layer_0[354]; 
    assign layer_1[872] = ~layer_0[819]; 
    assign layer_1[873] = ~(layer_0[82] & layer_0[131]); 
    assign layer_1[874] = ~(layer_0[1183] | layer_0[1190]); 
    assign layer_1[875] = ~(layer_0[1170] | layer_0[69]); 
    assign layer_1[876] = ~layer_0[1299]; 
    assign layer_1[877] = ~layer_0[1112]; 
    assign layer_1[878] = ~layer_0[606]; 
    assign layer_1[879] = ~(layer_0[314] | layer_0[589]); 
    assign layer_1[880] = ~layer_0[1149]; 
    assign layer_1[881] = ~layer_0[1212]; 
    assign layer_1[882] = ~layer_0[1099]; 
    assign layer_1[883] = ~layer_0[1267]; 
    assign layer_1[884] = ~layer_0[1149]; 
    assign layer_1[885] = ~layer_0[581]; 
    assign layer_1[886] = ~(layer_0[52] & layer_0[597]); 
    assign layer_1[887] = ~(layer_0[751] & layer_0[706]); 
    assign layer_1[888] = ~layer_0[236]; 
    assign layer_1[889] = ~layer_0[392]; 
    assign layer_1[890] = ~layer_0[967]; 
    assign layer_1[891] = ~layer_0[1030]; 
    assign layer_1[892] = ~layer_0[1087]; 
    assign layer_1[893] = ~layer_0[168]; 
    assign layer_1[894] = ~layer_0[443]; 
    assign layer_1[895] = ~layer_0[141]; 
    assign layer_1[896] = ~layer_0[1099]; 
    assign layer_1[897] = ~(layer_0[700] & layer_0[1048]); 
    assign layer_1[898] = ~layer_0[64]; 
    assign layer_1[899] = ~layer_0[681]; 
    assign layer_1[900] = ~layer_0[781]; 
    assign layer_1[901] = ~layer_0[236]; 
    assign layer_1[902] = ~layer_0[1045]; 
    assign layer_1[903] = ~layer_0[1015]; 
    assign layer_1[904] = ~(layer_0[943] & layer_0[863]); 
    assign layer_1[905] = ~layer_0[786]; 
    assign layer_1[906] = ~layer_0[1125]; 
    assign layer_1[907] = ~layer_0[1085]; 
    assign layer_1[908] = ~layer_0[806]; 
    assign layer_1[909] = ~layer_0[606]; 
    assign layer_1[910] = ~layer_0[314]; 
    assign layer_1[911] = ~layer_0[1241]; 
    assign layer_1[912] = ~layer_0[855]; 
    assign layer_1[913] = ~layer_0[740]; 
    assign layer_1[914] = ~layer_0[446]; 
    assign layer_1[915] = ~layer_0[581]; 
    assign layer_1[916] = ~layer_0[589]; 
    assign layer_1[917] = ~(layer_0[1046] | layer_0[35]); 
    assign layer_1[918] = ~layer_0[392]; 
    assign layer_1[919] = ~layer_0[353]; 
    assign layer_1[920] = ~layer_0[907]; 
    assign layer_1[921] = ~layer_0[1259]; 
    assign layer_1[922] = ~layer_0[147]; 
    assign layer_1[923] = ~(layer_0[1079] | layer_0[597]); 
    assign layer_1[924] = ~layer_0[82]; 
    assign layer_1[925] = ~layer_0[283]; 
    assign layer_1[926] = ~layer_0[1299]; 
    assign layer_1[927] = ~layer_0[543]; 
    assign layer_1[928] = ~layer_0[694]; 
    assign layer_1[929] = ~layer_0[898]; 
    assign layer_1[930] = ~layer_0[652]; 
    assign layer_1[931] = ~(layer_0[87] | layer_0[612]); 
    assign layer_1[932] = ~layer_0[1085]; 
    assign layer_1[933] = ~layer_0[406]; 
    assign layer_1[934] = ~layer_0[943]; 
    assign layer_1[935] = ~layer_0[1081]; 
    assign layer_1[936] = ~layer_0[1238]; 
    assign layer_1[937] = ~(layer_0[747] | layer_0[555]); 
    assign layer_1[938] = ~layer_0[656]; 
    assign layer_1[939] = ~layer_0[565]; 
    assign layer_1[940] = ~layer_0[219]; 
    assign layer_1[941] = ~layer_0[597]; 
    assign layer_1[942] = ~layer_0[415]; 
    assign layer_1[943] = ~(layer_0[1015] & layer_0[1292]); 
    assign layer_1[944] = ~(layer_0[910] & layer_0[972]); 
    assign layer_1[945] = ~layer_0[1287]; 
    assign layer_1[946] = ~layer_0[308]; 
    assign layer_1[947] = ~layer_0[1190]; 
    assign layer_1[948] = ~layer_0[606]; 
    assign layer_1[949] = ~layer_0[167]; 
    assign layer_1[950] = ~layer_0[426]; 
    assign layer_1[951] = ~layer_0[236]; 
    assign layer_1[952] = ~layer_0[1113]; 
    assign layer_1[953] = ~layer_0[874]; 
    assign layer_1[954] = ~layer_0[996]; 
    assign layer_1[955] = ~(layer_0[1087] & layer_0[694]); 
    assign layer_1[956] = ~layer_0[861]; 
    assign layer_1[957] = ~layer_0[446]; 
    assign layer_1[958] = ~layer_0[970]; 
    assign layer_1[959] = ~layer_0[1194]; 
    assign layer_1[960] = ~layer_0[51]; 
    assign layer_1[961] = ~layer_0[1212]; 
    assign layer_1[962] = ~layer_0[589]; 
    assign layer_1[963] = ~layer_0[1149]; 
    assign layer_1[964] = ~layer_0[851]; 
    assign layer_1[965] = ~layer_0[375]; 
    assign layer_1[966] = ~layer_0[1267]; 
    assign layer_1[967] = ~layer_0[113]; 
    assign layer_1[968] = ~layer_0[371]; 
    assign layer_1[969] = ~(layer_0[38] & layer_0[168]); 
    assign layer_1[970] = ~layer_0[856]; 
    assign layer_1[971] = ~layer_0[1081]; 
    assign layer_1[972] = ~layer_0[682]; 
    assign layer_1[973] = ~(layer_0[1004] ^ layer_0[941]); 
    assign layer_1[974] = ~layer_0[1230]; 
    assign layer_1[975] = ~(layer_0[254] & layer_0[962]); 
    assign layer_1[976] = ~layer_0[1142]; 
    assign layer_1[977] = ~layer_0[1193]; 
    assign layer_1[978] = ~layer_0[700]; 
    assign layer_1[979] = ~layer_0[415]; 
    assign layer_1[980] = ~layer_0[113]; 
    assign layer_1[981] = ~layer_0[308]; 
    assign layer_1[982] = ~layer_0[691]; 
    assign layer_1[983] = ~layer_0[768]; 
    assign layer_1[984] = ~layer_0[861]; 
    assign layer_1[985] = ~layer_0[606]; 
    assign layer_1[986] = ~layer_0[606]; 
    assign layer_1[987] = ~layer_0[652]; 
    assign layer_1[988] = ~layer_0[446]; 
    assign layer_1[989] = ~layer_0[639]; 
    assign layer_1[990] = ~layer_0[845]; 
    assign layer_1[991] = ~layer_0[460]; 
    assign layer_1[992] = ~layer_0[2]; 
    assign layer_1[993] = ~layer_0[606]; 
    assign layer_1[994] = ~layer_0[314]; 
    assign layer_1[995] = ~layer_0[139]; 
    assign layer_1[996] = ~layer_0[457]; 
    assign layer_1[997] = ~(layer_0[1183] | layer_0[202]); 
    assign layer_1[998] = ~layer_0[167]; 
    assign layer_1[999] = ~layer_0[682]; 
    assign layer_1[1000] = ~layer_0[126]; 
    assign layer_1[1001] = ~layer_0[835]; 
    assign layer_1[1002] = ~layer_0[314]; 
    assign layer_1[1003] = ~layer_0[999]; 
    assign layer_1[1004] = ~layer_0[76]; 
    assign layer_1[1005] = ~layer_0[90]; 
    assign layer_1[1006] = ~layer_0[731]; 
    assign layer_1[1007] = ~layer_0[996]; 
    assign layer_1[1008] = ~layer_0[1292]; 
    assign layer_1[1009] = ~layer_0[139]; 
    assign layer_1[1010] = ~layer_0[1247]; 
    assign layer_1[1011] = ~(layer_0[1049] | layer_0[1278]); 
    assign layer_1[1012] = ~layer_0[652]; 
    assign layer_1[1013] = ~layer_0[139]; 
    assign layer_1[1014] = ~layer_0[652]; 
    assign layer_1[1015] = ~layer_0[82]; 
    assign layer_1[1016] = ~layer_0[1063]; 
    assign layer_1[1017] = ~layer_0[1226]; 
    assign layer_1[1018] = ~layer_0[1190]; 
    assign layer_1[1019] = ~(layer_0[783] | layer_0[504]); 
    assign layer_1[1020] = ~layer_0[398]; 
    assign layer_1[1021] = ~layer_0[1267]; 
    assign layer_1[1022] = ~layer_0[691]; 
    assign layer_1[1023] = ~layer_0[855]; 
    assign layer_1[1024] = ~layer_0[10]; 
    assign layer_1[1025] = ~layer_0[946]; 
    assign layer_1[1026] = ~layer_0[1154]; 
    assign layer_1[1027] = ~layer_0[139]; 
    assign layer_1[1028] = ~layer_0[1007]; 
    assign layer_1[1029] = ~(layer_0[1172] | layer_0[433]); 
    assign layer_1[1030] = ~layer_0[82]; 
    assign layer_1[1031] = ~layer_0[1055]; 
    assign layer_1[1032] = ~layer_0[799]; 
    assign layer_1[1033] = ~layer_0[996]; 
    assign layer_1[1034] = ~layer_0[644]; 
    assign layer_1[1035] = ~layer_0[1229]; 
    assign layer_1[1036] = ~layer_0[1292]; 
    assign layer_1[1037] = ~layer_0[1045]; 
    assign layer_1[1038] = ~layer_0[1081]; 
    assign layer_1[1039] = ~layer_0[400]; 
    assign layer_1[1040] = ~(layer_0[1183] | layer_0[589]); 
    assign layer_1[1041] = ~layer_0[943]; 
    assign layer_1[1042] = ~layer_0[943]; 
    assign layer_1[1043] = ~layer_0[54]; 
    assign layer_1[1044] = ~layer_0[1081]; 
    assign layer_1[1045] = ~layer_0[1084]; 
    assign layer_1[1046] = ~layer_0[1238]; 
    assign layer_1[1047] = ~layer_0[194]; 
    assign layer_1[1048] = ~layer_0[398]; 
    assign layer_1[1049] = ~layer_0[198]; 
    assign layer_1[1050] = ~layer_0[446]; 
    assign layer_1[1051] = ~layer_0[781]; 
    assign layer_1[1052] = ~layer_0[219]; 
    assign layer_1[1053] = ~layer_0[1054]; 
    assign layer_1[1054] = ~layer_0[1022]; 
    assign layer_1[1055] = ~layer_0[139]; 
    assign layer_1[1056] = ~layer_0[1194]; 
    assign layer_1[1057] = ~layer_0[571]; 
    assign layer_1[1058] = ~layer_0[691]; 
    assign layer_1[1059] = ~layer_0[371]; 
    assign layer_1[1060] = layer_0[997] & ~layer_0[934]; 
    assign layer_1[1061] = ~layer_0[82]; 
    assign layer_1[1062] = ~layer_0[644]; 
    assign layer_1[1063] = ~(layer_0[250] | layer_0[1046]); 
    assign layer_1[1064] = ~layer_0[114]; 
    assign layer_1[1065] = layer_0[1127] & ~layer_0[835]; 
    assign layer_1[1066] = ~layer_0[1237]; 
    assign layer_1[1067] = ~layer_0[907]; 
    assign layer_1[1068] = ~layer_0[658]; 
    assign layer_1[1069] = ~layer_0[90]; 
    assign layer_1[1070] = ~layer_0[786]; 
    assign layer_1[1071] = ~(layer_0[613] | layer_0[1139]); 
    assign layer_1[1072] = ~layer_0[82]; 
    assign layer_1[1073] = ~(layer_0[1275] | layer_0[868]); 
    assign layer_1[1074] = ~(layer_0[1171] | layer_0[691]); 
    assign layer_1[1075] = ~layer_0[606]; 
    assign layer_1[1076] = ~layer_0[1183]; 
    assign layer_1[1077] = ~layer_0[524]; 
    assign layer_1[1078] = ~layer_0[139]; 
    assign layer_1[1079] = ~layer_0[82]; 
    assign layer_1[1080] = ~layer_0[947]; 
    assign layer_1[1081] = ~layer_0[415]; 
    assign layer_1[1082] = ~layer_0[1067]; 
    assign layer_1[1083] = ~layer_0[1299]; 
    assign layer_1[1084] = ~layer_0[781]; 
    assign layer_1[1085] = ~layer_0[236]; 
    assign layer_1[1086] = ~layer_0[1299]; 
    assign layer_1[1087] = ~layer_0[1085]; 
    assign layer_1[1088] = ~layer_0[731]; 
    assign layer_1[1089] = ~layer_0[785]; 
    assign layer_1[1090] = ~layer_0[345]; 
    assign layer_1[1091] = ~layer_0[972]; 
    assign layer_1[1092] = ~layer_0[691]; 
    assign layer_1[1093] = ~layer_0[907]; 
    assign layer_1[1094] = ~layer_0[1190]; 
    assign layer_1[1095] = ~layer_0[656]; 
    assign layer_1[1096] = ~layer_0[1292]; 
    assign layer_1[1097] = ~layer_0[644]; 
    assign layer_1[1098] = ~layer_0[499]; 
    assign layer_1[1099] = ~layer_0[806]; 
    assign layer_1[1100] = ~layer_0[1299]; 
    assign layer_1[1101] = ~layer_0[652]; 
    assign layer_1[1102] = ~layer_0[406]; 
    assign layer_1[1103] = ~(layer_0[1015] & layer_0[485]); 
    assign layer_1[1104] = ~layer_0[524]; 
    assign layer_1[1105] = ~(layer_0[774] & layer_0[804]); 
    assign layer_1[1106] = ~layer_0[426]; 
    assign layer_1[1107] = ~layer_0[581]; 
    assign layer_1[1108] = ~layer_0[1081]; 
    assign layer_1[1109] = ~layer_0[390]; 
    assign layer_1[1110] = ~layer_0[898]; 
    assign layer_1[1111] = ~layer_0[113]; 
    assign layer_1[1112] = ~layer_0[1081]; 
    assign layer_1[1113] = ~layer_0[1054]; 
    assign layer_1[1114] = ~layer_0[395]; 
    assign layer_1[1115] = ~layer_0[934]; 
    assign layer_1[1116] = ~layer_0[308]; 
    assign layer_1[1117] = ~layer_0[785]; 
    assign layer_1[1118] = ~layer_0[835]; 
    assign layer_1[1119] = ~layer_0[874]; 
    assign layer_1[1120] = ~layer_0[687]; 
    assign layer_1[1121] = ~layer_0[1134]; 
    assign layer_1[1122] = ~layer_0[1297]; 
    assign layer_1[1123] = ~layer_0[1292]; 
    assign layer_1[1124] = ~layer_0[1125]; 
    assign layer_1[1125] = ~layer_0[818]; 
    assign layer_1[1126] = ~layer_0[65]; 
    assign layer_1[1127] = ~(layer_0[113] | layer_0[1046]); 
    assign layer_1[1128] = ~layer_0[652]; 
    assign layer_1[1129] = ~layer_0[781]; 
    assign layer_1[1130] = ~layer_0[168]; 
    assign layer_1[1131] = ~layer_0[1067]; 
    assign layer_1[1132] = ~layer_0[1081]; 
    assign layer_1[1133] = ~layer_0[122]; 
    assign layer_1[1134] = ~layer_0[167]; 
    assign layer_1[1135] = ~layer_0[575]; 
    assign layer_1[1136] = ~layer_0[82]; 
    assign layer_1[1137] = ~layer_0[1230]; 
    assign layer_1[1138] = ~(layer_0[782] ^ layer_0[82]); 
    assign layer_1[1139] = ~layer_0[304]; 
    assign layer_1[1140] = ~layer_0[1015]; 
    assign layer_1[1141] = 1'b1; 
    assign layer_1[1142] = ~layer_0[82]; 
    assign layer_1[1143] = ~layer_0[493]; 
    assign layer_1[1144] = ~layer_0[371]; 
    assign layer_1[1145] = ~layer_0[457]; 
    assign layer_1[1146] = ~layer_0[48]; 
    assign layer_1[1147] = ~(layer_0[943] & layer_0[524]); 
    assign layer_1[1148] = ~layer_0[52]; 
    assign layer_1[1149] = ~layer_0[552]; 
    assign layer_1[1150] = ~(layer_0[1065] | layer_0[1111]); 
    assign layer_1[1151] = ~layer_0[806]; 
    assign layer_1[1152] = ~(layer_0[177] | layer_0[243]); 
    assign layer_1[1153] = ~layer_0[33]; 
    assign layer_1[1154] = ~layer_0[371]; 
    assign layer_1[1155] = ~layer_0[644]; 
    assign layer_1[1156] = ~layer_0[785]; 
    assign layer_1[1157] = ~(layer_0[620] ^ layer_0[578]); 
    assign layer_1[1158] = ~layer_0[532]; 
    assign layer_1[1159] = ~layer_0[581]; 
    assign layer_1[1160] = ~layer_0[371]; 
    assign layer_1[1161] = ~layer_0[934]; 
    assign layer_1[1162] = ~layer_0[1113]; 
    assign layer_1[1163] = ~layer_0[652]; 
    assign layer_1[1164] = ~layer_0[168]; 
    assign layer_1[1165] = ~layer_0[457]; 
    assign layer_1[1166] = ~layer_0[236]; 
    assign layer_1[1167] = ~layer_0[76]; 
    assign layer_1[1168] = ~layer_0[972]; 
    assign layer_1[1169] = ~layer_0[382]; 
    assign layer_1[1170] = ~layer_0[433]; 
    assign layer_1[1171] = ~layer_0[82]; 
    assign layer_1[1172] = ~layer_0[652]; 
    assign layer_1[1173] = ~layer_0[1054]; 
    assign layer_1[1174] = ~layer_0[691]; 
    assign layer_1[1175] = ~layer_0[541]; 
    assign layer_1[1176] = ~layer_0[691]; 
    assign layer_1[1177] = ~layer_0[855]; 
    assign layer_1[1178] = ~layer_0[700]; 
    assign layer_1[1179] = ~layer_0[644]; 
    assign layer_1[1180] = ~layer_0[639]; 
    assign layer_1[1181] = ~layer_0[139]; 
    assign layer_1[1182] = ~layer_0[231]; 
    assign layer_1[1183] = ~layer_0[652]; 
    assign layer_1[1184] = ~layer_0[1287]; 
    assign layer_1[1185] = ~layer_0[691]; 
    assign layer_1[1186] = ~layer_0[1160]; 
    assign layer_1[1187] = ~layer_0[1045]; 
    assign layer_1[1188] = ~layer_0[597]; 
    assign layer_1[1189] = ~layer_0[1099]; 
    assign layer_1[1190] = ~(layer_0[555] & layer_0[996]); 
    assign layer_1[1191] = 1'b0; 
    assign layer_1[1192] = ~layer_0[167]; 
    assign layer_1[1193] = ~layer_0[571]; 
    assign layer_1[1194] = ~layer_0[64]; 
    assign layer_1[1195] = ~(layer_0[579] & layer_0[962]); 
    assign layer_1[1196] = ~layer_0[709]; 
    assign layer_1[1197] = ~layer_0[855]; 
    assign layer_1[1198] = ~layer_0[652]; 
    assign layer_1[1199] = ~layer_0[1160]; 
    assign layer_1[1200] = ~layer_0[1194]; 
    assign layer_1[1201] = ~layer_0[691]; 
    assign layer_1[1202] = ~layer_0[652]; 
    assign layer_1[1203] = ~layer_0[208]; 
    assign layer_1[1204] = ~layer_0[1007]; 
    assign layer_1[1205] = ~layer_0[606]; 
    assign layer_1[1206] = ~layer_0[1081]; 
    assign layer_1[1207] = ~layer_0[577]; 
    assign layer_1[1208] = ~layer_0[443]; 
    assign layer_1[1209] = ~layer_0[1202]; 
    assign layer_1[1210] = ~(layer_0[208] & layer_0[52]); 
    assign layer_1[1211] = ~layer_0[589]; 
    assign layer_1[1212] = ~(layer_0[199] | layer_0[508]); 
    assign layer_1[1213] = ~layer_0[406]; 
    assign layer_1[1214] = ~layer_0[212]; 
    assign layer_1[1215] = ~layer_0[283]; 
    assign layer_1[1216] = ~layer_0[1267]; 
    assign layer_1[1217] = ~layer_0[856]; 
    assign layer_1[1218] = ~layer_0[1007]; 
    assign layer_1[1219] = ~layer_0[446]; 
    assign layer_1[1220] = ~layer_0[898]; 
    assign layer_1[1221] = ~layer_0[225]; 
    assign layer_1[1222] = ~(layer_0[202] | layer_0[575]); 
    assign layer_1[1223] = ~layer_0[1259]; 
    assign layer_1[1224] = ~layer_0[706]; 
    assign layer_1[1225] = ~layer_0[38]; 
    assign layer_1[1226] = ~layer_0[855]; 
    assign layer_1[1227] = ~layer_0[446]; 
    assign layer_1[1228] = ~layer_0[655]; 
    assign layer_1[1229] = ~layer_0[1085]; 
    assign layer_1[1230] = ~layer_0[768]; 
    assign layer_1[1231] = ~layer_0[1054]; 
    assign layer_1[1232] = ~(layer_0[996] | layer_0[700]); 
    assign layer_1[1233] = ~layer_0[433]; 
    assign layer_1[1234] = ~layer_0[1134]; 
    assign layer_1[1235] = ~layer_0[76]; 
    assign layer_1[1236] = ~layer_0[524]; 
    assign layer_1[1237] = ~layer_0[775]; 
    assign layer_1[1238] = ~layer_0[253]; 
    assign layer_1[1239] = ~layer_0[781]; 
    assign layer_1[1240] = ~layer_0[304]; 
    assign layer_1[1241] = layer_0[1079]; 
    assign layer_1[1242] = ~layer_0[657]; 
    assign layer_1[1243] = ~layer_0[371]; 
    assign layer_1[1244] = ~layer_0[652]; 
    assign layer_1[1245] = ~layer_0[470]; 
    assign layer_1[1246] = ~layer_0[354]; 
    assign layer_1[1247] = ~layer_0[589]; 
    assign layer_1[1248] = ~layer_0[799]; 
    assign layer_1[1249] = ~layer_0[1217]; 
    assign layer_1[1250] = ~layer_0[861]; 
    assign layer_1[1251] = ~layer_0[338]; 
    assign layer_1[1252] = ~layer_0[1081]; 
    assign layer_1[1253] = ~layer_0[2]; 
    assign layer_1[1254] = ~layer_0[90]; 
    assign layer_1[1255] = ~layer_0[781]; 
    assign layer_1[1256] = ~layer_0[90]; 
    assign layer_1[1257] = ~(layer_0[818] | layer_0[948]); 
    assign layer_1[1258] = ~layer_0[481]; 
    assign layer_1[1259] = ~layer_0[139]; 
    assign layer_1[1260] = ~layer_0[48]; 
    assign layer_1[1261] = ~layer_0[606]; 
    assign layer_1[1262] = ~layer_0[1190]; 
    assign layer_1[1263] = ~layer_0[569]; 
    assign layer_1[1264] = ~layer_0[1162]; 
    assign layer_1[1265] = ~(layer_0[218] & layer_0[495]); 
    assign layer_1[1266] = ~(layer_0[106] ^ layer_0[1042]); 
    assign layer_1[1267] = ~layer_0[820]; 
    assign layer_1[1268] = ~layer_0[652]; 
    assign layer_1[1269] = ~layer_0[168]; 
    assign layer_1[1270] = ~layer_0[1230]; 
    assign layer_1[1271] = ~(layer_0[1290] & layer_0[33]); 
    assign layer_1[1272] = ~layer_0[51]; 
    assign layer_1[1273] = ~layer_0[855]; 
    assign layer_1[1274] = ~layer_0[691]; 
    assign layer_1[1275] = layer_0[368]; 
    assign layer_1[1276] = ~layer_0[898]; 
    assign layer_1[1277] = ~layer_0[66]; 
    assign layer_1[1278] = ~layer_0[415]; 
    assign layer_1[1279] = ~layer_0[835]; 
    assign layer_1[1280] = ~layer_0[700]; 
    assign layer_1[1281] = ~layer_0[643]; 
    assign layer_1[1282] = ~layer_0[371]; 
    assign layer_1[1283] = ~layer_0[250]; 
    assign layer_1[1284] = ~layer_0[1190]; 
    assign layer_1[1285] = ~layer_0[1236]; 
    assign layer_1[1286] = ~layer_0[1022]; 
    assign layer_1[1287] = ~layer_0[1054]; 
    assign layer_1[1288] = ~layer_0[41]; 
    assign layer_1[1289] = ~layer_0[731]; 
    assign layer_1[1290] = ~layer_0[194]; 
    assign layer_1[1291] = ~layer_0[781]; 
    assign layer_1[1292] = ~layer_0[1054]; 
    assign layer_1[1293] = ~layer_0[111]; 
    assign layer_1[1294] = ~layer_0[1067]; 
    assign layer_1[1295] = ~layer_0[76]; 
    assign layer_1[1296] = ~layer_0[38]; 
    assign layer_1[1297] = ~layer_0[855]; 
    assign layer_1[1298] = ~layer_0[781]; 
    assign layer_1[1299] = ~layer_0[644]; 
    // Layer 2 ============================================================
    assign out[0] = ~(layer_1[151] & layer_1[546]); 
    assign out[1] = layer_1[646] ^ layer_1[914]; 
    assign out[2] = ~(layer_1[1187] | layer_1[100]); 
    assign out[3] = ~layer_1[462]; 
    assign out[4] = ~(layer_1[12] | layer_1[130]); 
    assign out[5] = ~layer_1[546]; 
    assign out[6] = ~layer_1[268]; 
    assign out[7] = ~layer_1[268]; 
    assign out[8] = ~layer_1[546]; 
    assign out[9] = ~layer_1[268]; 
    assign out[10] = ~layer_1[208]; 
    assign out[11] = ~layer_1[546]; 
    assign out[12] = ~layer_1[546]; 
    assign out[13] = ~layer_1[535]; 
    assign out[14] = ~(layer_1[642] | layer_1[284]); 
    assign out[15] = ~layer_1[535]; 
    assign out[16] = ~layer_1[130]; 
    assign out[17] = ~(layer_1[899] | layer_1[441]); 
    assign out[18] = ~(layer_1[349] & layer_1[208]); 
    assign out[19] = ~(layer_1[642] | layer_1[1046]); 
    assign out[20] = layer_1[135] & ~layer_1[268]; 
    assign out[21] = layer_1[1102] & ~layer_1[899]; 
    assign out[22] = ~layer_1[268]; 
    assign out[23] = ~(layer_1[642] | layer_1[535]); 
    assign out[24] = ~layer_1[130]; 
    assign out[25] = ~layer_1[642]; 
    assign out[26] = ~layer_1[546]; 
    assign out[27] = ~layer_1[535]; 
    assign out[28] = ~layer_1[535]; 
    assign out[29] = ~layer_1[535]; 
    assign out[30] = ~layer_1[546]; 
    assign out[31] = ~(layer_1[268] | layer_1[936]); 
    assign out[32] = ~layer_1[268]; 
    assign out[33] = ~(layer_1[130] | layer_1[268]); 
    assign out[34] = ~layer_1[268]; 
    assign out[35] = ~(layer_1[984] | layer_1[268]); 
    assign out[36] = ~(layer_1[268] | layer_1[130]); 
    assign out[37] = ~layer_1[268]; 
    assign out[38] = ~layer_1[535]; 
    assign out[39] = ~layer_1[535]; 
    assign out[40] = ~layer_1[546]; 
    assign out[41] = ~(layer_1[642] | layer_1[452]); 
    assign out[42] = ~layer_1[452]; 
    assign out[43] = ~(layer_1[12] | layer_1[535]); 
    assign out[44] = ~layer_1[535]; 
    assign out[45] = ~(layer_1[535] | layer_1[1197]); 
    assign out[46] = ~(layer_1[1046] | layer_1[546]); 
    assign out[47] = ~(layer_1[642] & layer_1[687]); 
    assign out[48] = ~layer_1[535]; 
    assign out[49] = ~layer_1[268]; 
    assign out[50] = ~layer_1[535]; 
    assign out[51] = ~layer_1[268]; 
    assign out[52] = layer_1[345] ^ layer_1[193]; 
    assign out[53] = ~layer_1[100]; 
    assign out[54] = ~layer_1[130]; 
    assign out[55] = layer_1[1213] & ~layer_1[113]; 
    assign out[56] = ~layer_1[268]; 
    assign out[57] = layer_1[567] ^ layer_1[464]; 
    assign out[58] = layer_1[1213] & ~layer_1[130]; 
    assign out[59] = ~layer_1[535]; 
    assign out[60] = ~(layer_1[208] & layer_1[151]); 
    assign out[61] = ~layer_1[535]; 
    assign out[62] = layer_1[809] & ~layer_1[130]; 
    assign out[63] = ~layer_1[535]; 
    assign out[64] = ~layer_1[268]; 
    assign out[65] = ~(layer_1[130] | layer_1[268]); 
    assign out[66] = ~layer_1[546]; 
    assign out[67] = ~layer_1[268]; 
    assign out[68] = ~layer_1[268]; 
    assign out[69] = ~(layer_1[151] | layer_1[1046]); 
    assign out[70] = layer_1[109] ^ layer_1[160]; 
    assign out[71] = ~(layer_1[151] & layer_1[208]); 
    assign out[72] = ~(layer_1[208] & layer_1[151]); 
    assign out[73] = ~layer_1[546]; 
    assign out[74] = ~layer_1[268]; 
    assign out[75] = layer_1[837] & ~layer_1[130]; 
    assign out[76] = ~layer_1[268]; 
    assign out[77] = layer_1[1276] & ~layer_1[268]; 
    assign out[78] = layer_1[837] & ~layer_1[546]; 
    assign out[79] = ~layer_1[546]; 
    assign out[80] = ~layer_1[546]; 
    assign out[81] = layer_1[1276] & ~layer_1[852]; 
    assign out[82] = ~layer_1[268]; 
    assign out[83] = layer_1[205] & ~layer_1[130]; 
    assign out[84] = ~(layer_1[208] & layer_1[452]); 
    assign out[85] = ~layer_1[535]; 
    assign out[86] = ~(layer_1[113] & layer_1[243]); 
    assign out[87] = ~layer_1[546]; 
    assign out[88] = ~layer_1[208]; 
    assign out[89] = ~layer_1[208]; 
    assign out[90] = ~layer_1[268]; 
    assign out[91] = ~(layer_1[441] | layer_1[105]); 
    assign out[92] = ~(layer_1[956] | layer_1[268]); 
    assign out[93] = ~layer_1[535]; 
    assign out[94] = ~layer_1[130]; 
    assign out[95] = ~(layer_1[208] & layer_1[208]); 
    assign out[96] = ~(layer_1[130] | layer_1[12]); 
    assign out[97] = ~layer_1[268]; 
    assign out[98] = ~layer_1[535]; 
    assign out[99] = ~(layer_1[268] | layer_1[130]); 
    assign out[100] = ~(layer_1[687] & layer_1[86]); 
    assign out[101] = ~(layer_1[86] | layer_1[311]); 
    assign out[102] = ~(layer_1[535] | layer_1[912]); 
    assign out[103] = ~layer_1[268]; 
    assign out[104] = ~(layer_1[452] | layer_1[460]); 
    assign out[105] = ~layer_1[535]; 
    assign out[106] = ~layer_1[546]; 
    assign out[107] = ~(layer_1[130] | layer_1[206]); 
    assign out[108] = ~layer_1[268]; 
    assign out[109] = ~layer_1[268]; 
    assign out[110] = ~layer_1[546]; 
    assign out[111] = ~(layer_1[1197] | layer_1[20]); 
    assign out[112] = ~(layer_1[130] | layer_1[326]); 
    assign out[113] = ~(layer_1[12] | layer_1[130]); 
    assign out[114] = ~(layer_1[546] & layer_1[535]); 
    assign out[115] = layer_1[464] ^ layer_1[567]; 
    assign out[116] = ~(layer_1[222] | layer_1[268]); 
    assign out[117] = ~(layer_1[441] | layer_1[268]); 
    assign out[118] = ~layer_1[268]; 
    assign out[119] = ~layer_1[268]; 
    assign out[120] = ~layer_1[546]; 
    assign out[121] = ~layer_1[268]; 
    assign out[122] = ~layer_1[208]; 
    assign out[123] = ~(layer_1[130] | layer_1[514]); 
    assign out[124] = ~layer_1[208]; 
    assign out[125] = ~layer_1[610]; 
    assign out[126] = layer_1[1102] & ~layer_1[105]; 
    assign out[127] = layer_1[567] ^ layer_1[464]; 
    assign out[128] = ~layer_1[535]; 
    assign out[129] = ~layer_1[535]; 
    assign out[130] = layer_1[747]; 
    assign out[131] = layer_1[715] | layer_1[276]; 
    assign out[132] = layer_1[997] | layer_1[77]; 
    assign out[133] = layer_1[1046] & layer_1[609]; 
    assign out[134] = layer_1[997]; 
    assign out[135] = layer_1[715] | layer_1[351]; 
    assign out[136] = layer_1[1105]; 
    assign out[137] = layer_1[1071] | layer_1[77]; 
    assign out[138] = layer_1[822] & layer_1[609]; 
    assign out[139] = layer_1[1222]; 
    assign out[140] = layer_1[1073]; 
    assign out[141] = layer_1[609]; 
    assign out[142] = layer_1[310] & layer_1[311]; 
    assign out[143] = layer_1[555] & layer_1[641]; 
    assign out[144] = layer_1[213] | layer_1[1073]; 
    assign out[145] = layer_1[609]; 
    assign out[146] = layer_1[609]; 
    assign out[147] = layer_1[170]; 
    assign out[148] = layer_1[715] | layer_1[515]; 
    assign out[149] = layer_1[170] & layer_1[1105]; 
    assign out[150] = layer_1[747]; 
    assign out[151] = layer_1[77] | layer_1[616]; 
    assign out[152] = layer_1[170]; 
    assign out[153] = ~layer_1[1241] | (layer_1[140] & layer_1[1241]); 
    assign out[154] = layer_1[213] | layer_1[276]; 
    assign out[155] = layer_1[1222] | layer_1[213]; 
    assign out[156] = layer_1[406]; 
    assign out[157] = ~layer_1[769] | (layer_1[769] & layer_1[1073]); 
    assign out[158] = layer_1[170] & layer_1[854]; 
    assign out[159] = layer_1[1073]; 
    assign out[160] = layer_1[555] & layer_1[387]; 
    assign out[161] = layer_1[204]; 
    assign out[162] = layer_1[977] & layer_1[822]; 
    assign out[163] = layer_1[747]; 
    assign out[164] = layer_1[822]; 
    assign out[165] = layer_1[555]; 
    assign out[166] = layer_1[609]; 
    assign out[167] = layer_1[555]; 
    assign out[168] = layer_1[1222] | layer_1[77]; 
    assign out[169] = layer_1[170]; 
    assign out[170] = layer_1[895] & layer_1[843]; 
    assign out[171] = layer_1[77] | layer_1[1222]; 
    assign out[172] = layer_1[715] | layer_1[276]; 
    assign out[173] = layer_1[1071] | layer_1[78]; 
    assign out[174] = layer_1[854] & layer_1[822]; 
    assign out[175] = layer_1[786]; 
    assign out[176] = layer_1[609] & layer_1[822]; 
    assign out[177] = layer_1[1145] | layer_1[60]; 
    assign out[178] = layer_1[1143]; 
    assign out[179] = layer_1[387] & layer_1[911]; 
    assign out[180] = layer_1[170] & layer_1[1145]; 
    assign out[181] = layer_1[1233] & layer_1[95]; 
    assign out[182] = layer_1[22] & layer_1[137]; 
    assign out[183] = layer_1[609]; 
    assign out[184] = layer_1[609]; 
    assign out[185] = layer_1[609]; 
    assign out[186] = ~(layer_1[1221] ^ layer_1[445]); 
    assign out[187] = layer_1[311] & layer_1[822]; 
    assign out[188] = layer_1[747]; 
    assign out[189] = layer_1[482]; 
    assign out[190] = layer_1[715]; 
    assign out[191] = layer_1[609]; 
    assign out[192] = layer_1[1222]; 
    assign out[193] = ~layer_1[104] | (layer_1[104] & layer_1[77]); 
    assign out[194] = layer_1[170]; 
    assign out[195] = layer_1[213] | layer_1[1071]; 
    assign out[196] = layer_1[1105]; 
    assign out[197] = layer_1[276] | layer_1[555]; 
    assign out[198] = layer_1[822] & layer_1[966]; 
    assign out[199] = layer_1[170] & layer_1[311]; 
    assign out[200] = layer_1[1145]; 
    assign out[201] = layer_1[406] & layer_1[1221]; 
    assign out[202] = layer_1[1145]; 
    assign out[203] = layer_1[60] & layer_1[1222]; 
    assign out[204] = layer_1[310] & layer_1[609]; 
    assign out[205] = layer_1[1145] | layer_1[482]; 
    assign out[206] = layer_1[609]; 
    assign out[207] = layer_1[170] & layer_1[310]; 
    assign out[208] = layer_1[1127] & layer_1[822]; 
    assign out[209] = layer_1[170] & layer_1[854]; 
    assign out[210] = layer_1[747]; 
    assign out[211] = layer_1[170]; 
    assign out[212] = layer_1[822] & layer_1[1073]; 
    assign out[213] = layer_1[747]; 
    assign out[214] = ~layer_1[1241] | (layer_1[1241] & layer_1[1143]); 
    assign out[215] = layer_1[213] | layer_1[655]; 
    assign out[216] = layer_1[77] | layer_1[997]; 
    assign out[217] = layer_1[170]; 
    assign out[218] = layer_1[822] & layer_1[609]; 
    assign out[219] = layer_1[77] | layer_1[60]; 
    assign out[220] = layer_1[170]; 
    assign out[221] = layer_1[822] & layer_1[1233]; 
    assign out[222] = layer_1[609]; 
    assign out[223] = layer_1[794] & layer_1[843]; 
    assign out[224] = layer_1[997] | layer_1[747]; 
    assign out[225] = ~layer_1[727] | (layer_1[213] & layer_1[727]); 
    assign out[226] = layer_1[237] & layer_1[1286]; 
    assign out[227] = layer_1[609]; 
    assign out[228] = ~layer_1[1241] | (layer_1[655] & layer_1[1241]); 
    assign out[229] = layer_1[609] & layer_1[834]; 
    assign out[230] = layer_1[60] & layer_1[736]; 
    assign out[231] = layer_1[715] & layer_1[581]; 
    assign out[232] = layer_1[895] & layer_1[843]; 
    assign out[233] = layer_1[822]; 
    assign out[234] = layer_1[609] & layer_1[1105]; 
    assign out[235] = layer_1[78] | layer_1[997]; 
    assign out[236] = layer_1[715] | layer_1[1222]; 
    assign out[237] = layer_1[1145]; 
    assign out[238] = layer_1[60] & layer_1[723]; 
    assign out[239] = layer_1[1063] & layer_1[854]; 
    assign out[240] = ~(layer_1[1271] ^ layer_1[895]); 
    assign out[241] = layer_1[1221] & layer_1[996]; 
    assign out[242] = layer_1[60] & layer_1[237]; 
    assign out[243] = layer_1[77] | layer_1[701]; 
    assign out[244] = layer_1[609]; 
    assign out[245] = layer_1[77] | layer_1[1222]; 
    assign out[246] = layer_1[609]; 
    assign out[247] = layer_1[170]; 
    assign out[248] = layer_1[325]; 
    assign out[249] = layer_1[822]; 
    assign out[250] = ~layer_1[898] | (layer_1[898] & layer_1[715]); 
    assign out[251] = layer_1[609]; 
    assign out[252] = layer_1[482]; 
    assign out[253] = layer_1[1200] & layer_1[715]; 
    assign out[254] = layer_1[555]; 
    assign out[255] = layer_1[1222] | layer_1[213]; 
    assign out[256] = ~layer_1[727] | (layer_1[77] & layer_1[727]); 
    assign out[257] = layer_1[1145] & layer_1[431]; 
    assign out[258] = layer_1[170]; 
    assign out[259] = layer_1[60] & layer_1[734]; 
    assign out[260] = ~layer_1[188]; 
    assign out[261] = layer_1[904] & ~layer_1[89]; 
    assign out[262] = layer_1[536] ^ layer_1[716]; 
    assign out[263] = layer_1[790]; 
    assign out[264] = layer_1[958] & ~layer_1[325]; 
    assign out[265] = ~(layer_1[188] & layer_1[460]); 
    assign out[266] = layer_1[551] & ~layer_1[356]; 
    assign out[267] = layer_1[581] ^ layer_1[1197]; 
    assign out[268] = layer_1[427]; 
    assign out[269] = layer_1[500] ^ layer_1[729]; 
    assign out[270] = layer_1[427]; 
    assign out[271] = layer_1[790]; 
    assign out[272] = layer_1[877] & ~layer_1[188]; 
    assign out[273] = layer_1[1225] & layer_1[944]; 
    assign out[274] = layer_1[1057] & ~layer_1[188]; 
    assign out[275] = layer_1[904] & ~layer_1[188]; 
    assign out[276] = layer_1[877] & ~layer_1[188]; 
    assign out[277] = layer_1[427]; 
    assign out[278] = layer_1[1125]; 
    assign out[279] = layer_1[356] ^ layer_1[436]; 
    assign out[280] = layer_1[995] & ~layer_1[356]; 
    assign out[281] = layer_1[283] | layer_1[321]; 
    assign out[282] = layer_1[944] & ~layer_1[188]; 
    assign out[283] = layer_1[1225] & ~layer_1[356]; 
    assign out[284] = layer_1[480]; 
    assign out[285] = layer_1[157] | layer_1[283]; 
    assign out[286] = layer_1[120] & ~layer_1[188]; 
    assign out[287] = layer_1[877] & layer_1[428]; 
    assign out[288] = layer_1[436] & ~layer_1[188]; 
    assign out[289] = layer_1[513] & layer_1[917]; 
    assign out[290] = layer_1[1288] ^ layer_1[581]; 
    assign out[291] = layer_1[551] ^ layer_1[188]; 
    assign out[292] = layer_1[904] ^ layer_1[188]; 
    assign out[293] = layer_1[427]; 
    assign out[294] = layer_1[1225] ^ layer_1[410]; 
    assign out[295] = layer_1[334]; 
    assign out[296] = layer_1[958]; 
    assign out[297] = layer_1[1170] ^ layer_1[581]; 
    assign out[298] = layer_1[836]; 
    assign out[299] = layer_1[904] & ~layer_1[188]; 
    assign out[300] = ~(layer_1[915] & layer_1[356]); 
    assign out[301] = layer_1[864] & ~layer_1[188]; 
    assign out[302] = layer_1[436] & ~layer_1[188]; 
    assign out[303] = layer_1[877] & layer_1[436]; 
    assign out[304] = ~layer_1[356]; 
    assign out[305] = layer_1[581] ^ layer_1[407]; 
    assign out[306] = layer_1[427]; 
    assign out[307] = layer_1[427]; 
    assign out[308] = layer_1[157] | layer_1[1023]; 
    assign out[309] = layer_1[1206] | layer_1[1226]; 
    assign out[310] = ~(layer_1[356] & layer_1[460]); 
    assign out[311] = layer_1[427]; 
    assign out[312] = layer_1[1225] & ~layer_1[543]; 
    assign out[313] = layer_1[843] ^ layer_1[699]; 
    assign out[314] = ~layer_1[188]; 
    assign out[315] = layer_1[356] ^ layer_1[904]; 
    assign out[316] = ~(layer_1[188] & layer_1[45]); 
    assign out[317] = layer_1[356] ^ layer_1[436]; 
    assign out[318] = layer_1[551] ^ layer_1[543]; 
    assign out[319] = layer_1[139] & layer_1[732]; 
    assign out[320] = layer_1[1170] ^ layer_1[581]; 
    assign out[321] = layer_1[944] & ~layer_1[543]; 
    assign out[322] = layer_1[427]; 
    assign out[323] = layer_1[904] & ~layer_1[188]; 
    assign out[324] = layer_1[851] ^ layer_1[517]; 
    assign out[325] = layer_1[1226] ^ layer_1[581]; 
    assign out[326] = layer_1[904] & ~layer_1[356]; 
    assign out[327] = layer_1[1297] ^ layer_1[581]; 
    assign out[328] = layer_1[201] ^ layer_1[581]; 
    assign out[329] = layer_1[1271] & ~layer_1[356]; 
    assign out[330] = layer_1[334]; 
    assign out[331] = layer_1[904] & ~layer_1[356]; 
    assign out[332] = layer_1[117] ^ layer_1[1071]; 
    assign out[333] = layer_1[618] | layer_1[1197]; 
    assign out[334] = layer_1[1180] & ~layer_1[915]; 
    assign out[335] = layer_1[1282] ^ layer_1[729]; 
    assign out[336] = layer_1[245] ^ layer_1[581]; 
    assign out[337] = layer_1[427] | layer_1[427]; 
    assign out[338] = ~layer_1[188]; 
    assign out[339] = layer_1[100]; 
    assign out[340] = layer_1[904] ^ layer_1[356]; 
    assign out[341] = layer_1[866] & layer_1[877]; 
    assign out[342] = layer_1[238]; 
    assign out[343] = layer_1[238] & layer_1[513]; 
    assign out[344] = layer_1[581] ^ layer_1[1226]; 
    assign out[345] = layer_1[409] & ~layer_1[356]; 
    assign out[346] = layer_1[513] & ~layer_1[855]; 
    assign out[347] = layer_1[877] & layer_1[157]; 
    assign out[348] = layer_1[407] ^ layer_1[581]; 
    assign out[349] = ~layer_1[188]; 
    assign out[350] = layer_1[944] & ~layer_1[188]; 
    assign out[351] = layer_1[259] | layer_1[788]; 
    assign out[352] = layer_1[581] ^ layer_1[245]; 
    assign out[353] = layer_1[124] & layer_1[971]; 
    assign out[354] = layer_1[427]; 
    assign out[355] = layer_1[877] & layer_1[904]; 
    assign out[356] = layer_1[1225] & ~layer_1[1232]; 
    assign out[357] = ~(layer_1[885] & layer_1[432]); 
    assign out[358] = layer_1[904] & ~layer_1[188]; 
    assign out[359] = layer_1[230] | layer_1[892]; 
    assign out[360] = layer_1[1163] & ~layer_1[188]; 
    assign out[361] = layer_1[428] & ~layer_1[715]; 
    assign out[362] = layer_1[26] ^ layer_1[117]; 
    assign out[363] = layer_1[877] & layer_1[1095]; 
    assign out[364] = ~(layer_1[233] & layer_1[188]); 
    assign out[365] = layer_1[859] ^ layer_1[624]; 
    assign out[366] = layer_1[245] ^ layer_1[581]; 
    assign out[367] = layer_1[1125]; 
    assign out[368] = ~layer_1[188] | (layer_1[188] & layer_1[428]); 
    assign out[369] = layer_1[356] ^ layer_1[904]; 
    assign out[370] = layer_1[1197] | layer_1[1206]; 
    assign out[371] = layer_1[1197] ^ layer_1[581]; 
    assign out[372] = layer_1[798] ^ layer_1[320]; 
    assign out[373] = layer_1[359]; 
    assign out[374] = layer_1[729] ^ layer_1[500]; 
    assign out[375] = ~layer_1[45]; 
    assign out[376] = layer_1[320]; 
    assign out[377] = layer_1[1197] ^ layer_1[581]; 
    assign out[378] = layer_1[359]; 
    assign out[379] = layer_1[436] & ~layer_1[188]; 
    assign out[380] = ~(layer_1[188] & layer_1[188]); 
    assign out[381] = layer_1[427]; 
    assign out[382] = layer_1[904] & ~layer_1[356]; 
    assign out[383] = layer_1[1125]; 
    assign out[384] = layer_1[427] | layer_1[863]; 
    assign out[385] = layer_1[359] | layer_1[1233]; 
    assign out[386] = layer_1[188] ^ layer_1[904]; 
    assign out[387] = layer_1[1205] ^ layer_1[26]; 
    assign out[388] = layer_1[995] & layer_1[124]; 
    assign out[389] = layer_1[581] ^ layer_1[120]; 
    assign out[390] = layer_1[106] & ~layer_1[415]; 
    assign out[391] = layer_1[798] ^ layer_1[914]; 
    assign out[392] = ~layer_1[866]; 
    assign out[393] = ~(layer_1[18] & layer_1[1283]); 
    assign out[394] = layer_1[904] ^ layer_1[937]; 
    assign out[395] = layer_1[937] ^ layer_1[436]; 
    assign out[396] = layer_1[189] ^ layer_1[109]; 
    assign out[397] = layer_1[436] & ~layer_1[76]; 
    assign out[398] = layer_1[321]; 
    assign out[399] = layer_1[208] ^ layer_1[866]; 
    assign out[400] = layer_1[100] ^ layer_1[682]; 
    assign out[401] = layer_1[72] & ~layer_1[1232]; 
    assign out[402] = layer_1[851] & ~layer_1[76]; 
    assign out[403] = layer_1[786] ^ layer_1[312]; 
    assign out[404] = layer_1[72]; 
    assign out[405] = layer_1[72] & ~layer_1[76]; 
    assign out[406] = layer_1[72] & ~layer_1[76]; 
    assign out[407] = layer_1[755] ^ layer_1[312]; 
    assign out[408] = layer_1[834] & ~layer_1[415]; 
    assign out[409] = layer_1[1298] & ~layer_1[866]; 
    assign out[410] = ~layer_1[100]; 
    assign out[411] = layer_1[72] & ~layer_1[76]; 
    assign out[412] = layer_1[456] ^ layer_1[937]; 
    assign out[413] = layer_1[937] ^ layer_1[160]; 
    assign out[414] = ~(layer_1[100] | layer_1[768]); 
    assign out[415] = layer_1[263] ^ layer_1[211]; 
    assign out[416] = layer_1[72]; 
    assign out[417] = layer_1[937] ^ layer_1[436]; 
    assign out[418] = layer_1[359] | layer_1[291]; 
    assign out[419] = layer_1[1037] & ~layer_1[866]; 
    assign out[420] = layer_1[618]; 
    assign out[421] = layer_1[538] ^ layer_1[758]; 
    assign out[422] = layer_1[46] ^ layer_1[442]; 
    assign out[423] = ~layer_1[415]; 
    assign out[424] = layer_1[875] ^ layer_1[1163]; 
    assign out[425] = layer_1[1234] & ~layer_1[866]; 
    assign out[426] = layer_1[937] ^ layer_1[496]; 
    assign out[427] = layer_1[436] ^ layer_1[937]; 
    assign out[428] = layer_1[321] & ~layer_1[387]; 
    assign out[429] = layer_1[834] ^ layer_1[854]; 
    assign out[430] = layer_1[316] ^ layer_1[786]; 
    assign out[431] = layer_1[186] ^ layer_1[76]; 
    assign out[432] = layer_1[76] ^ layer_1[1255]; 
    assign out[433] = layer_1[72] & ~layer_1[415]; 
    assign out[434] = layer_1[72]; 
    assign out[435] = layer_1[436] ^ layer_1[76]; 
    assign out[436] = layer_1[76] ^ layer_1[414]; 
    assign out[437] = layer_1[312] & ~layer_1[76]; 
    assign out[438] = layer_1[798] ^ layer_1[1234]; 
    assign out[439] = ~(layer_1[113] & layer_1[768]); 
    assign out[440] = layer_1[834] & ~layer_1[866]; 
    assign out[441] = layer_1[416] | layer_1[428]; 
    assign out[442] = layer_1[72]; 
    assign out[443] = layer_1[1101] ^ layer_1[353]; 
    assign out[444] = layer_1[875] ^ layer_1[987]; 
    assign out[445] = layer_1[442] | layer_1[146]; 
    assign out[446] = ~layer_1[100]; 
    assign out[447] = layer_1[353] ^ layer_1[257]; 
    assign out[448] = layer_1[937] ^ layer_1[904]; 
    assign out[449] = layer_1[146] | layer_1[442]; 
    assign out[450] = layer_1[186] ^ layer_1[1232]; 
    assign out[451] = layer_1[66] ^ layer_1[937]; 
    assign out[452] = layer_1[1234] ^ layer_1[937]; 
    assign out[453] = layer_1[109] ^ layer_1[189]; 
    assign out[454] = layer_1[443] & ~layer_1[100]; 
    assign out[455] = layer_1[1234] ^ layer_1[937]; 
    assign out[456] = layer_1[1239] ^ layer_1[818]; 
    assign out[457] = layer_1[321]; 
    assign out[458] = layer_1[1234] & ~layer_1[76]; 
    assign out[459] = layer_1[386] & ~layer_1[866]; 
    assign out[460] = layer_1[937] ^ layer_1[436]; 
    assign out[461] = layer_1[100] ^ layer_1[546]; 
    assign out[462] = layer_1[641] ^ layer_1[316]; 
    assign out[463] = layer_1[76] ^ layer_1[436]; 
    assign out[464] = layer_1[641] ^ layer_1[331]; 
    assign out[465] = ~layer_1[1283]; 
    assign out[466] = layer_1[146] | layer_1[153]; 
    assign out[467] = layer_1[442] | layer_1[252]; 
    assign out[468] = layer_1[1121] & ~layer_1[866]; 
    assign out[469] = layer_1[1234] ^ layer_1[76]; 
    assign out[470] = layer_1[321]; 
    assign out[471] = layer_1[72] & layer_1[72]; 
    assign out[472] = layer_1[1129] & ~layer_1[866]; 
    assign out[473] = layer_1[618]; 
    assign out[474] = layer_1[72] & ~layer_1[76]; 
    assign out[475] = layer_1[987] ^ layer_1[353]; 
    assign out[476] = ~(layer_1[866] & layer_1[243]); 
    assign out[477] = layer_1[937] ^ layer_1[456]; 
    assign out[478] = layer_1[1017] ^ layer_1[753]; 
    assign out[479] = layer_1[633] | layer_1[153]; 
    assign out[480] = layer_1[186] & ~layer_1[76]; 
    assign out[481] = layer_1[321] & ~layer_1[387]; 
    assign out[482] = layer_1[1234] & ~layer_1[76]; 
    assign out[483] = layer_1[252] | layer_1[153]; 
    assign out[484] = layer_1[1234] ^ layer_1[76]; 
    assign out[485] = layer_1[146] | layer_1[785]; 
    assign out[486] = layer_1[875] ^ layer_1[987]; 
    assign out[487] = layer_1[613] ^ layer_1[72]; 
    assign out[488] = layer_1[252] | layer_1[442]; 
    assign out[489] = ~(layer_1[171] & layer_1[1283]); 
    assign out[490] = layer_1[1163] ^ layer_1[875]; 
    assign out[491] = layer_1[386] & ~layer_1[100]; 
    assign out[492] = layer_1[72] & ~layer_1[301]; 
    assign out[493] = layer_1[987] ^ layer_1[353]; 
    assign out[494] = layer_1[64] | layer_1[146]; 
    assign out[495] = layer_1[889] ^ layer_1[874]; 
    assign out[496] = ~(layer_1[100] | layer_1[346]); 
    assign out[497] = layer_1[153] | layer_1[526]; 
    assign out[498] = layer_1[436] ^ layer_1[937]; 
    assign out[499] = layer_1[937] ^ layer_1[904]; 
    assign out[500] = layer_1[42] ^ layer_1[1040]; 
    assign out[501] = layer_1[914] & ~layer_1[798]; 
    assign out[502] = layer_1[72]; 
    assign out[503] = layer_1[798] ^ layer_1[645]; 
    assign out[504] = layer_1[1121] & ~layer_1[100]; 
    assign out[505] = layer_1[987] ^ layer_1[353]; 
    assign out[506] = layer_1[441] & ~layer_1[866]; 
    assign out[507] = layer_1[866] ^ layer_1[637]; 
    assign out[508] = layer_1[591] ^ layer_1[1246]; 
    assign out[509] = layer_1[353] ^ layer_1[1163]; 
    assign out[510] = layer_1[1121] & ~layer_1[76]; 
    assign out[511] = layer_1[1159] & layer_1[1153]; 
    assign out[512] = layer_1[72] & layer_1[72]; 
    assign out[513] = layer_1[1121] & ~layer_1[76]; 
    assign out[514] = layer_1[1234]; 
    assign out[515] = layer_1[415] ^ layer_1[208]; 
    assign out[516] = layer_1[353] ^ layer_1[987]; 
    assign out[517] = layer_1[76] ^ layer_1[186]; 
    assign out[518] = layer_1[428] | layer_1[334]; 
    assign out[519] = layer_1[618] | layer_1[428]; 
    assign out[520] = layer_1[866] & ~layer_1[184]; 
    assign out[521] = layer_1[216] & ~layer_1[1163]; 
    assign out[522] = layer_1[50] & ~layer_1[670]; 
    assign out[523] = layer_1[404] ^ layer_1[184]; 
    assign out[524] = layer_1[194] ^ layer_1[941]; 
    assign out[525] = ~(layer_1[489] | layer_1[1157]); 
    assign out[526] = layer_1[1210] & ~layer_1[556]; 
    assign out[527] = ~(layer_1[1146] | layer_1[139]); 
    assign out[528] = layer_1[113] & ~layer_1[977]; 
    assign out[529] = ~layer_1[883]; 
    assign out[530] = ~layer_1[139]; 
    assign out[531] = layer_1[886] & ~layer_1[139]; 
    assign out[532] = ~layer_1[708]; 
    assign out[533] = ~(layer_1[736] | layer_1[469]); 
    assign out[534] = layer_1[372] & ~layer_1[1021]; 
    assign out[535] = layer_1[933] & ~layer_1[139]; 
    assign out[536] = layer_1[113] & ~layer_1[977]; 
    assign out[537] = ~layer_1[139]; 
    assign out[538] = ~(layer_1[1260] | layer_1[139]); 
    assign out[539] = ~(layer_1[966] | layer_1[1118]); 
    assign out[540] = ~(layer_1[1157] | layer_1[139]); 
    assign out[541] = layer_1[385] & ~layer_1[139]; 
    assign out[542] = ~layer_1[139]; 
    assign out[543] = ~layer_1[139]; 
    assign out[544] = layer_1[1175] & ~layer_1[1053]; 
    assign out[545] = ~(layer_1[195] | layer_1[766]); 
    assign out[546] = ~(layer_1[1061] | layer_1[888]); 
    assign out[547] = ~(layer_1[708] | layer_1[1139]); 
    assign out[548] = ~(layer_1[724] | layer_1[708]); 
    assign out[549] = ~layer_1[382]; 
    assign out[550] = ~(layer_1[653] | layer_1[1157]); 
    assign out[551] = ~(layer_1[757] | layer_1[708]); 
    assign out[552] = layer_1[1210] & ~layer_1[139]; 
    assign out[553] = ~layer_1[929]; 
    assign out[554] = layer_1[322] & ~layer_1[184]; 
    assign out[555] = layer_1[113] & ~layer_1[1251]; 
    assign out[556] = ~layer_1[139]; 
    assign out[557] = layer_1[591] & ~layer_1[685]; 
    assign out[558] = layer_1[216] & ~layer_1[218]; 
    assign out[559] = layer_1[952] & ~layer_1[199]; 
    assign out[560] = layer_1[1210] & ~layer_1[924]; 
    assign out[561] = ~(layer_1[676] | layer_1[1007]); 
    assign out[562] = layer_1[898] & ~layer_1[724]; 
    assign out[563] = ~(layer_1[345] | layer_1[1157]); 
    assign out[564] = ~(layer_1[1139] | layer_1[640]); 
    assign out[565] = layer_1[113] & ~layer_1[653]; 
    assign out[566] = layer_1[1210] & ~layer_1[1053]; 
    assign out[567] = layer_1[1210] & ~layer_1[653]; 
    assign out[568] = ~(layer_1[139] | layer_1[657]); 
    assign out[569] = layer_1[886] & ~layer_1[85]; 
    assign out[570] = ~layer_1[139]; 
    assign out[571] = layer_1[1224] & ~layer_1[17]; 
    assign out[572] = layer_1[422] & ~layer_1[802]; 
    assign out[573] = layer_1[22] ^ layer_1[310]; 
    assign out[574] = ~(layer_1[139] | layer_1[1157]); 
    assign out[575] = layer_1[249] & ~layer_1[724]; 
    assign out[576] = ~(layer_1[139] | layer_1[195]); 
    assign out[577] = layer_1[1210] & ~layer_1[653]; 
    assign out[578] = ~(layer_1[1118] | layer_1[195]); 
    assign out[579] = ~layer_1[139]; 
    assign out[580] = layer_1[898] & ~layer_1[470]; 
    assign out[581] = layer_1[1224] & ~layer_1[1045]; 
    assign out[582] = ~layer_1[1099]; 
    assign out[583] = layer_1[1210] & ~layer_1[653]; 
    assign out[584] = ~(layer_1[451] | layer_1[139]); 
    assign out[585] = layer_1[1217] ^ layer_1[1167]; 
    assign out[586] = ~(layer_1[1146] | layer_1[195]); 
    assign out[587] = ~(layer_1[184] | layer_1[139]); 
    assign out[588] = layer_1[275] & ~layer_1[929]; 
    assign out[589] = ~layer_1[708]; 
    assign out[590] = ~(layer_1[966] & layer_1[966]); 
    assign out[591] = layer_1[422] & ~layer_1[17]; 
    assign out[592] = ~(layer_1[195] | layer_1[708]); 
    assign out[593] = layer_1[1162] & ~layer_1[195]; 
    assign out[594] = ~(layer_1[924] | layer_1[451]); 
    assign out[595] = layer_1[698] & ~layer_1[1264]; 
    assign out[596] = ~layer_1[139]; 
    assign out[597] = layer_1[169] & ~layer_1[1125]; 
    assign out[598] = ~layer_1[1157]; 
    assign out[599] = ~(layer_1[324] | layer_1[708]); 
    assign out[600] = ~(layer_1[195] | layer_1[1146]); 
    assign out[601] = ~layer_1[908]; 
    assign out[602] = layer_1[1224] & ~layer_1[632]; 
    assign out[603] = layer_1[1053] ^ layer_1[372]; 
    assign out[604] = ~layer_1[139]; 
    assign out[605] = ~(layer_1[883] | layer_1[494]); 
    assign out[606] = ~(layer_1[883] | layer_1[278]); 
    assign out[607] = ~(layer_1[977] | layer_1[708]); 
    assign out[608] = layer_1[1210] & ~layer_1[653]; 
    assign out[609] = ~(layer_1[1276] | layer_1[1146]); 
    assign out[610] = ~(layer_1[1007] | layer_1[139]); 
    assign out[611] = ~layer_1[708]; 
    assign out[612] = layer_1[422] & ~layer_1[1265]; 
    assign out[613] = ~(layer_1[1276] & layer_1[1241]); 
    assign out[614] = layer_1[632] ^ layer_1[767]; 
    assign out[615] = layer_1[1175] & ~layer_1[17]; 
    assign out[616] = ~(layer_1[199] | layer_1[1157]); 
    assign out[617] = layer_1[105] & ~layer_1[582]; 
    assign out[618] = ~(layer_1[908] | layer_1[1139]); 
    assign out[619] = ~(layer_1[1072] | layer_1[1146]); 
    assign out[620] = ~(layer_1[1146] | layer_1[1030]); 
    assign out[621] = layer_1[1217] ^ layer_1[591]; 
    assign out[622] = ~(layer_1[1139] | layer_1[1146]); 
    assign out[623] = layer_1[591] & ~layer_1[502]; 
    assign out[624] = ~(layer_1[1146] | layer_1[1139]); 
    assign out[625] = layer_1[886] & ~layer_1[409]; 
    assign out[626] = ~(layer_1[139] | layer_1[708]); 
    assign out[627] = layer_1[18] ^ layer_1[929]; 
    assign out[628] = ~layer_1[1007]; 
    assign out[629] = ~layer_1[139]; 
    assign out[630] = ~(layer_1[139] | layer_1[708]); 
    assign out[631] = ~(layer_1[1139] | layer_1[708]); 
    assign out[632] = layer_1[113] & ~layer_1[280]; 
    assign out[633] = layer_1[113] & ~layer_1[17]; 
    assign out[634] = ~(layer_1[708] | layer_1[280]); 
    assign out[635] = layer_1[113] & ~layer_1[17]; 
    assign out[636] = layer_1[169] & ~layer_1[220]; 
    assign out[637] = ~(layer_1[883] | layer_1[426]); 
    assign out[638] = ~layer_1[883]; 
    assign out[639] = layer_1[290] & ~layer_1[966]; 
    assign out[640] = ~layer_1[139]; 
    assign out[641] = ~(layer_1[195] | layer_1[708]); 
    assign out[642] = layer_1[1188] ^ layer_1[531]; 
    assign out[643] = ~layer_1[1099]; 
    assign out[644] = layer_1[113] & ~layer_1[363]; 
    assign out[645] = layer_1[591] & ~layer_1[1139]; 
    assign out[646] = ~layer_1[1099]; 
    assign out[647] = ~(layer_1[842] | layer_1[1007]); 
    assign out[648] = ~layer_1[924]; 
    assign out[649] = layer_1[886] & ~layer_1[802]; 
    assign out[650] = layer_1[814] & ~layer_1[1063]; 
    assign out[651] = layer_1[189] ^ layer_1[40]; 
    assign out[652] = layer_1[1280]; 
    assign out[653] = layer_1[53] & ~layer_1[866]; 
    assign out[654] = layer_1[940] & ~layer_1[530]; 
    assign out[655] = ~(layer_1[937] | layer_1[526]); 
    assign out[656] = layer_1[1232]; 
    assign out[657] = layer_1[814] & ~layer_1[917]; 
    assign out[658] = layer_1[494]; 
    assign out[659] = layer_1[761] & ~layer_1[92]; 
    assign out[660] = layer_1[814] & ~layer_1[1071]; 
    assign out[661] = layer_1[40] ^ layer_1[834]; 
    assign out[662] = layer_1[144] & ~layer_1[987]; 
    assign out[663] = layer_1[897] & ~layer_1[1275]; 
    assign out[664] = layer_1[1232] & ~layer_1[17]; 
    assign out[665] = layer_1[959] & ~layer_1[1063]; 
    assign out[666] = ~(layer_1[160] & layer_1[793]); 
    assign out[667] = layer_1[175] & ~layer_1[396]; 
    assign out[668] = layer_1[823] & ~layer_1[526]; 
    assign out[669] = layer_1[670] & ~layer_1[1065]; 
    assign out[670] = layer_1[59] & ~layer_1[1101]; 
    assign out[671] = layer_1[1265] & ~layer_1[937]; 
    assign out[672] = ~(layer_1[937] | layer_1[1071]); 
    assign out[673] = layer_1[1033] & ~layer_1[938]; 
    assign out[674] = ~(layer_1[610] & layer_1[817]); 
    assign out[675] = layer_1[954] & ~layer_1[1126]; 
    assign out[676] = layer_1[1200] & ~layer_1[1063]; 
    assign out[677] = layer_1[1265] & ~layer_1[1071]; 
    assign out[678] = layer_1[852] & ~layer_1[816]; 
    assign out[679] = layer_1[452] & ~layer_1[794]; 
    assign out[680] = layer_1[670] & ~layer_1[298]; 
    assign out[681] = layer_1[1265] & ~layer_1[1071]; 
    assign out[682] = ~(layer_1[937] | layer_1[1071]); 
    assign out[683] = layer_1[814] & ~layer_1[408]; 
    assign out[684] = layer_1[573] & ~layer_1[937]; 
    assign out[685] = layer_1[59] & ~layer_1[530]; 
    assign out[686] = layer_1[1265] & ~layer_1[832]; 
    assign out[687] = ~layer_1[861] | (layer_1[861] & layer_1[531]); 
    assign out[688] = layer_1[814] & ~layer_1[326]; 
    assign out[689] = layer_1[814] & ~layer_1[1071]; 
    assign out[690] = ~(layer_1[917] | layer_1[194]); 
    assign out[691] = layer_1[29] & ~layer_1[110]; 
    assign out[692] = layer_1[959] & ~layer_1[1063]; 
    assign out[693] = layer_1[382] & ~layer_1[703]; 
    assign out[694] = layer_1[1265] & ~layer_1[938]; 
    assign out[695] = ~layer_1[1063]; 
    assign out[696] = layer_1[175] & ~layer_1[530]; 
    assign out[697] = layer_1[814] & ~layer_1[917]; 
    assign out[698] = layer_1[823] & ~layer_1[1071]; 
    assign out[699] = layer_1[823] & ~layer_1[1071]; 
    assign out[700] = layer_1[814] & ~layer_1[778]; 
    assign out[701] = layer_1[959] & ~layer_1[1095]; 
    assign out[702] = layer_1[1265] & ~layer_1[1071]; 
    assign out[703] = layer_1[814] & ~layer_1[565]; 
    assign out[704] = layer_1[897] & ~layer_1[937]; 
    assign out[705] = layer_1[803]; 
    assign out[706] = layer_1[386] & ~layer_1[1267]; 
    assign out[707] = ~(layer_1[703] | layer_1[1071]); 
    assign out[708] = layer_1[452] & ~layer_1[794]; 
    assign out[709] = layer_1[670] & ~layer_1[1275]; 
    assign out[710] = layer_1[99]; 
    assign out[711] = ~layer_1[159] | (layer_1[159] & layer_1[343]); 
    assign out[712] = layer_1[1182]; 
    assign out[713] = ~layer_1[962] | (layer_1[1265] & layer_1[962]); 
    assign out[714] = layer_1[320] & ~layer_1[917]; 
    assign out[715] = layer_1[206] & ~layer_1[565]; 
    assign out[716] = layer_1[823] & ~layer_1[817]; 
    assign out[717] = layer_1[814] & ~layer_1[937]; 
    assign out[718] = layer_1[1294] & ~layer_1[110]; 
    assign out[719] = layer_1[946] & ~layer_1[704]; 
    assign out[720] = layer_1[538] & ~layer_1[1267]; 
    assign out[721] = layer_1[814] & ~layer_1[917]; 
    assign out[722] = layer_1[515] & ~layer_1[832]; 
    assign out[723] = layer_1[53] & ~layer_1[1065]; 
    assign out[724] = layer_1[814] & ~layer_1[1063]; 
    assign out[725] = layer_1[1232] & ~layer_1[92]; 
    assign out[726] = layer_1[368] & ~layer_1[298]; 
    assign out[727] = layer_1[112] & ~layer_1[1063]; 
    assign out[728] = layer_1[1265] & ~layer_1[866]; 
    assign out[729] = layer_1[420] & ~layer_1[1071]; 
    assign out[730] = layer_1[814] & ~layer_1[1063]; 
    assign out[731] = layer_1[183] & ~layer_1[346]; 
    assign out[732] = layer_1[897] & ~layer_1[925]; 
    assign out[733] = ~(layer_1[1221] & layer_1[883]); 
    assign out[734] = layer_1[1265] & ~layer_1[110]; 
    assign out[735] = ~layer_1[1090]; 
    assign out[736] = layer_1[682] & ~layer_1[794]; 
    assign out[737] = layer_1[814] & ~layer_1[565]; 
    assign out[738] = layer_1[189] & ~layer_1[782]; 
    assign out[739] = layer_1[814] & ~layer_1[1063]; 
    assign out[740] = layer_1[823]; 
    assign out[741] = layer_1[761] & ~layer_1[1063]; 
    assign out[742] = layer_1[1265] & ~layer_1[1071]; 
    assign out[743] = layer_1[1265] & ~layer_1[526]; 
    assign out[744] = layer_1[823] & ~layer_1[1071]; 
    assign out[745] = ~(layer_1[888] | layer_1[328]); 
    assign out[746] = layer_1[538] & ~layer_1[283]; 
    assign out[747] = layer_1[29] & ~layer_1[1071]; 
    assign out[748] = layer_1[386] & ~layer_1[1194]; 
    assign out[749] = layer_1[897] & ~layer_1[863]; 
    assign out[750] = ~(layer_1[1071] | layer_1[1063]); 
    assign out[751] = layer_1[538] & ~layer_1[76]; 
    assign out[752] = layer_1[1056] & ~layer_1[1063]; 
    assign out[753] = layer_1[761] & ~layer_1[565]; 
    assign out[754] = layer_1[839] & ~layer_1[1063]; 
    assign out[755] = ~layer_1[346] | (layer_1[236] & layer_1[346]); 
    assign out[756] = layer_1[1265] & ~layer_1[565]; 
    assign out[757] = layer_1[1265] & ~layer_1[212]; 
    assign out[758] = layer_1[761] & ~layer_1[346]; 
    assign out[759] = layer_1[999] & ~layer_1[100]; 
    assign out[760] = layer_1[917] ^ layer_1[400]; 
    assign out[761] = layer_1[897] & ~layer_1[703]; 
    assign out[762] = layer_1[1265] & ~layer_1[1071]; 
    assign out[763] = layer_1[823] & ~layer_1[1095]; 
    assign out[764] = layer_1[823] ^ layer_1[907]; 
    assign out[765] = ~layer_1[1071]; 
    assign out[766] = layer_1[1265]; 
    assign out[767] = layer_1[400] & ~layer_1[917]; 
    assign out[768] = layer_1[1265] & ~layer_1[76]; 
    assign out[769] = layer_1[866] ^ layer_1[666]; 
    assign out[770] = layer_1[707] & ~layer_1[866]; 
    assign out[771] = layer_1[946] & ~layer_1[76]; 
    assign out[772] = layer_1[452] & ~layer_1[1221]; 
    assign out[773] = layer_1[162] & ~layer_1[1060]; 
    assign out[774] = layer_1[856] & ~layer_1[1063]; 
    assign out[775] = layer_1[1030] & ~layer_1[703]; 
    assign out[776] = layer_1[1131] & ~layer_1[937]; 
    assign out[777] = ~(layer_1[105] & layer_1[1090]); 
    assign out[778] = layer_1[897] & ~layer_1[159]; 
    assign out[779] = layer_1[691]; 
    assign out[780] = layer_1[1212] ^ layer_1[870]; 
    assign out[781] = layer_1[1152] | layer_1[602]; 
    assign out[782] = ~layer_1[1199]; 
    assign out[783] = ~layer_1[1199]; 
    assign out[784] = layer_1[578] | layer_1[830]; 
    assign out[785] = layer_1[844] ^ layer_1[532]; 
    assign out[786] = layer_1[276] ^ layer_1[685]; 
    assign out[787] = layer_1[674] & ~layer_1[441]; 
    assign out[788] = layer_1[1074]; 
    assign out[789] = layer_1[1212] & ~layer_1[60]; 
    assign out[790] = layer_1[1212] & ~layer_1[514]; 
    assign out[791] = layer_1[716]; 
    assign out[792] = layer_1[411] ^ layer_1[864]; 
    assign out[793] = layer_1[1212] & ~layer_1[1187]; 
    assign out[794] = layer_1[127] & layer_1[830]; 
    assign out[795] = ~layer_1[1199]; 
    assign out[796] = layer_1[653] ^ layer_1[411]; 
    assign out[797] = ~layer_1[1199]; 
    assign out[798] = layer_1[716]; 
    assign out[799] = layer_1[1074]; 
    assign out[800] = ~layer_1[1199]; 
    assign out[801] = layer_1[716] | layer_1[541]; 
    assign out[802] = ~layer_1[1187]; 
    assign out[803] = layer_1[830] | layer_1[756]; 
    assign out[804] = layer_1[923] ^ layer_1[756]; 
    assign out[805] = layer_1[923] ^ layer_1[1294]; 
    assign out[806] = layer_1[852] ^ layer_1[276]; 
    assign out[807] = layer_1[844] ^ layer_1[547]; 
    assign out[808] = layer_1[1207] ^ layer_1[958]; 
    assign out[809] = layer_1[276] ^ layer_1[685]; 
    assign out[810] = layer_1[852] & ~layer_1[1187]; 
    assign out[811] = layer_1[532]; 
    assign out[812] = layer_1[236] ^ layer_1[1212]; 
    assign out[813] = layer_1[1185] & ~layer_1[1187]; 
    assign out[814] = ~(layer_1[1199] & layer_1[284]); 
    assign out[815] = layer_1[1212] & ~layer_1[992]; 
    assign out[816] = ~layer_1[1199]; 
    assign out[817] = layer_1[276] ^ layer_1[685]; 
    assign out[818] = layer_1[515] & ~layer_1[441]; 
    assign out[819] = layer_1[1212] & ~layer_1[938]; 
    assign out[820] = layer_1[1212] & ~layer_1[411]; 
    assign out[821] = layer_1[923] ^ layer_1[1188]; 
    assign out[822] = layer_1[653]; 
    assign out[823] = layer_1[4] ^ layer_1[31]; 
    assign out[824] = layer_1[325] | layer_1[68]; 
    assign out[825] = layer_1[254] & layer_1[685]; 
    assign out[826] = layer_1[870] ^ layer_1[941]; 
    assign out[827] = ~layer_1[1199]; 
    assign out[828] = ~layer_1[1199]; 
    assign out[829] = layer_1[852] ^ layer_1[276]; 
    assign out[830] = layer_1[1212] & ~layer_1[514]; 
    assign out[831] = layer_1[532]; 
    assign out[832] = layer_1[1074]; 
    assign out[833] = layer_1[756] ^ layer_1[779]; 
    assign out[834] = layer_1[532]; 
    assign out[835] = ~(layer_1[750] & layer_1[246]); 
    assign out[836] = layer_1[653]; 
    assign out[837] = layer_1[937] & ~layer_1[799]; 
    assign out[838] = layer_1[1210] & ~layer_1[411]; 
    assign out[839] = ~(layer_1[1199] & layer_1[297]); 
    assign out[840] = layer_1[1210] & ~layer_1[1187]; 
    assign out[841] = layer_1[716] & ~layer_1[411]; 
    assign out[842] = layer_1[744] & ~layer_1[441]; 
    assign out[843] = layer_1[685] & ~layer_1[441]; 
    assign out[844] = layer_1[1212] ^ layer_1[997]; 
    assign out[845] = ~layer_1[1199]; 
    assign out[846] = layer_1[937] & ~layer_1[728]; 
    assign out[847] = layer_1[278] ^ layer_1[430]; 
    assign out[848] = layer_1[1210] ^ layer_1[514]; 
    assign out[849] = layer_1[844] ^ layer_1[532]; 
    assign out[850] = layer_1[539] & ~layer_1[284]; 
    assign out[851] = layer_1[430] ^ layer_1[278]; 
    assign out[852] = ~layer_1[108]; 
    assign out[853] = layer_1[1212] & ~layer_1[514]; 
    assign out[854] = layer_1[703] & layer_1[756]; 
    assign out[855] = layer_1[201] ^ layer_1[882]; 
    assign out[856] = layer_1[1210] & ~layer_1[237]; 
    assign out[857] = layer_1[716] & ~layer_1[514]; 
    assign out[858] = ~layer_1[108]; 
    assign out[859] = layer_1[716]; 
    assign out[860] = layer_1[756] ^ layer_1[1019]; 
    assign out[861] = layer_1[602]; 
    assign out[862] = layer_1[602]; 
    assign out[863] = ~layer_1[1199]; 
    assign out[864] = layer_1[9] ^ layer_1[1240]; 
    assign out[865] = layer_1[937] ^ layer_1[799]; 
    assign out[866] = layer_1[552] | layer_1[830]; 
    assign out[867] = layer_1[844] ^ layer_1[532]; 
    assign out[868] = layer_1[716]; 
    assign out[869] = ~(layer_1[1187] | layer_1[463]); 
    assign out[870] = ~layer_1[1199]; 
    assign out[871] = layer_1[685]; 
    assign out[872] = layer_1[256] ^ layer_1[923]; 
    assign out[873] = layer_1[552] | layer_1[830]; 
    assign out[874] = layer_1[1082] & ~layer_1[441]; 
    assign out[875] = layer_1[716]; 
    assign out[876] = layer_1[1143] ^ layer_1[532]; 
    assign out[877] = layer_1[532] | layer_1[716]; 
    assign out[878] = layer_1[228] ^ layer_1[217]; 
    assign out[879] = layer_1[653]; 
    assign out[880] = layer_1[1212] & ~layer_1[236]; 
    assign out[881] = layer_1[1212]; 
    assign out[882] = layer_1[941] & layer_1[1212]; 
    assign out[883] = layer_1[254] ^ layer_1[514]; 
    assign out[884] = layer_1[941] ^ layer_1[923]; 
    assign out[885] = ~(layer_1[441] | layer_1[1197]); 
    assign out[886] = layer_1[514] ^ layer_1[254]; 
    assign out[887] = layer_1[602]; 
    assign out[888] = layer_1[1210] & ~layer_1[514]; 
    assign out[889] = layer_1[1212] ^ layer_1[411]; 
    assign out[890] = layer_1[532] & ~layer_1[992]; 
    assign out[891] = layer_1[552] | layer_1[830]; 
    assign out[892] = layer_1[1029] ^ layer_1[716]; 
    assign out[893] = layer_1[236] ^ layer_1[1212]; 
    assign out[894] = layer_1[547]; 
    assign out[895] = layer_1[923] ^ layer_1[756]; 
    assign out[896] = layer_1[756] | layer_1[779]; 
    assign out[897] = layer_1[602] & ~layer_1[463]; 
    assign out[898] = ~layer_1[108]; 
    assign out[899] = ~layer_1[1199]; 
    assign out[900] = ~(layer_1[888] & layer_1[283]); 
    assign out[901] = layer_1[236] ^ layer_1[1212]; 
    assign out[902] = layer_1[1212]; 
    assign out[903] = layer_1[653] & ~layer_1[1187]; 
    assign out[904] = layer_1[716]; 
    assign out[905] = layer_1[716]; 
    assign out[906] = layer_1[532] | layer_1[716]; 
    assign out[907] = layer_1[1212] & ~layer_1[750]; 
    assign out[908] = layer_1[653] & ~layer_1[938]; 
    assign out[909] = layer_1[1212] & ~layer_1[441]; 
    assign out[910] = ~(layer_1[771] & layer_1[352]); 
    assign out[911] = ~(layer_1[871] & layer_1[242]); 
    assign out[912] = ~layer_1[1195]; 
    assign out[913] = ~(layer_1[837] & layer_1[439]); 
    assign out[914] = ~layer_1[879]; 
    assign out[915] = ~layer_1[419]; 
    assign out[916] = ~layer_1[879] | (layer_1[788] & layer_1[879]); 
    assign out[917] = ~layer_1[1195]; 
    assign out[918] = ~(layer_1[1002] & layer_1[965]); 
    assign out[919] = ~layer_1[1002]; 
    assign out[920] = ~(layer_1[447] & layer_1[242]); 
    assign out[921] = ~layer_1[1195]; 
    assign out[922] = ~layer_1[1103]; 
    assign out[923] = ~(layer_1[191] & layer_1[837]); 
    assign out[924] = ~layer_1[1103]; 
    assign out[925] = ~(layer_1[1103] | layer_1[1103]); 
    assign out[926] = ~layer_1[1103]; 
    assign out[927] = ~(layer_1[943] & layer_1[1057]); 
    assign out[928] = ~layer_1[1195]; 
    assign out[929] = ~(layer_1[205] | layer_1[903]); 
    assign out[930] = ~layer_1[943]; 
    assign out[931] = ~layer_1[879]; 
    assign out[932] = ~(layer_1[1230] & layer_1[1002]); 
    assign out[933] = ~layer_1[1230] | (layer_1[1038] & layer_1[1230]); 
    assign out[934] = ~(layer_1[1036] | layer_1[879]); 
    assign out[935] = ~(layer_1[1002] & layer_1[126]); 
    assign out[936] = ~(layer_1[466] | layer_1[205]); 
    assign out[937] = ~(layer_1[1020] & layer_1[461]); 
    assign out[938] = ~layer_1[1195]; 
    assign out[939] = ~layer_1[1103]; 
    assign out[940] = ~(layer_1[710] | layer_1[1048]); 
    assign out[941] = ~(layer_1[1036] | layer_1[461]); 
    assign out[942] = ~(layer_1[124] | layer_1[114]); 
    assign out[943] = ~(layer_1[447] & layer_1[983]); 
    assign out[944] = ~layer_1[1195]; 
    assign out[945] = ~layer_1[1103]; 
    assign out[946] = ~(layer_1[989] & layer_1[1002]); 
    assign out[947] = ~(layer_1[742] & layer_1[352]); 
    assign out[948] = ~layer_1[879]; 
    assign out[949] = ~(layer_1[1002] & layer_1[75]); 
    assign out[950] = ~layer_1[943]; 
    assign out[951] = ~(layer_1[837] & layer_1[1193]); 
    assign out[952] = ~(layer_1[461] & layer_1[123]); 
    assign out[953] = ~(layer_1[1195] & layer_1[1162]); 
    assign out[954] = ~layer_1[1103]; 
    assign out[955] = ~layer_1[205]; 
    assign out[956] = ~(layer_1[952] & layer_1[352]); 
    assign out[957] = ~(layer_1[1195] & layer_1[983]); 
    assign out[958] = ~layer_1[943]; 
    assign out[959] = ~layer_1[1195]; 
    assign out[960] = ~(layer_1[965] & layer_1[994]); 
    assign out[961] = ~(layer_1[965] & layer_1[1193]); 
    assign out[962] = ~(layer_1[1103] | layer_1[124]); 
    assign out[963] = ~(layer_1[1002] & layer_1[1230]); 
    assign out[964] = ~layer_1[1195]; 
    assign out[965] = ~(layer_1[879] | layer_1[943]); 
    assign out[966] = ~layer_1[1103]; 
    assign out[967] = ~layer_1[1195]; 
    assign out[968] = ~layer_1[943]; 
    assign out[969] = ~(layer_1[945] | layer_1[450]); 
    assign out[970] = ~(layer_1[1103] | layer_1[205]); 
    assign out[971] = ~(layer_1[983] & layer_1[38]); 
    assign out[972] = ~(layer_1[879] | layer_1[450]); 
    assign out[973] = ~layer_1[745]; 
    assign out[974] = ~layer_1[745]; 
    assign out[975] = ~(layer_1[318] & layer_1[952]); 
    assign out[976] = ~(layer_1[1002] & layer_1[983]); 
    assign out[977] = ~layer_1[18]; 
    assign out[978] = ~(layer_1[376] & layer_1[571]); 
    assign out[979] = ~(layer_1[62] | layer_1[965]); 
    assign out[980] = ~layer_1[1103]; 
    assign out[981] = ~layer_1[1002]; 
    assign out[982] = ~(layer_1[726] & layer_1[593]); 
    assign out[983] = ~(layer_1[1103] | layer_1[1103]); 
    assign out[984] = ~layer_1[879]; 
    assign out[985] = ~layer_1[1103]; 
    assign out[986] = ~layer_1[879]; 
    assign out[987] = ~layer_1[1195]; 
    assign out[988] = ~(layer_1[38] & layer_1[1002]); 
    assign out[989] = ~(layer_1[1036] | layer_1[121]); 
    assign out[990] = ~layer_1[879]; 
    assign out[991] = ~layer_1[1195]; 
    assign out[992] = ~(layer_1[75] & layer_1[1002]); 
    assign out[993] = ~(layer_1[191] & layer_1[38]); 
    assign out[994] = ~layer_1[1103]; 
    assign out[995] = ~layer_1[943]; 
    assign out[996] = ~layer_1[1230] | (layer_1[1230] & layer_1[1277]); 
    assign out[997] = ~layer_1[1195]; 
    assign out[998] = ~layer_1[943]; 
    assign out[999] = ~layer_1[1103]; 
    assign out[1000] = ~layer_1[1195]; 
    assign out[1001] = ~(layer_1[352] & layer_1[983]); 
    assign out[1002] = ~(layer_1[1002] & layer_1[447]); 
    assign out[1003] = ~(layer_1[461] & layer_1[352]); 
    assign out[1004] = ~layer_1[943]; 
    assign out[1005] = ~(layer_1[124] | layer_1[121]); 
    assign out[1006] = ~(layer_1[1002] & layer_1[983]); 
    assign out[1007] = ~(layer_1[1002] & layer_1[983]); 
    assign out[1008] = ~layer_1[1195]; 
    assign out[1009] = ~layer_1[1103]; 
    assign out[1010] = ~layer_1[1103]; 
    assign out[1011] = ~(layer_1[193] | layer_1[1195]); 
    assign out[1012] = ~(layer_1[965] & layer_1[191]); 
    assign out[1013] = ~(layer_1[742] & layer_1[1002]); 
    assign out[1014] = ~(layer_1[726] & layer_1[965]); 
    assign out[1015] = ~(layer_1[879] | layer_1[308]); 
    assign out[1016] = ~(layer_1[1103] | layer_1[943]); 
    assign out[1017] = ~(layer_1[983] & layer_1[994]); 
    assign out[1018] = ~(layer_1[447] & layer_1[983]); 
    assign out[1019] = ~(layer_1[879] | layer_1[158]); 
    assign out[1020] = ~(layer_1[975] & layer_1[1057]); 
    assign out[1021] = ~layer_1[943]; 
    assign out[1022] = ~(layer_1[541] | layer_1[1103]); 
    assign out[1023] = ~layer_1[1103]; 
    assign out[1024] = ~(layer_1[1002] & layer_1[983]); 
    assign out[1025] = ~(layer_1[551] & layer_1[1057]); 
    assign out[1026] = ~(layer_1[1002] & layer_1[983]); 
    assign out[1027] = ~(layer_1[1195] | layer_1[997]); 
    assign out[1028] = ~layer_1[943]; 
    assign out[1029] = ~layer_1[1195]; 
    assign out[1030] = ~(layer_1[1193] & layer_1[952]); 
    assign out[1031] = ~layer_1[943]; 
    assign out[1032] = ~layer_1[1103]; 
    assign out[1033] = ~(layer_1[879] & layer_1[1002]); 
    assign out[1034] = ~(layer_1[742] & layer_1[447]); 
    assign out[1035] = ~(layer_1[762] & layer_1[352]); 
    assign out[1036] = ~layer_1[879]; 
    assign out[1037] = ~layer_1[1195]; 
    assign out[1038] = ~(layer_1[1137] & layer_1[983]); 
    assign out[1039] = ~layer_1[879]; 
    assign out[1040] = layer_1[577] & ~layer_1[789]; 
    assign out[1041] = layer_1[81] ^ layer_1[64]; 
    assign out[1042] = layer_1[1271] & ~layer_1[626]; 
    assign out[1043] = layer_1[181] ^ layer_1[746]; 
    assign out[1044] = layer_1[332] & ~layer_1[626]; 
    assign out[1045] = layer_1[1105] ^ layer_1[112]; 
    assign out[1046] = layer_1[758] | layer_1[858]; 
    assign out[1047] = ~layer_1[626]; 
    assign out[1048] = layer_1[291] ^ layer_1[3]; 
    assign out[1049] = layer_1[147] & ~layer_1[518]; 
    assign out[1050] = layer_1[301]; 
    assign out[1051] = layer_1[1271] ^ layer_1[25]; 
    assign out[1052] = layer_1[529] ^ layer_1[550]; 
    assign out[1053] = layer_1[81] ^ layer_1[476]; 
    assign out[1054] = layer_1[81]; 
    assign out[1055] = layer_1[153] ^ layer_1[378]; 
    assign out[1056] = layer_1[758]; 
    assign out[1057] = layer_1[1026] ^ layer_1[467]; 
    assign out[1058] = layer_1[905] ^ layer_1[892]; 
    assign out[1059] = layer_1[960] | layer_1[858]; 
    assign out[1060] = layer_1[770] | layer_1[581]; 
    assign out[1061] = layer_1[64] ^ layer_1[81]; 
    assign out[1062] = layer_1[58]; 
    assign out[1063] = layer_1[858]; 
    assign out[1064] = layer_1[9] ^ layer_1[81]; 
    assign out[1065] = layer_1[64] ^ layer_1[81]; 
    assign out[1066] = layer_1[1064] & ~layer_1[931]; 
    assign out[1067] = layer_1[147] ^ layer_1[1257]; 
    assign out[1068] = layer_1[58] | layer_1[858]; 
    assign out[1069] = layer_1[706] & ~layer_1[1026]; 
    assign out[1070] = ~layer_1[1054]; 
    assign out[1071] = layer_1[892] ^ layer_1[905]; 
    assign out[1072] = layer_1[428] ^ layer_1[658]; 
    assign out[1073] = layer_1[577] ^ layer_1[550]; 
    assign out[1074] = layer_1[550] ^ layer_1[577]; 
    assign out[1075] = layer_1[529] ^ layer_1[550]; 
    assign out[1076] = layer_1[322] ^ layer_1[1221]; 
    assign out[1077] = ~(layer_1[955] & layer_1[1200]); 
    assign out[1078] = layer_1[404] & ~layer_1[626]; 
    assign out[1079] = layer_1[301]; 
    assign out[1080] = layer_1[237] ^ layer_1[77]; 
    assign out[1081] = layer_1[847] ^ layer_1[81]; 
    assign out[1082] = layer_1[813] ^ layer_1[605]; 
    assign out[1083] = ~(layer_1[914] & layer_1[889]); 
    assign out[1084] = layer_1[81] & ~layer_1[587]; 
    assign out[1085] = layer_1[997] ^ layer_1[81]; 
    assign out[1086] = layer_1[1271] ^ layer_1[857]; 
    assign out[1087] = layer_1[81] ^ layer_1[64]; 
    assign out[1088] = layer_1[565] ^ layer_1[322]; 
    assign out[1089] = layer_1[213] ^ layer_1[758]; 
    assign out[1090] = layer_1[1064] & ~layer_1[362]; 
    assign out[1091] = layer_1[647] | layer_1[1196]; 
    assign out[1092] = layer_1[9] ^ layer_1[81]; 
    assign out[1093] = layer_1[416] ^ layer_1[1271]; 
    assign out[1094] = layer_1[931] ^ layer_1[499]; 
    assign out[1095] = layer_1[872] & ~layer_1[816]; 
    assign out[1096] = layer_1[81] ^ layer_1[565]; 
    assign out[1097] = ~(layer_1[64] | layer_1[857]); 
    assign out[1098] = layer_1[428] ^ layer_1[81]; 
    assign out[1099] = layer_1[58] | layer_1[858]; 
    assign out[1100] = layer_1[1271] ^ layer_1[416]; 
    assign out[1101] = layer_1[175] ^ layer_1[189]; 
    assign out[1102] = layer_1[626] ^ layer_1[767]; 
    assign out[1103] = layer_1[469] & ~layer_1[362]; 
    assign out[1104] = layer_1[813] ^ layer_1[81]; 
    assign out[1105] = layer_1[467] ^ layer_1[857]; 
    assign out[1106] = layer_1[64] ^ layer_1[831]; 
    assign out[1107] = layer_1[147] & ~layer_1[1026]; 
    assign out[1108] = layer_1[1276] & ~layer_1[416]; 
    assign out[1109] = layer_1[931] ^ layer_1[81]; 
    assign out[1110] = layer_1[110] ^ layer_1[346]; 
    assign out[1111] = layer_1[1271] & ~layer_1[626]; 
    assign out[1112] = layer_1[967] ^ layer_1[109]; 
    assign out[1113] = layer_1[550] ^ layer_1[81]; 
    assign out[1114] = ~(layer_1[682] & layer_1[955]); 
    assign out[1115] = layer_1[147] ^ layer_1[626]; 
    assign out[1116] = layer_1[322] & ~layer_1[1221]; 
    assign out[1117] = layer_1[958] & ~layer_1[857]; 
    assign out[1118] = layer_1[1253] ^ layer_1[291]; 
    assign out[1119] = layer_1[416] ^ layer_1[1276]; 
    assign out[1120] = layer_1[980] ^ layer_1[787]; 
    assign out[1121] = ~(layer_1[1026] & layer_1[553]); 
    assign out[1122] = layer_1[58] & ~layer_1[980]; 
    assign out[1123] = layer_1[858] | layer_1[58]; 
    assign out[1124] = layer_1[813] ^ layer_1[81]; 
    assign out[1125] = layer_1[81] ^ layer_1[813]; 
    assign out[1126] = layer_1[587] ^ layer_1[81]; 
    assign out[1127] = layer_1[64] ^ layer_1[81]; 
    assign out[1128] = layer_1[1271] ^ layer_1[321]; 
    assign out[1129] = layer_1[81] ^ layer_1[64]; 
    assign out[1130] = layer_1[109] ^ layer_1[1127]; 
    assign out[1131] = layer_1[378] ^ layer_1[1237]; 
    assign out[1132] = layer_1[811] ^ layer_1[64]; 
    assign out[1133] = layer_1[313] ^ layer_1[813]; 
    assign out[1134] = layer_1[813] ^ layer_1[81]; 
    assign out[1135] = ~(layer_1[349] & layer_1[1200]); 
    assign out[1136] = layer_1[813] ^ layer_1[1223]; 
    assign out[1137] = layer_1[81] ^ layer_1[1016]; 
    assign out[1138] = ~layer_1[645]; 
    assign out[1139] = layer_1[147]; 
    assign out[1140] = layer_1[967] ^ layer_1[109]; 
    assign out[1141] = layer_1[266] ^ layer_1[869]; 
    assign out[1142] = layer_1[1209] ^ layer_1[605]; 
    assign out[1143] = layer_1[291] ^ layer_1[1253]; 
    assign out[1144] = layer_1[235] ^ layer_1[84]; 
    assign out[1145] = layer_1[858] | layer_1[58]; 
    assign out[1146] = layer_1[1175] & ~layer_1[64]; 
    assign out[1147] = layer_1[301]; 
    assign out[1148] = layer_1[858] | layer_1[1165]; 
    assign out[1149] = layer_1[64] ^ layer_1[301]; 
    assign out[1150] = layer_1[550] ^ layer_1[566]; 
    assign out[1151] = layer_1[967] ^ layer_1[109]; 
    assign out[1152] = layer_1[1271] ^ layer_1[813]; 
    assign out[1153] = layer_1[81] ^ layer_1[64]; 
    assign out[1154] = layer_1[658] ^ layer_1[869]; 
    assign out[1155] = layer_1[278] ^ layer_1[1196]; 
    assign out[1156] = layer_1[64] ^ layer_1[81]; 
    assign out[1157] = ~layer_1[914]; 
    assign out[1158] = layer_1[58] | layer_1[858]; 
    assign out[1159] = layer_1[147] & ~layer_1[212]; 
    assign out[1160] = layer_1[746] ^ layer_1[587]; 
    assign out[1161] = layer_1[109] ^ layer_1[967]; 
    assign out[1162] = layer_1[1196] ^ layer_1[1139]; 
    assign out[1163] = layer_1[531] ^ layer_1[339]; 
    assign out[1164] = layer_1[84] ^ layer_1[892]; 
    assign out[1165] = layer_1[733] ^ layer_1[1237]; 
    assign out[1166] = ~layer_1[626]; 
    assign out[1167] = layer_1[278] ^ layer_1[1196]; 
    assign out[1168] = layer_1[321] ^ layer_1[1271]; 
    assign out[1169] = layer_1[921] & ~layer_1[564]; 
    assign out[1170] = ~(layer_1[598] | layer_1[648]); 
    assign out[1171] = ~(layer_1[598] | layer_1[943]); 
    assign out[1172] = ~(layer_1[50] | layer_1[139]); 
    assign out[1173] = ~(layer_1[598] | layer_1[50]); 
    assign out[1174] = ~(layer_1[887] | layer_1[648]); 
    assign out[1175] = ~(layer_1[590] | layer_1[1005]); 
    assign out[1176] = ~(layer_1[1005] | layer_1[139]); 
    assign out[1177] = ~layer_1[648]; 
    assign out[1178] = ~(layer_1[22] | layer_1[289]); 
    assign out[1179] = layer_1[290] & ~layer_1[943]; 
    assign out[1180] = ~(layer_1[943] | layer_1[943]); 
    assign out[1181] = ~(layer_1[22] | layer_1[598]); 
    assign out[1182] = ~(layer_1[590] | layer_1[22]); 
    assign out[1183] = layer_1[742] & ~layer_1[904]; 
    assign out[1184] = ~(layer_1[943] | layer_1[453]); 
    assign out[1185] = layer_1[275] & ~layer_1[22]; 
    assign out[1186] = layer_1[553] ^ layer_1[700]; 
    assign out[1187] = ~(layer_1[598] | layer_1[590]); 
    assign out[1188] = ~layer_1[598]; 
    assign out[1189] = ~layer_1[598]; 
    assign out[1190] = layer_1[742] & ~layer_1[22]; 
    assign out[1191] = layer_1[1194] ^ layer_1[436]; 
    assign out[1192] = ~(layer_1[648] | layer_1[50]); 
    assign out[1193] = ~layer_1[598]; 
    assign out[1194] = ~layer_1[22]; 
    assign out[1195] = layer_1[742] & ~layer_1[598]; 
    assign out[1196] = ~layer_1[648]; 
    assign out[1197] = ~(layer_1[904] | layer_1[4]); 
    assign out[1198] = ~layer_1[598]; 
    assign out[1199] = ~(layer_1[943] | layer_1[446]); 
    assign out[1200] = ~(layer_1[598] | layer_1[139]); 
    assign out[1201] = layer_1[551] ^ layer_1[439]; 
    assign out[1202] = ~(layer_1[22] | layer_1[598]); 
    assign out[1203] = ~(layer_1[943] | layer_1[598]); 
    assign out[1204] = ~(layer_1[1289] | layer_1[648]); 
    assign out[1205] = ~(layer_1[598] | layer_1[887]); 
    assign out[1206] = ~(layer_1[453] | layer_1[598]); 
    assign out[1207] = ~layer_1[598]; 
    assign out[1208] = ~(layer_1[887] | layer_1[305]); 
    assign out[1209] = ~(layer_1[139] | layer_1[495]); 
    assign out[1210] = ~(layer_1[50] | layer_1[329]); 
    assign out[1211] = ~(layer_1[943] | layer_1[598]); 
    assign out[1212] = layer_1[898] & ~layer_1[810]; 
    assign out[1213] = ~(layer_1[598] | layer_1[648]); 
    assign out[1214] = layer_1[944] ^ layer_1[742]; 
    assign out[1215] = layer_1[983] & ~layer_1[943]; 
    assign out[1216] = ~layer_1[139]; 
    assign out[1217] = ~(layer_1[129] | layer_1[810]); 
    assign out[1218] = ~(layer_1[279] & layer_1[191]); 
    assign out[1219] = ~(layer_1[50] | layer_1[700]); 
    assign out[1220] = ~(layer_1[22] | layer_1[700]); 
    assign out[1221] = ~layer_1[279]; 
    assign out[1222] = ~(layer_1[887] | layer_1[590]); 
    assign out[1223] = ~(layer_1[139] | layer_1[50]); 
    assign out[1224] = ~(layer_1[1208] & layer_1[887]); 
    assign out[1225] = ~(layer_1[598] | layer_1[842]); 
    assign out[1226] = ~(layer_1[810] | layer_1[139]); 
    assign out[1227] = layer_1[383] & ~layer_1[160]; 
    assign out[1228] = ~(layer_1[50] | layer_1[139]); 
    assign out[1229] = ~(layer_1[139] | layer_1[598]); 
    assign out[1230] = ~(layer_1[598] | layer_1[1225]); 
    assign out[1231] = ~layer_1[887]; 
    assign out[1232] = ~(layer_1[648] | layer_1[22]); 
    assign out[1233] = ~(layer_1[598] | layer_1[139]); 
    assign out[1234] = ~(layer_1[590] | layer_1[887]); 
    assign out[1235] = ~layer_1[139]; 
    assign out[1236] = ~(layer_1[886] | layer_1[139]); 
    assign out[1237] = ~layer_1[598]; 
    assign out[1238] = ~(layer_1[139] | layer_1[886]); 
    assign out[1239] = ~layer_1[598]; 
    assign out[1240] = ~(layer_1[598] | layer_1[139]); 
    assign out[1241] = layer_1[983] & ~layer_1[837]; 
    assign out[1242] = layer_1[460] & ~layer_1[598]; 
    assign out[1243] = layer_1[943] ^ layer_1[983]; 
    assign out[1244] = ~(layer_1[598] | layer_1[598]); 
    assign out[1245] = ~(layer_1[577] | layer_1[50]); 
    assign out[1246] = ~(layer_1[810] | layer_1[598]); 
    assign out[1247] = layer_1[742] & ~layer_1[22]; 
    assign out[1248] = ~(layer_1[590] | layer_1[648]); 
    assign out[1249] = layer_1[837] ^ layer_1[372]; 
    assign out[1250] = ~layer_1[887]; 
    assign out[1251] = ~(layer_1[598] | layer_1[598]); 
    assign out[1252] = ~(layer_1[873] | layer_1[590]); 
    assign out[1253] = ~layer_1[598]; 
    assign out[1254] = layer_1[742] & ~layer_1[598]; 
    assign out[1255] = ~(layer_1[139] | layer_1[50]); 
    assign out[1256] = ~(layer_1[22] | layer_1[495]); 
    assign out[1257] = ~(layer_1[598] | layer_1[1069]); 
    assign out[1258] = ~(layer_1[50] | layer_1[139]); 
    assign out[1259] = ~(layer_1[139] | layer_1[598]); 
    assign out[1260] = ~(layer_1[648] | layer_1[22]); 
    assign out[1261] = ~(layer_1[904] & layer_1[18]); 
    assign out[1262] = layer_1[1002] & ~layer_1[22]; 
    assign out[1263] = layer_1[837] ^ layer_1[1230]; 
    assign out[1264] = layer_1[297] & ~layer_1[598]; 
    assign out[1265] = ~(layer_1[886] | layer_1[810]); 
    assign out[1266] = ~layer_1[887]; 
    assign out[1267] = ~(layer_1[598] | layer_1[648]); 
    assign out[1268] = layer_1[983] & ~layer_1[22]; 
    assign out[1269] = ~layer_1[422]; 
    assign out[1270] = ~(layer_1[598] | layer_1[887]); 
    assign out[1271] = ~(layer_1[216] | layer_1[160]); 
    assign out[1272] = ~layer_1[598]; 
    assign out[1273] = ~(layer_1[887] & layer_1[279]); 
    assign out[1274] = ~layer_1[887]; 
    assign out[1275] = ~layer_1[648]; 
    assign out[1276] = ~(layer_1[590] | layer_1[598]); 
    assign out[1277] = ~(layer_1[50] | layer_1[598]); 
    assign out[1278] = layer_1[916] ^ layer_1[1271]; 
    assign out[1279] = ~(layer_1[598] | layer_1[801]); 
    assign out[1280] = ~(layer_1[22] | layer_1[598]); 
    assign out[1281] = ~(layer_1[289] | layer_1[887]); 
    assign out[1282] = ~(layer_1[598] | layer_1[22]); 
    assign out[1283] = ~(layer_1[139] | layer_1[50]); 
    assign out[1284] = ~(layer_1[139] | layer_1[27]); 
    assign out[1285] = ~layer_1[648] | (layer_1[1191] & layer_1[648]); 
    assign out[1286] = ~(layer_1[648] | layer_1[673]); 
    assign out[1287] = ~layer_1[887]; 
    assign out[1288] = ~(layer_1[648] | layer_1[1256]); 
    assign out[1289] = layer_1[297] & ~layer_1[598]; 
    assign out[1290] = ~(layer_1[139] | layer_1[50]); 
    assign out[1291] = ~(layer_1[50] | layer_1[700]); 
    assign out[1292] = ~(layer_1[943] | layer_1[648]); 
    assign out[1293] = ~(layer_1[50] | layer_1[139]); 
    assign out[1294] = ~layer_1[139]; 
    assign out[1295] = layer_1[848] ^ layer_1[879]; 
    assign out[1296] = ~(layer_1[887] | layer_1[305]); 
    assign out[1297] = ~(layer_1[191] & layer_1[1208]); 
    assign out[1298] = ~(layer_1[943] | layer_1[732]); 
    assign out[1299] = ~(layer_1[50] | layer_1[302]); 
    // Arrange outputs in categories ================================================
    assign categories[129:0] = out[129:0];
    assign categories[254:130] = 0;
    assign categories[384:255] = out[259:130];
    assign categories[509:385] = 0;
    assign categories[639:510] = out[389:260];
    assign categories[764:640] = 0;
    assign categories[894:765] = out[519:390];
    assign categories[1019:895] = 0;
    assign categories[1149:1020] = out[649:520];
    assign categories[1274:1150] = 0;
    assign categories[1404:1275] = out[779:650];
    assign categories[1529:1405] = 0;
    assign categories[1659:1530] = out[909:780];
    assign categories[1784:1660] = 0;
    assign categories[1914:1785] = out[1039:910];
    assign categories[2039:1915] = 0;
    assign categories[2169:2040] = out[1169:1040];
    assign categories[2294:2170] = 0;
    assign categories[2424:2295] = out[1299:1170];
    assign categories[2549:2425] = 0;

endmodule
