// Generated from: baralizm_20250116-123948_acc9424_seed1022128_epochs50_dsp128_3x4000_b256_lrm5-1with_dataset.npz
module net (
    input wire  [255:0] in,
    output wire [3999:0] out
);
    wire [4000:0] layer_0;
    wire [4000:0] layer_1;

    // Layer 0 ============================================================
    assign layer_0[0] = ~in[248] | (in[234] & in[248]); 
    assign layer_0[1] = ~(in[194] | in[191]); 
    assign layer_0[2] = ~in[142] | (in[253] & in[142]); 
    assign layer_0[3] = in[231]; 
    assign layer_0[4] = in[73] & ~in[110]; 
    assign layer_0[5] = ~in[107]; 
    assign layer_0[6] = ~in[212] | (in[228] & in[212]); 
    assign layer_0[7] = in[60] | in[164]; 
    assign layer_0[8] = ~in[13]; 
    assign layer_0[9] = in[248]; 
    assign layer_0[10] = ~(in[1] | in[115]); 
    assign layer_0[11] = in[69] & ~in[132]; 
    assign layer_0[12] = in[141] & ~in[35]; 
    assign layer_0[13] = in[155] | in[28]; 
    assign layer_0[14] = in[183] & ~in[211]; 
    assign layer_0[15] = ~in[89] | (in[89] & in[17]); 
    assign layer_0[16] = in[127]; 
    assign layer_0[17] = ~in[137] | (in[128] & in[137]); 
    assign layer_0[18] = in[49] ^ in[149]; 
    assign layer_0[19] = ~in[107]; 
    assign layer_0[20] = ~(in[23] ^ in[20]); 
    assign layer_0[21] = ~in[148]; 
    assign layer_0[22] = in[204] ^ in[172]; 
    assign layer_0[23] = in[35]; 
    assign layer_0[24] = in[56] & ~in[140]; 
    assign layer_0[25] = ~in[165] | (in[176] & in[165]); 
    assign layer_0[26] = in[166] ^ in[228]; 
    assign layer_0[27] = ~in[165] | (in[225] & in[165]); 
    assign layer_0[28] = ~in[199]; 
    assign layer_0[29] = ~(in[183] & in[120]); 
    assign layer_0[30] = in[170] & in[180]; 
    assign layer_0[31] = in[17] ^ in[94]; 
    assign layer_0[32] = in[118]; 
    assign layer_0[33] = ~in[76]; 
    assign layer_0[34] = ~in[143] | (in[143] & in[135]); 
    assign layer_0[35] = ~in[73] | (in[13] & in[73]); 
    assign layer_0[36] = in[166] & ~in[195]; 
    assign layer_0[37] = ~in[190]; 
    assign layer_0[38] = in[168] & ~in[74]; 
    assign layer_0[39] = ~in[196] | (in[196] & in[98]); 
    assign layer_0[40] = ~(in[214] ^ in[199]); 
    assign layer_0[41] = in[230] ^ in[210]; 
    assign layer_0[42] = in[24] & ~in[17]; 
    assign layer_0[43] = ~in[217]; 
    assign layer_0[44] = in[70] | in[28]; 
    assign layer_0[45] = in[210]; 
    assign layer_0[46] = ~in[74]; 
    assign layer_0[47] = ~(in[106] ^ in[117]); 
    assign layer_0[48] = in[68] | in[60]; 
    assign layer_0[49] = ~in[173]; 
    assign layer_0[50] = in[135]; 
    assign layer_0[51] = in[149] & ~in[49]; 
    assign layer_0[52] = in[48] ^ in[130]; 
    assign layer_0[53] = ~(in[47] | in[76]); 
    assign layer_0[54] = ~(in[194] & in[213]); 
    assign layer_0[55] = in[144] & in[60]; 
    assign layer_0[56] = ~(in[8] | in[110]); 
    assign layer_0[57] = in[222] | in[195]; 
    assign layer_0[58] = ~(in[249] ^ in[220]); 
    assign layer_0[59] = ~(in[195] ^ in[250]); 
    assign layer_0[60] = in[226] | in[253]; 
    assign layer_0[61] = ~in[236]; 
    assign layer_0[62] = ~(in[80] | in[7]); 
    assign layer_0[63] = in[18] & in[145]; 
    assign layer_0[64] = in[18] | in[44]; 
    assign layer_0[65] = ~in[148] | (in[193] & in[148]); 
    assign layer_0[66] = in[78] ^ in[112]; 
    assign layer_0[67] = in[255]; 
    assign layer_0[68] = ~in[131] | (in[110] & in[131]); 
    assign layer_0[69] = in[26]; 
    assign layer_0[70] = in[224] & in[148]; 
    assign layer_0[71] = ~(in[124] ^ in[71]); 
    assign layer_0[72] = ~(in[202] ^ in[208]); 
    assign layer_0[73] = in[165] & ~in[79]; 
    assign layer_0[74] = in[240]; 
    assign layer_0[75] = ~(in[80] | in[155]); 
    assign layer_0[76] = in[210]; 
    assign layer_0[77] = ~in[26]; 
    assign layer_0[78] = in[30]; 
    assign layer_0[79] = in[149] & ~in[95]; 
    assign layer_0[80] = in[22] & ~in[11]; 
    assign layer_0[81] = ~in[134] | (in[134] & in[220]); 
    assign layer_0[82] = ~in[8] | (in[8] & in[111]); 
    assign layer_0[83] = ~in[139]; 
    assign layer_0[84] = ~in[75] | (in[17] & in[75]); 
    assign layer_0[85] = in[151] & in[43]; 
    assign layer_0[86] = in[152] & ~in[178]; 
    assign layer_0[87] = in[73]; 
    assign layer_0[88] = ~in[40] | (in[40] & in[114]); 
    assign layer_0[89] = in[88] ^ in[156]; 
    assign layer_0[90] = in[86] & ~in[186]; 
    assign layer_0[91] = in[34] & ~in[11]; 
    assign layer_0[92] = in[126] | in[163]; 
    assign layer_0[93] = in[21] | in[121]; 
    assign layer_0[94] = ~in[58] | (in[58] & in[44]); 
    assign layer_0[95] = in[88] & ~in[140]; 
    assign layer_0[96] = in[80] | in[187]; 
    assign layer_0[97] = ~(in[27] ^ in[26]); 
    assign layer_0[98] = ~(in[84] | in[56]); 
    assign layer_0[99] = in[253] ^ in[174]; 
    assign layer_0[100] = ~in[57]; 
    assign layer_0[101] = ~in[10]; 
    assign layer_0[102] = in[88] & ~in[29]; 
    assign layer_0[103] = ~(in[96] | in[64]); 
    assign layer_0[104] = ~(in[103] ^ in[157]); 
    assign layer_0[105] = ~(in[53] & in[8]); 
    assign layer_0[106] = in[44]; 
    assign layer_0[107] = in[116] & ~in[228]; 
    assign layer_0[108] = ~(in[46] | in[104]); 
    assign layer_0[109] = ~(in[255] | in[214]); 
    assign layer_0[110] = in[68]; 
    assign layer_0[111] = ~(in[37] | in[34]); 
    assign layer_0[112] = in[131] | in[185]; 
    assign layer_0[113] = ~in[96] | (in[96] & in[98]); 
    assign layer_0[114] = in[222] | in[190]; 
    assign layer_0[115] = in[247] ^ in[178]; 
    assign layer_0[116] = ~in[171] | (in[171] & in[246]); 
    assign layer_0[117] = in[185] ^ in[234]; 
    assign layer_0[118] = in[86] & ~in[161]; 
    assign layer_0[119] = in[119] ^ in[246]; 
    assign layer_0[120] = in[186] & in[100]; 
    assign layer_0[121] = ~(in[52] ^ in[141]); 
    assign layer_0[122] = in[170] | in[111]; 
    assign layer_0[123] = in[192] & ~in[129]; 
    assign layer_0[124] = ~in[164]; 
    assign layer_0[125] = ~(in[42] | in[155]); 
    assign layer_0[126] = ~(in[180] & in[151]); 
    assign layer_0[127] = ~(in[177] ^ in[181]); 
    assign layer_0[128] = ~in[216]; 
    assign layer_0[129] = ~in[78] | (in[78] & in[127]); 
    assign layer_0[130] = in[104] & ~in[190]; 
    assign layer_0[131] = ~in[196]; 
    assign layer_0[132] = in[119] & ~in[147]; 
    assign layer_0[133] = in[94] & ~in[212]; 
    assign layer_0[134] = in[54] & ~in[81]; 
    assign layer_0[135] = ~in[106] | (in[210] & in[106]); 
    assign layer_0[136] = in[167] ^ in[113]; 
    assign layer_0[137] = ~(in[0] ^ in[122]); 
    assign layer_0[138] = ~(in[198] ^ in[143]); 
    assign layer_0[139] = in[177] ^ in[217]; 
    assign layer_0[140] = in[154] & ~in[30]; 
    assign layer_0[141] = ~in[135] | (in[135] & in[225]); 
    assign layer_0[142] = in[131]; 
    assign layer_0[143] = ~(in[0] | in[72]); 
    assign layer_0[144] = in[64] & ~in[182]; 
    assign layer_0[145] = ~in[166] | (in[80] & in[166]); 
    assign layer_0[146] = ~in[39]; 
    assign layer_0[147] = in[35] | in[109]; 
    assign layer_0[148] = in[59] & ~in[127]; 
    assign layer_0[149] = ~in[1]; 
    assign layer_0[150] = ~in[126] | (in[221] & in[126]); 
    assign layer_0[151] = ~(in[1] | in[36]); 
    assign layer_0[152] = in[137] & ~in[23]; 
    assign layer_0[153] = in[204] | in[188]; 
    assign layer_0[154] = ~(in[103] | in[231]); 
    assign layer_0[155] = ~(in[164] ^ in[223]); 
    assign layer_0[156] = ~in[236] | (in[140] & in[236]); 
    assign layer_0[157] = in[140]; 
    assign layer_0[158] = ~in[134] | (in[35] & in[134]); 
    assign layer_0[159] = ~in[91] | (in[15] & in[91]); 
    assign layer_0[160] = ~in[253]; 
    assign layer_0[161] = ~(in[137] ^ in[159]); 
    assign layer_0[162] = ~in[165] | (in[98] & in[165]); 
    assign layer_0[163] = in[156] | in[207]; 
    assign layer_0[164] = ~in[127] | (in[142] & in[127]); 
    assign layer_0[165] = ~(in[76] | in[91]); 
    assign layer_0[166] = in[91]; 
    assign layer_0[167] = ~in[70] | (in[70] & in[58]); 
    assign layer_0[168] = in[118]; 
    assign layer_0[169] = in[16] & ~in[31]; 
    assign layer_0[170] = in[145]; 
    assign layer_0[171] = ~(in[17] & in[83]); 
    assign layer_0[172] = ~(in[111] | in[78]); 
    assign layer_0[173] = ~(in[17] & in[14]); 
    assign layer_0[174] = in[80]; 
    assign layer_0[175] = in[178] & ~in[99]; 
    assign layer_0[176] = in[195]; 
    assign layer_0[177] = ~(in[99] & in[87]); 
    assign layer_0[178] = in[195] | in[222]; 
    assign layer_0[179] = ~(in[83] | in[144]); 
    assign layer_0[180] = in[170]; 
    assign layer_0[181] = in[165]; 
    assign layer_0[182] = in[198]; 
    assign layer_0[183] = in[103]; 
    assign layer_0[184] = ~(in[129] | in[243]); 
    assign layer_0[185] = in[151]; 
    assign layer_0[186] = ~(in[142] | in[186]); 
    assign layer_0[187] = ~(in[41] | in[21]); 
    assign layer_0[188] = in[80] & ~in[175]; 
    assign layer_0[189] = ~in[127] | (in[127] & in[8]); 
    assign layer_0[190] = in[157] & ~in[79]; 
    assign layer_0[191] = ~(in[201] ^ in[218]); 
    assign layer_0[192] = ~in[181] | (in[181] & in[227]); 
    assign layer_0[193] = ~(in[12] ^ in[9]); 
    assign layer_0[194] = in[116] ^ in[209]; 
    assign layer_0[195] = ~in[175] | (in[242] & in[175]); 
    assign layer_0[196] = in[28] ^ in[155]; 
    assign layer_0[197] = in[21] | in[95]; 
    assign layer_0[198] = ~(in[210] | in[159]); 
    assign layer_0[199] = in[54] & in[158]; 
    assign layer_0[200] = ~in[27]; 
    assign layer_0[201] = ~in[62] | (in[142] & in[62]); 
    assign layer_0[202] = in[200] ^ in[213]; 
    assign layer_0[203] = in[131]; 
    assign layer_0[204] = in[178]; 
    assign layer_0[205] = in[232] & ~in[147]; 
    assign layer_0[206] = in[148] & ~in[207]; 
    assign layer_0[207] = in[227] | in[229]; 
    assign layer_0[208] = ~in[106] | (in[106] & in[196]); 
    assign layer_0[209] = in[103] & ~in[170]; 
    assign layer_0[210] = in[127] ^ in[80]; 
    assign layer_0[211] = in[158] & ~in[35]; 
    assign layer_0[212] = ~in[194]; 
    assign layer_0[213] = ~in[211] | (in[142] & in[211]); 
    assign layer_0[214] = in[233] ^ in[176]; 
    assign layer_0[215] = ~(in[242] ^ in[255]); 
    assign layer_0[216] = in[110] & ~in[185]; 
    assign layer_0[217] = in[175]; 
    assign layer_0[218] = ~(in[129] & in[243]); 
    assign layer_0[219] = ~(in[190] ^ in[227]); 
    assign layer_0[220] = ~in[56] | (in[56] & in[140]); 
    assign layer_0[221] = in[208] & in[144]; 
    assign layer_0[222] = ~in[101] | (in[12] & in[101]); 
    assign layer_0[223] = in[108]; 
    assign layer_0[224] = ~(in[60] ^ in[110]); 
    assign layer_0[225] = ~in[193] | (in[255] & in[193]); 
    assign layer_0[226] = in[52] & ~in[59]; 
    assign layer_0[227] = in[88] & ~in[3]; 
    assign layer_0[228] = in[68] ^ in[58]; 
    assign layer_0[229] = ~in[104]; 
    assign layer_0[230] = in[73] & ~in[118]; 
    assign layer_0[231] = ~(in[185] & in[131]); 
    assign layer_0[232] = in[114] & ~in[239]; 
    assign layer_0[233] = ~in[61]; 
    assign layer_0[234] = in[218]; 
    assign layer_0[235] = in[125]; 
    assign layer_0[236] = in[90]; 
    assign layer_0[237] = ~(in[54] ^ in[58]); 
    assign layer_0[238] = in[1] ^ in[82]; 
    assign layer_0[239] = ~(in[177] | in[225]); 
    assign layer_0[240] = in[40]; 
    assign layer_0[241] = ~in[196] | (in[196] & in[80]); 
    assign layer_0[242] = in[10] | in[95]; 
    assign layer_0[243] = in[107]; 
    assign layer_0[244] = ~in[92]; 
    assign layer_0[245] = ~in[229]; 
    assign layer_0[246] = ~in[146] | (in[146] & in[242]); 
    assign layer_0[247] = ~in[107]; 
    assign layer_0[248] = ~(in[177] ^ in[165]); 
    assign layer_0[249] = in[242] | in[209]; 
    assign layer_0[250] = in[203] | in[242]; 
    assign layer_0[251] = in[7]; 
    assign layer_0[252] = in[177]; 
    assign layer_0[253] = ~in[132]; 
    assign layer_0[254] = ~in[133] | (in[173] & in[133]); 
    assign layer_0[255] = in[48] & ~in[103]; 
    assign layer_0[256] = in[217]; 
    assign layer_0[257] = in[100] | in[126]; 
    assign layer_0[258] = in[67]; 
    assign layer_0[259] = in[224] | in[230]; 
    assign layer_0[260] = in[88] | in[176]; 
    assign layer_0[261] = in[98]; 
    assign layer_0[262] = ~(in[205] & in[175]); 
    assign layer_0[263] = in[144] | in[155]; 
    assign layer_0[264] = ~(in[32] | in[88]); 
    assign layer_0[265] = in[243] & ~in[254]; 
    assign layer_0[266] = ~in[215] | (in[215] & in[222]); 
    assign layer_0[267] = ~in[181]; 
    assign layer_0[268] = ~(in[13] | in[10]); 
    assign layer_0[269] = in[205] ^ in[78]; 
    assign layer_0[270] = in[112] & in[72]; 
    assign layer_0[271] = in[144]; 
    assign layer_0[272] = in[101] & ~in[129]; 
    assign layer_0[273] = in[49] & in[6]; 
    assign layer_0[274] = in[176] & in[51]; 
    assign layer_0[275] = ~(in[65] | in[175]); 
    assign layer_0[276] = in[109] & ~in[52]; 
    assign layer_0[277] = in[22] | in[21]; 
    assign layer_0[278] = ~in[18]; 
    assign layer_0[279] = ~in[87]; 
    assign layer_0[280] = in[16] | in[61]; 
    assign layer_0[281] = ~in[21]; 
    assign layer_0[282] = in[91] ^ in[194]; 
    assign layer_0[283] = ~(in[5] ^ in[18]); 
    assign layer_0[284] = in[189]; 
    assign layer_0[285] = ~(in[154] | in[79]); 
    assign layer_0[286] = in[204] ^ in[245]; 
    assign layer_0[287] = ~(in[92] | in[30]); 
    assign layer_0[288] = ~(in[124] ^ in[162]); 
    assign layer_0[289] = in[150] ^ in[99]; 
    assign layer_0[290] = ~(in[213] | in[112]); 
    assign layer_0[291] = in[165] ^ in[198]; 
    assign layer_0[292] = in[78] | in[195]; 
    assign layer_0[293] = ~in[54]; 
    assign layer_0[294] = in[153] & ~in[32]; 
    assign layer_0[295] = in[209] ^ in[187]; 
    assign layer_0[296] = in[128] ^ in[94]; 
    assign layer_0[297] = in[20] & in[10]; 
    assign layer_0[298] = in[62] & ~in[23]; 
    assign layer_0[299] = in[82] & ~in[58]; 
    assign layer_0[300] = ~in[168] | (in[168] & in[235]); 
    assign layer_0[301] = ~(in[87] | in[155]); 
    assign layer_0[302] = ~in[180]; 
    assign layer_0[303] = ~(in[230] ^ in[226]); 
    assign layer_0[304] = ~in[142] | (in[59] & in[142]); 
    assign layer_0[305] = ~in[118] | (in[118] & in[126]); 
    assign layer_0[306] = in[39]; 
    assign layer_0[307] = ~(in[142] | in[150]); 
    assign layer_0[308] = in[119] & ~in[140]; 
    assign layer_0[309] = ~(in[110] | in[169]); 
    assign layer_0[310] = in[73] & in[134]; 
    assign layer_0[311] = in[54] & ~in[50]; 
    assign layer_0[312] = ~(in[46] ^ in[151]); 
    assign layer_0[313] = in[113] ^ in[203]; 
    assign layer_0[314] = ~(in[80] | in[76]); 
    assign layer_0[315] = in[135] & ~in[243]; 
    assign layer_0[316] = ~in[131] | (in[205] & in[131]); 
    assign layer_0[317] = ~in[245] | (in[245] & in[160]); 
    assign layer_0[318] = ~(in[125] | in[126]); 
    assign layer_0[319] = ~(in[72] ^ in[64]); 
    assign layer_0[320] = ~(in[71] & in[181]); 
    assign layer_0[321] = in[198] | in[173]; 
    assign layer_0[322] = ~in[233]; 
    assign layer_0[323] = in[197] & ~in[206]; 
    assign layer_0[324] = in[20] | in[10]; 
    assign layer_0[325] = in[166] & ~in[210]; 
    assign layer_0[326] = in[66]; 
    assign layer_0[327] = ~(in[253] ^ in[190]); 
    assign layer_0[328] = in[106]; 
    assign layer_0[329] = in[51] & ~in[34]; 
    assign layer_0[330] = ~(in[153] & in[107]); 
    assign layer_0[331] = in[36]; 
    assign layer_0[332] = in[120]; 
    assign layer_0[333] = ~(in[246] & in[215]); 
    assign layer_0[334] = ~in[202] | (in[202] & in[85]); 
    assign layer_0[335] = ~in[54]; 
    assign layer_0[336] = ~in[184]; 
    assign layer_0[337] = ~in[123] | (in[128] & in[123]); 
    assign layer_0[338] = in[56]; 
    assign layer_0[339] = ~(in[247] | in[227]); 
    assign layer_0[340] = ~in[84]; 
    assign layer_0[341] = in[106] & ~in[195]; 
    assign layer_0[342] = ~(in[167] | in[66]); 
    assign layer_0[343] = ~(in[86] ^ in[58]); 
    assign layer_0[344] = ~in[100]; 
    assign layer_0[345] = ~(in[78] ^ in[123]); 
    assign layer_0[346] = ~in[101]; 
    assign layer_0[347] = in[214] & ~in[146]; 
    assign layer_0[348] = ~(in[38] | in[163]); 
    assign layer_0[349] = in[172] & ~in[210]; 
    assign layer_0[350] = in[227] & in[174]; 
    assign layer_0[351] = in[148]; 
    assign layer_0[352] = ~in[225] | (in[184] & in[225]); 
    assign layer_0[353] = ~in[143]; 
    assign layer_0[354] = in[27] ^ in[133]; 
    assign layer_0[355] = ~in[104] | (in[165] & in[104]); 
    assign layer_0[356] = ~in[21]; 
    assign layer_0[357] = in[178] & ~in[82]; 
    assign layer_0[358] = ~(in[24] ^ in[5]); 
    assign layer_0[359] = ~(in[64] | in[154]); 
    assign layer_0[360] = in[79]; 
    assign layer_0[361] = in[75] & ~in[3]; 
    assign layer_0[362] = in[64] ^ in[134]; 
    assign layer_0[363] = in[144] ^ in[109]; 
    assign layer_0[364] = in[103] & ~in[132]; 
    assign layer_0[365] = in[71] | in[17]; 
    assign layer_0[366] = in[247] & ~in[158]; 
    assign layer_0[367] = ~in[171]; 
    assign layer_0[368] = ~in[98]; 
    assign layer_0[369] = in[198]; 
    assign layer_0[370] = in[15] | in[44]; 
    assign layer_0[371] = in[45] | in[14]; 
    assign layer_0[372] = ~in[82]; 
    assign layer_0[373] = ~(in[220] ^ in[98]); 
    assign layer_0[374] = in[36] | in[121]; 
    assign layer_0[375] = in[79] ^ in[141]; 
    assign layer_0[376] = ~(in[151] ^ in[69]); 
    assign layer_0[377] = in[59]; 
    assign layer_0[378] = ~in[55]; 
    assign layer_0[379] = ~in[113] | (in[113] & in[56]); 
    assign layer_0[380] = ~in[120] | (in[80] & in[120]); 
    assign layer_0[381] = in[242] & ~in[173]; 
    assign layer_0[382] = in[103]; 
    assign layer_0[383] = in[118] & in[75]; 
    assign layer_0[384] = ~(in[107] & in[169]); 
    assign layer_0[385] = in[215]; 
    assign layer_0[386] = ~in[135]; 
    assign layer_0[387] = ~in[190] | (in[253] & in[190]); 
    assign layer_0[388] = ~in[238]; 
    assign layer_0[389] = ~(in[55] ^ in[150]); 
    assign layer_0[390] = in[236] | in[175]; 
    assign layer_0[391] = ~(in[217] | in[224]); 
    assign layer_0[392] = in[85] & ~in[126]; 
    assign layer_0[393] = ~in[209] | (in[209] & in[184]); 
    assign layer_0[394] = ~in[123]; 
    assign layer_0[395] = in[121]; 
    assign layer_0[396] = ~(in[237] | in[218]); 
    assign layer_0[397] = in[165]; 
    assign layer_0[398] = in[12] ^ in[73]; 
    assign layer_0[399] = in[42] | in[106]; 
    assign layer_0[400] = ~in[182] | (in[136] & in[182]); 
    assign layer_0[401] = ~(in[205] ^ in[110]); 
    assign layer_0[402] = ~(in[44] ^ in[106]); 
    assign layer_0[403] = ~(in[147] & in[76]); 
    assign layer_0[404] = ~(in[104] | in[174]); 
    assign layer_0[405] = ~in[125] | (in[67] & in[125]); 
    assign layer_0[406] = in[32]; 
    assign layer_0[407] = in[154] ^ in[199]; 
    assign layer_0[408] = ~(in[6] | in[91]); 
    assign layer_0[409] = ~(in[19] ^ in[28]); 
    assign layer_0[410] = in[204]; 
    assign layer_0[411] = in[179] & ~in[222]; 
    assign layer_0[412] = ~(in[93] | in[104]); 
    assign layer_0[413] = ~(in[175] | in[67]); 
    assign layer_0[414] = in[222] ^ in[184]; 
    assign layer_0[415] = ~(in[21] ^ in[108]); 
    assign layer_0[416] = ~(in[36] & in[95]); 
    assign layer_0[417] = ~(in[138] | in[45]); 
    assign layer_0[418] = ~in[215] | (in[215] & in[255]); 
    assign layer_0[419] = ~(in[0] | in[41]); 
    assign layer_0[420] = in[145] & ~in[30]; 
    assign layer_0[421] = ~(in[55] | in[76]); 
    assign layer_0[422] = ~(in[213] ^ in[169]); 
    assign layer_0[423] = ~(in[164] ^ in[183]); 
    assign layer_0[424] = ~(in[249] ^ in[201]); 
    assign layer_0[425] = ~(in[252] | in[128]); 
    assign layer_0[426] = ~in[195]; 
    assign layer_0[427] = ~(in[253] | in[203]); 
    assign layer_0[428] = ~(in[188] | in[165]); 
    assign layer_0[429] = ~in[74]; 
    assign layer_0[430] = in[98] & ~in[59]; 
    assign layer_0[431] = in[67] | in[121]; 
    assign layer_0[432] = in[186] | in[124]; 
    assign layer_0[433] = ~(in[43] | in[25]); 
    assign layer_0[434] = ~in[101] | (in[111] & in[101]); 
    assign layer_0[435] = ~(in[149] ^ in[163]); 
    assign layer_0[436] = ~(in[134] | in[138]); 
    assign layer_0[437] = ~(in[135] | in[153]); 
    assign layer_0[438] = ~in[146] | (in[146] & in[192]); 
    assign layer_0[439] = in[35] & in[54]; 
    assign layer_0[440] = in[148] & in[74]; 
    assign layer_0[441] = ~in[232] | (in[203] & in[232]); 
    assign layer_0[442] = in[119]; 
    assign layer_0[443] = in[87]; 
    assign layer_0[444] = ~in[186]; 
    assign layer_0[445] = ~in[73] | (in[166] & in[73]); 
    assign layer_0[446] = ~in[102]; 
    assign layer_0[447] = ~in[125] | (in[248] & in[125]); 
    assign layer_0[448] = in[198] & in[99]; 
    assign layer_0[449] = ~(in[247] & in[176]); 
    assign layer_0[450] = ~(in[37] | in[104]); 
    assign layer_0[451] = ~in[187]; 
    assign layer_0[452] = ~(in[69] ^ in[83]); 
    assign layer_0[453] = in[231] | in[248]; 
    assign layer_0[454] = in[67] ^ in[5]; 
    assign layer_0[455] = ~in[155] | (in[155] & in[94]); 
    assign layer_0[456] = ~(in[219] | in[210]); 
    assign layer_0[457] = in[232]; 
    assign layer_0[458] = in[102]; 
    assign layer_0[459] = in[90] | in[36]; 
    assign layer_0[460] = ~(in[141] ^ in[77]); 
    assign layer_0[461] = ~in[255] | (in[246] & in[255]); 
    assign layer_0[462] = ~in[144]; 
    assign layer_0[463] = ~(in[46] ^ in[40]); 
    assign layer_0[464] = ~(in[247] ^ in[241]); 
    assign layer_0[465] = in[57] & ~in[88]; 
    assign layer_0[466] = ~in[201] | (in[233] & in[201]); 
    assign layer_0[467] = ~in[152] | (in[33] & in[152]); 
    assign layer_0[468] = ~in[131]; 
    assign layer_0[469] = in[163] ^ in[67]; 
    assign layer_0[470] = in[139] ^ in[157]; 
    assign layer_0[471] = in[49]; 
    assign layer_0[472] = ~(in[149] | in[146]); 
    assign layer_0[473] = ~in[133] | (in[243] & in[133]); 
    assign layer_0[474] = in[24] ^ in[65]; 
    assign layer_0[475] = in[27] | in[140]; 
    assign layer_0[476] = in[201] & ~in[167]; 
    assign layer_0[477] = ~(in[218] & in[207]); 
    assign layer_0[478] = in[174]; 
    assign layer_0[479] = ~in[225] | (in[199] & in[225]); 
    assign layer_0[480] = ~(in[69] | in[61]); 
    assign layer_0[481] = in[209]; 
    assign layer_0[482] = in[61] ^ in[108]; 
    assign layer_0[483] = ~in[42] | (in[169] & in[42]); 
    assign layer_0[484] = in[91] & ~in[1]; 
    assign layer_0[485] = ~in[180]; 
    assign layer_0[486] = in[56]; 
    assign layer_0[487] = in[79]; 
    assign layer_0[488] = ~in[195] | (in[195] & in[198]); 
    assign layer_0[489] = in[196]; 
    assign layer_0[490] = ~in[132]; 
    assign layer_0[491] = ~(in[213] ^ in[164]); 
    assign layer_0[492] = ~in[90]; 
    assign layer_0[493] = in[223]; 
    assign layer_0[494] = ~(in[176] ^ in[67]); 
    assign layer_0[495] = in[164] & ~in[52]; 
    assign layer_0[496] = in[194]; 
    assign layer_0[497] = ~in[107]; 
    assign layer_0[498] = ~(in[235] | in[208]); 
    assign layer_0[499] = in[73] | in[133]; 
    assign layer_0[500] = ~(in[98] | in[71]); 
    assign layer_0[501] = in[29] ^ in[139]; 
    assign layer_0[502] = in[57] & ~in[2]; 
    assign layer_0[503] = ~in[92] | (in[7] & in[92]); 
    assign layer_0[504] = in[138] & ~in[38]; 
    assign layer_0[505] = in[127] ^ in[18]; 
    assign layer_0[506] = in[134] & ~in[38]; 
    assign layer_0[507] = ~in[227]; 
    assign layer_0[508] = ~in[198]; 
    assign layer_0[509] = in[233] ^ in[167]; 
    assign layer_0[510] = in[136]; 
    assign layer_0[511] = ~(in[125] & in[240]); 
    assign layer_0[512] = ~(in[35] & in[126]); 
    assign layer_0[513] = ~in[170]; 
    assign layer_0[514] = ~(in[67] ^ in[132]); 
    assign layer_0[515] = in[89]; 
    assign layer_0[516] = ~(in[54] | in[93]); 
    assign layer_0[517] = in[234]; 
    assign layer_0[518] = in[193] & ~in[178]; 
    assign layer_0[519] = in[119] & ~in[64]; 
    assign layer_0[520] = ~in[252]; 
    assign layer_0[521] = ~in[63] | (in[56] & in[63]); 
    assign layer_0[522] = ~(in[202] | in[105]); 
    assign layer_0[523] = in[225]; 
    assign layer_0[524] = in[173]; 
    assign layer_0[525] = ~(in[79] ^ in[202]); 
    assign layer_0[526] = ~in[108]; 
    assign layer_0[527] = ~(in[36] | in[143]); 
    assign layer_0[528] = in[219] | in[145]; 
    assign layer_0[529] = ~(in[13] | in[21]); 
    assign layer_0[530] = ~(in[219] ^ in[230]); 
    assign layer_0[531] = ~(in[193] & in[243]); 
    assign layer_0[532] = in[122] & ~in[189]; 
    assign layer_0[533] = in[88] & ~in[1]; 
    assign layer_0[534] = in[68] ^ in[36]; 
    assign layer_0[535] = in[203]; 
    assign layer_0[536] = in[182]; 
    assign layer_0[537] = in[123]; 
    assign layer_0[538] = in[182]; 
    assign layer_0[539] = ~in[72] | (in[72] & in[83]); 
    assign layer_0[540] = in[230] | in[251]; 
    assign layer_0[541] = in[161] & ~in[95]; 
    assign layer_0[542] = ~in[216] | (in[216] & in[160]); 
    assign layer_0[543] = ~in[56] | (in[130] & in[56]); 
    assign layer_0[544] = ~(in[108] | in[174]); 
    assign layer_0[545] = in[73] & ~in[197]; 
    assign layer_0[546] = ~in[104]; 
    assign layer_0[547] = in[167]; 
    assign layer_0[548] = ~(in[165] ^ in[239]); 
    assign layer_0[549] = ~in[14] | (in[14] & in[47]); 
    assign layer_0[550] = in[152] & ~in[28]; 
    assign layer_0[551] = ~in[108]; 
    assign layer_0[552] = ~in[219] | (in[255] & in[219]); 
    assign layer_0[553] = ~in[64] | (in[35] & in[64]); 
    assign layer_0[554] = ~in[173]; 
    assign layer_0[555] = in[119] ^ in[0]; 
    assign layer_0[556] = in[182]; 
    assign layer_0[557] = in[61] | in[164]; 
    assign layer_0[558] = ~in[69]; 
    assign layer_0[559] = ~in[46] | (in[152] & in[46]); 
    assign layer_0[560] = in[144] | in[148]; 
    assign layer_0[561] = in[246] & ~in[180]; 
    assign layer_0[562] = ~(in[220] ^ in[225]); 
    assign layer_0[563] = in[154] & in[232]; 
    assign layer_0[564] = in[170] & ~in[174]; 
    assign layer_0[565] = in[121] & ~in[38]; 
    assign layer_0[566] = in[214] & ~in[90]; 
    assign layer_0[567] = in[248] & in[128]; 
    assign layer_0[568] = ~in[138]; 
    assign layer_0[569] = in[133] | in[94]; 
    assign layer_0[570] = in[88] & ~in[114]; 
    assign layer_0[571] = ~(in[6] & in[23]); 
    assign layer_0[572] = in[74] & ~in[134]; 
    assign layer_0[573] = ~(in[94] | in[5]); 
    assign layer_0[574] = ~(in[190] | in[179]); 
    assign layer_0[575] = in[189]; 
    assign layer_0[576] = in[149] & ~in[62]; 
    assign layer_0[577] = ~(in[106] ^ in[134]); 
    assign layer_0[578] = ~(in[141] | in[65]); 
    assign layer_0[579] = ~in[110] | (in[33] & in[110]); 
    assign layer_0[580] = in[102]; 
    assign layer_0[581] = in[106] & ~in[88]; 
    assign layer_0[582] = ~(in[28] | in[52]); 
    assign layer_0[583] = in[184] | in[150]; 
    assign layer_0[584] = in[185]; 
    assign layer_0[585] = ~in[52] | (in[52] & in[13]); 
    assign layer_0[586] = ~(in[99] ^ in[183]); 
    assign layer_0[587] = ~in[197] | (in[197] & in[118]); 
    assign layer_0[588] = ~in[118]; 
    assign layer_0[589] = ~in[96] | (in[96] & in[71]); 
    assign layer_0[590] = ~(in[200] & in[143]); 
    assign layer_0[591] = in[181] ^ in[91]; 
    assign layer_0[592] = ~in[170]; 
    assign layer_0[593] = in[120] & ~in[17]; 
    assign layer_0[594] = in[175] ^ in[250]; 
    assign layer_0[595] = ~(in[155] | in[156]); 
    assign layer_0[596] = ~in[55] | (in[124] & in[55]); 
    assign layer_0[597] = ~in[116] | (in[231] & in[116]); 
    assign layer_0[598] = in[190]; 
    assign layer_0[599] = ~in[90]; 
    assign layer_0[600] = ~(in[38] ^ in[95]); 
    assign layer_0[601] = ~in[116]; 
    assign layer_0[602] = ~in[170] | (in[220] & in[170]); 
    assign layer_0[603] = in[141] & ~in[181]; 
    assign layer_0[604] = in[234] & in[248]; 
    assign layer_0[605] = in[135]; 
    assign layer_0[606] = in[151] & ~in[159]; 
    assign layer_0[607] = ~in[138]; 
    assign layer_0[608] = ~(in[248] ^ in[138]); 
    assign layer_0[609] = in[215] & ~in[97]; 
    assign layer_0[610] = ~in[116] | (in[116] & in[42]); 
    assign layer_0[611] = ~in[197] | (in[78] & in[197]); 
    assign layer_0[612] = in[119]; 
    assign layer_0[613] = ~in[32] | (in[32] & in[57]); 
    assign layer_0[614] = ~in[70]; 
    assign layer_0[615] = in[205] | in[191]; 
    assign layer_0[616] = ~in[138] | (in[80] & in[138]); 
    assign layer_0[617] = in[117] & ~in[81]; 
    assign layer_0[618] = ~in[122]; 
    assign layer_0[619] = in[224] | in[195]; 
    assign layer_0[620] = in[10] & in[92]; 
    assign layer_0[621] = ~in[56] | (in[56] & in[168]); 
    assign layer_0[622] = ~(in[115] | in[20]); 
    assign layer_0[623] = ~in[184] | (in[154] & in[184]); 
    assign layer_0[624] = in[106]; 
    assign layer_0[625] = ~in[36] | (in[17] & in[36]); 
    assign layer_0[626] = ~(in[96] | in[192]); 
    assign layer_0[627] = ~(in[209] | in[178]); 
    assign layer_0[628] = in[174]; 
    assign layer_0[629] = in[37] & ~in[27]; 
    assign layer_0[630] = in[121] ^ in[204]; 
    assign layer_0[631] = ~in[141] | (in[141] & in[38]); 
    assign layer_0[632] = in[213] | in[92]; 
    assign layer_0[633] = in[60]; 
    assign layer_0[634] = in[60] & ~in[1]; 
    assign layer_0[635] = in[6] ^ in[63]; 
    assign layer_0[636] = in[172] & ~in[62]; 
    assign layer_0[637] = ~(in[80] ^ in[145]); 
    assign layer_0[638] = ~(in[214] ^ in[93]); 
    assign layer_0[639] = ~in[37] | (in[37] & in[51]); 
    assign layer_0[640] = in[91] ^ in[47]; 
    assign layer_0[641] = in[112] ^ in[127]; 
    assign layer_0[642] = ~in[107] | (in[28] & in[107]); 
    assign layer_0[643] = ~(in[163] ^ in[183]); 
    assign layer_0[644] = ~in[91]; 
    assign layer_0[645] = in[54] & ~in[167]; 
    assign layer_0[646] = ~in[197]; 
    assign layer_0[647] = ~(in[180] | in[125]); 
    assign layer_0[648] = in[28] & in[10]; 
    assign layer_0[649] = in[204]; 
    assign layer_0[650] = in[195] | in[111]; 
    assign layer_0[651] = ~in[52] | (in[7] & in[52]); 
    assign layer_0[652] = ~in[152] | (in[63] & in[152]); 
    assign layer_0[653] = ~(in[249] | in[195]); 
    assign layer_0[654] = ~in[52] | (in[52] & in[106]); 
    assign layer_0[655] = in[70] ^ in[136]; 
    assign layer_0[656] = in[140]; 
    assign layer_0[657] = ~in[57]; 
    assign layer_0[658] = in[194] & in[189]; 
    assign layer_0[659] = in[40] & ~in[139]; 
    assign layer_0[660] = ~in[254] | (in[254] & in[209]); 
    assign layer_0[661] = ~in[157]; 
    assign layer_0[662] = in[16] | in[15]; 
    assign layer_0[663] = ~(in[138] & in[105]); 
    assign layer_0[664] = ~in[136] | (in[78] & in[136]); 
    assign layer_0[665] = in[109] & ~in[149]; 
    assign layer_0[666] = ~in[38]; 
    assign layer_0[667] = ~(in[213] ^ in[227]); 
    assign layer_0[668] = ~in[176] | (in[118] & in[176]); 
    assign layer_0[669] = in[134] ^ in[93]; 
    assign layer_0[670] = in[93] & in[42]; 
    assign layer_0[671] = in[108]; 
    assign layer_0[672] = ~in[122]; 
    assign layer_0[673] = ~in[104] | (in[133] & in[104]); 
    assign layer_0[674] = in[48] | in[73]; 
    assign layer_0[675] = ~in[99] | (in[21] & in[99]); 
    assign layer_0[676] = in[11] | in[128]; 
    assign layer_0[677] = ~(in[146] & in[129]); 
    assign layer_0[678] = in[48]; 
    assign layer_0[679] = ~(in[197] & in[142]); 
    assign layer_0[680] = ~in[147] | (in[147] & in[206]); 
    assign layer_0[681] = in[93] | in[213]; 
    assign layer_0[682] = ~in[167] | (in[196] & in[167]); 
    assign layer_0[683] = ~(in[7] | in[125]); 
    assign layer_0[684] = in[72] | in[85]; 
    assign layer_0[685] = in[70] & in[106]; 
    assign layer_0[686] = ~(in[41] | in[149]); 
    assign layer_0[687] = in[147]; 
    assign layer_0[688] = in[135]; 
    assign layer_0[689] = in[61] & ~in[161]; 
    assign layer_0[690] = ~(in[28] | in[87]); 
    assign layer_0[691] = in[83]; 
    assign layer_0[692] = ~in[155] | (in[155] & in[234]); 
    assign layer_0[693] = in[46]; 
    assign layer_0[694] = in[70] & ~in[79]; 
    assign layer_0[695] = in[149] & ~in[192]; 
    assign layer_0[696] = in[1] ^ in[42]; 
    assign layer_0[697] = in[141]; 
    assign layer_0[698] = ~in[101] | (in[101] & in[177]); 
    assign layer_0[699] = in[47] ^ in[22]; 
    assign layer_0[700] = ~(in[138] | in[244]); 
    assign layer_0[701] = ~in[118]; 
    assign layer_0[702] = ~(in[255] ^ in[128]); 
    assign layer_0[703] = ~(in[224] | in[117]); 
    assign layer_0[704] = ~in[90] | (in[22] & in[90]); 
    assign layer_0[705] = ~(in[61] ^ in[188]); 
    assign layer_0[706] = in[137] & in[74]; 
    assign layer_0[707] = in[39] | in[23]; 
    assign layer_0[708] = in[151] ^ in[172]; 
    assign layer_0[709] = in[93] | in[80]; 
    assign layer_0[710] = in[25] ^ in[98]; 
    assign layer_0[711] = ~(in[215] ^ in[223]); 
    assign layer_0[712] = ~(in[244] | in[226]); 
    assign layer_0[713] = ~in[147]; 
    assign layer_0[714] = ~in[203] | (in[110] & in[203]); 
    assign layer_0[715] = in[79]; 
    assign layer_0[716] = in[127] ^ in[82]; 
    assign layer_0[717] = ~(in[50] ^ in[34]); 
    assign layer_0[718] = in[152] & ~in[77]; 
    assign layer_0[719] = ~in[104]; 
    assign layer_0[720] = in[139] & ~in[46]; 
    assign layer_0[721] = in[157] & ~in[250]; 
    assign layer_0[722] = ~in[127] | (in[219] & in[127]); 
    assign layer_0[723] = ~(in[75] | in[94]); 
    assign layer_0[724] = ~(in[210] & in[137]); 
    assign layer_0[725] = in[111]; 
    assign layer_0[726] = in[229]; 
    assign layer_0[727] = in[226] & ~in[222]; 
    assign layer_0[728] = in[27] | in[55]; 
    assign layer_0[729] = in[195] | in[165]; 
    assign layer_0[730] = ~in[179] | (in[179] & in[100]); 
    assign layer_0[731] = ~in[74]; 
    assign layer_0[732] = ~in[101]; 
    assign layer_0[733] = ~(in[227] | in[120]); 
    assign layer_0[734] = ~in[199] | (in[249] & in[199]); 
    assign layer_0[735] = in[128] ^ in[73]; 
    assign layer_0[736] = in[245]; 
    assign layer_0[737] = in[67] | in[80]; 
    assign layer_0[738] = in[137] | in[62]; 
    assign layer_0[739] = ~in[135]; 
    assign layer_0[740] = ~(in[194] ^ in[222]); 
    assign layer_0[741] = ~(in[48] | in[155]); 
    assign layer_0[742] = in[134]; 
    assign layer_0[743] = in[255] | in[244]; 
    assign layer_0[744] = in[42] ^ in[5]; 
    assign layer_0[745] = in[201] ^ in[234]; 
    assign layer_0[746] = in[198]; 
    assign layer_0[747] = ~(in[121] & in[215]); 
    assign layer_0[748] = ~(in[217] | in[212]); 
    assign layer_0[749] = ~in[254] | (in[197] & in[254]); 
    assign layer_0[750] = in[7] & in[15]; 
    assign layer_0[751] = ~(in[198] ^ in[165]); 
    assign layer_0[752] = ~in[118]; 
    assign layer_0[753] = ~in[108] | (in[108] & in[22]); 
    assign layer_0[754] = in[88]; 
    assign layer_0[755] = in[95] ^ in[183]; 
    assign layer_0[756] = in[245] | in[218]; 
    assign layer_0[757] = in[126] | in[113]; 
    assign layer_0[758] = in[163] ^ in[219]; 
    assign layer_0[759] = ~(in[136] | in[109]); 
    assign layer_0[760] = in[87]; 
    assign layer_0[761] = in[92] & ~in[162]; 
    assign layer_0[762] = ~in[131]; 
    assign layer_0[763] = in[89]; 
    assign layer_0[764] = ~(in[203] | in[219]); 
    assign layer_0[765] = in[64] & in[86]; 
    assign layer_0[766] = ~in[132]; 
    assign layer_0[767] = ~in[53]; 
    assign layer_0[768] = ~in[149] | (in[149] & in[50]); 
    assign layer_0[769] = in[139] ^ in[206]; 
    assign layer_0[770] = ~in[18] | (in[18] & in[64]); 
    assign layer_0[771] = in[3] | in[43]; 
    assign layer_0[772] = ~(in[149] ^ in[190]); 
    assign layer_0[773] = ~in[84] | (in[121] & in[84]); 
    assign layer_0[774] = ~(in[255] | in[209]); 
    assign layer_0[775] = in[86] | in[112]; 
    assign layer_0[776] = in[39] & ~in[128]; 
    assign layer_0[777] = ~in[9] | (in[28] & in[9]); 
    assign layer_0[778] = in[31] ^ in[53]; 
    assign layer_0[779] = ~(in[25] | in[23]); 
    assign layer_0[780] = in[183] ^ in[132]; 
    assign layer_0[781] = ~in[131] | (in[131] & in[44]); 
    assign layer_0[782] = in[210]; 
    assign layer_0[783] = ~in[199]; 
    assign layer_0[784] = ~(in[79] & in[54]); 
    assign layer_0[785] = in[212] | in[178]; 
    assign layer_0[786] = ~in[205]; 
    assign layer_0[787] = in[82] | in[203]; 
    assign layer_0[788] = ~in[5]; 
    assign layer_0[789] = ~(in[235] ^ in[165]); 
    assign layer_0[790] = ~in[102] | (in[147] & in[102]); 
    assign layer_0[791] = in[171] | in[67]; 
    assign layer_0[792] = ~(in[215] ^ in[199]); 
    assign layer_0[793] = ~(in[55] & in[84]); 
    assign layer_0[794] = ~in[148] | (in[92] & in[148]); 
    assign layer_0[795] = ~in[187]; 
    assign layer_0[796] = ~in[76]; 
    assign layer_0[797] = in[102] & in[65]; 
    assign layer_0[798] = in[230] & ~in[238]; 
    assign layer_0[799] = in[228]; 
    assign layer_0[800] = ~in[143] | (in[35] & in[143]); 
    assign layer_0[801] = in[44] | in[19]; 
    assign layer_0[802] = ~(in[241] | in[249]); 
    assign layer_0[803] = ~in[219] | (in[252] & in[219]); 
    assign layer_0[804] = in[26] | in[123]; 
    assign layer_0[805] = in[196] & in[164]; 
    assign layer_0[806] = in[18] ^ in[95]; 
    assign layer_0[807] = in[134] | in[219]; 
    assign layer_0[808] = in[23] | in[39]; 
    assign layer_0[809] = ~(in[31] | in[129]); 
    assign layer_0[810] = in[168] ^ in[52]; 
    assign layer_0[811] = ~in[82] | (in[21] & in[82]); 
    assign layer_0[812] = ~in[143] | (in[31] & in[143]); 
    assign layer_0[813] = in[192] ^ in[135]; 
    assign layer_0[814] = in[118] & in[58]; 
    assign layer_0[815] = in[226]; 
    assign layer_0[816] = ~in[172]; 
    assign layer_0[817] = ~(in[48] | in[101]); 
    assign layer_0[818] = ~in[121] | (in[121] & in[65]); 
    assign layer_0[819] = ~(in[142] ^ in[204]); 
    assign layer_0[820] = in[209] | in[140]; 
    assign layer_0[821] = ~in[137] | (in[193] & in[137]); 
    assign layer_0[822] = in[204] | in[236]; 
    assign layer_0[823] = ~(in[16] & in[81]); 
    assign layer_0[824] = in[178] | in[91]; 
    assign layer_0[825] = in[140]; 
    assign layer_0[826] = ~(in[200] & in[196]); 
    assign layer_0[827] = in[40] ^ in[74]; 
    assign layer_0[828] = ~in[8]; 
    assign layer_0[829] = in[35] & ~in[81]; 
    assign layer_0[830] = in[168]; 
    assign layer_0[831] = ~(in[80] ^ in[119]); 
    assign layer_0[832] = in[89]; 
    assign layer_0[833] = in[158] ^ in[105]; 
    assign layer_0[834] = in[120] & ~in[233]; 
    assign layer_0[835] = in[194] & ~in[200]; 
    assign layer_0[836] = ~(in[76] | in[170]); 
    assign layer_0[837] = in[161]; 
    assign layer_0[838] = in[175] & in[91]; 
    assign layer_0[839] = in[3] | in[0]; 
    assign layer_0[840] = ~in[163] | (in[206] & in[163]); 
    assign layer_0[841] = ~in[117]; 
    assign layer_0[842] = in[138] & ~in[161]; 
    assign layer_0[843] = in[102] & ~in[127]; 
    assign layer_0[844] = in[156]; 
    assign layer_0[845] = ~(in[75] | in[96]); 
    assign layer_0[846] = ~(in[24] & in[144]); 
    assign layer_0[847] = ~in[91] | (in[94] & in[91]); 
    assign layer_0[848] = in[156] & ~in[63]; 
    assign layer_0[849] = ~in[66]; 
    assign layer_0[850] = ~in[211] | (in[211] & in[93]); 
    assign layer_0[851] = ~(in[105] & in[95]); 
    assign layer_0[852] = in[59]; 
    assign layer_0[853] = ~(in[15] ^ in[60]); 
    assign layer_0[854] = in[247]; 
    assign layer_0[855] = ~(in[23] | in[56]); 
    assign layer_0[856] = ~in[237]; 
    assign layer_0[857] = ~in[176] | (in[202] & in[176]); 
    assign layer_0[858] = in[148]; 
    assign layer_0[859] = ~in[156] | (in[50] & in[156]); 
    assign layer_0[860] = ~in[197]; 
    assign layer_0[861] = ~(in[178] ^ in[176]); 
    assign layer_0[862] = in[72] & ~in[2]; 
    assign layer_0[863] = ~in[125]; 
    assign layer_0[864] = in[199] & in[155]; 
    assign layer_0[865] = ~in[77]; 
    assign layer_0[866] = ~in[81] | (in[39] & in[81]); 
    assign layer_0[867] = ~in[135]; 
    assign layer_0[868] = ~in[2] | (in[2] & in[83]); 
    assign layer_0[869] = in[211] & ~in[251]; 
    assign layer_0[870] = in[160] | in[85]; 
    assign layer_0[871] = ~in[114] | (in[157] & in[114]); 
    assign layer_0[872] = ~(in[221] | in[252]); 
    assign layer_0[873] = in[177] & ~in[254]; 
    assign layer_0[874] = ~(in[235] ^ in[238]); 
    assign layer_0[875] = in[202] & ~in[114]; 
    assign layer_0[876] = in[142] & in[40]; 
    assign layer_0[877] = ~in[93] | (in[9] & in[93]); 
    assign layer_0[878] = in[228]; 
    assign layer_0[879] = in[40] ^ in[143]; 
    assign layer_0[880] = in[143] & ~in[163]; 
    assign layer_0[881] = in[132]; 
    assign layer_0[882] = in[119] & in[233]; 
    assign layer_0[883] = ~in[93]; 
    assign layer_0[884] = ~(in[12] | in[78]); 
    assign layer_0[885] = ~(in[203] & in[127]); 
    assign layer_0[886] = in[178] | in[122]; 
    assign layer_0[887] = in[38]; 
    assign layer_0[888] = in[70]; 
    assign layer_0[889] = in[21] & ~in[3]; 
    assign layer_0[890] = ~in[20]; 
    assign layer_0[891] = ~(in[123] ^ in[105]); 
    assign layer_0[892] = ~in[248]; 
    assign layer_0[893] = in[241] ^ in[176]; 
    assign layer_0[894] = in[121] ^ in[125]; 
    assign layer_0[895] = ~in[64] | (in[171] & in[64]); 
    assign layer_0[896] = in[180]; 
    assign layer_0[897] = in[11] & in[63]; 
    assign layer_0[898] = ~in[66]; 
    assign layer_0[899] = ~in[16] | (in[16] & in[135]); 
    assign layer_0[900] = ~(in[201] | in[226]); 
    assign layer_0[901] = ~in[238] | (in[194] & in[238]); 
    assign layer_0[902] = in[179]; 
    assign layer_0[903] = ~in[73] | (in[73] & in[143]); 
    assign layer_0[904] = in[168]; 
    assign layer_0[905] = ~in[151]; 
    assign layer_0[906] = in[244]; 
    assign layer_0[907] = in[92] & ~in[27]; 
    assign layer_0[908] = ~(in[51] | in[75]); 
    assign layer_0[909] = in[120]; 
    assign layer_0[910] = in[204] | in[138]; 
    assign layer_0[911] = in[75] & ~in[9]; 
    assign layer_0[912] = in[216] & ~in[156]; 
    assign layer_0[913] = in[141] ^ in[25]; 
    assign layer_0[914] = ~in[63]; 
    assign layer_0[915] = ~(in[96] | in[184]); 
    assign layer_0[916] = in[20] & ~in[76]; 
    assign layer_0[917] = ~(in[170] ^ in[173]); 
    assign layer_0[918] = in[58] & ~in[183]; 
    assign layer_0[919] = in[171] & ~in[89]; 
    assign layer_0[920] = in[25]; 
    assign layer_0[921] = in[109] | in[114]; 
    assign layer_0[922] = ~in[235]; 
    assign layer_0[923] = ~(in[93] | in[9]); 
    assign layer_0[924] = ~in[117]; 
    assign layer_0[925] = ~in[183]; 
    assign layer_0[926] = in[233]; 
    assign layer_0[927] = in[199]; 
    assign layer_0[928] = ~in[48]; 
    assign layer_0[929] = in[110] & ~in[226]; 
    assign layer_0[930] = in[118]; 
    assign layer_0[931] = ~in[77]; 
    assign layer_0[932] = in[92]; 
    assign layer_0[933] = ~(in[194] | in[67]); 
    assign layer_0[934] = in[116]; 
    assign layer_0[935] = ~in[48] | (in[48] & in[169]); 
    assign layer_0[936] = ~in[155] | (in[81] & in[155]); 
    assign layer_0[937] = ~(in[216] & in[142]); 
    assign layer_0[938] = in[215] ^ in[90]; 
    assign layer_0[939] = in[143]; 
    assign layer_0[940] = in[154] & in[73]; 
    assign layer_0[941] = in[241] & in[153]; 
    assign layer_0[942] = ~(in[244] & in[129]); 
    assign layer_0[943] = ~(in[157] ^ in[222]); 
    assign layer_0[944] = ~in[58] | (in[58] & in[1]); 
    assign layer_0[945] = in[120] & ~in[167]; 
    assign layer_0[946] = ~(in[249] ^ in[178]); 
    assign layer_0[947] = in[181]; 
    assign layer_0[948] = ~(in[11] ^ in[107]); 
    assign layer_0[949] = in[150] & ~in[171]; 
    assign layer_0[950] = ~(in[84] | in[149]); 
    assign layer_0[951] = ~in[182] | (in[246] & in[182]); 
    assign layer_0[952] = ~in[21] | (in[21] & in[58]); 
    assign layer_0[953] = in[53] & in[138]; 
    assign layer_0[954] = in[124]; 
    assign layer_0[955] = in[135] | in[94]; 
    assign layer_0[956] = ~in[104] | (in[104] & in[142]); 
    assign layer_0[957] = ~(in[235] | in[141]); 
    assign layer_0[958] = ~in[176]; 
    assign layer_0[959] = in[5]; 
    assign layer_0[960] = ~in[6] | (in[6] & in[48]); 
    assign layer_0[961] = ~in[118]; 
    assign layer_0[962] = ~(in[126] | in[115]); 
    assign layer_0[963] = in[224] & in[245]; 
    assign layer_0[964] = ~(in[153] ^ in[142]); 
    assign layer_0[965] = in[102] ^ in[5]; 
    assign layer_0[966] = in[232]; 
    assign layer_0[967] = ~(in[110] | in[87]); 
    assign layer_0[968] = ~in[251] | (in[255] & in[251]); 
    assign layer_0[969] = in[143]; 
    assign layer_0[970] = in[17] | in[60]; 
    assign layer_0[971] = ~(in[226] & in[182]); 
    assign layer_0[972] = ~in[56] | (in[153] & in[56]); 
    assign layer_0[973] = ~(in[169] & in[65]); 
    assign layer_0[974] = ~in[85]; 
    assign layer_0[975] = ~in[62]; 
    assign layer_0[976] = ~in[116]; 
    assign layer_0[977] = ~(in[248] ^ in[146]); 
    assign layer_0[978] = ~in[224] | (in[246] & in[224]); 
    assign layer_0[979] = ~(in[67] & in[2]); 
    assign layer_0[980] = in[203] | in[213]; 
    assign layer_0[981] = in[72] ^ in[37]; 
    assign layer_0[982] = in[111] ^ in[97]; 
    assign layer_0[983] = ~(in[112] | in[220]); 
    assign layer_0[984] = ~(in[63] | in[131]); 
    assign layer_0[985] = in[158] | in[204]; 
    assign layer_0[986] = ~(in[186] ^ in[250]); 
    assign layer_0[987] = in[151] & in[163]; 
    assign layer_0[988] = ~(in[13] | in[124]); 
    assign layer_0[989] = ~in[105]; 
    assign layer_0[990] = in[159] & in[74]; 
    assign layer_0[991] = in[32]; 
    assign layer_0[992] = in[168] | in[166]; 
    assign layer_0[993] = in[57] & ~in[7]; 
    assign layer_0[994] = ~in[65]; 
    assign layer_0[995] = in[218] & ~in[234]; 
    assign layer_0[996] = ~(in[38] | in[85]); 
    assign layer_0[997] = in[152] ^ in[168]; 
    assign layer_0[998] = ~in[145] | (in[145] & in[83]); 
    assign layer_0[999] = ~in[122]; 
    assign layer_0[1000] = in[160]; 
    assign layer_0[1001] = ~in[137] | (in[243] & in[137]); 
    assign layer_0[1002] = ~in[184] | (in[184] & in[91]); 
    assign layer_0[1003] = in[99] ^ in[102]; 
    assign layer_0[1004] = in[165]; 
    assign layer_0[1005] = ~(in[218] | in[227]); 
    assign layer_0[1006] = ~in[166] | (in[82] & in[166]); 
    assign layer_0[1007] = ~(in[104] ^ in[116]); 
    assign layer_0[1008] = ~(in[47] & in[143]); 
    assign layer_0[1009] = ~in[45] | (in[45] & in[48]); 
    assign layer_0[1010] = in[90]; 
    assign layer_0[1011] = ~(in[144] | in[168]); 
    assign layer_0[1012] = in[174]; 
    assign layer_0[1013] = in[76] | in[201]; 
    assign layer_0[1014] = in[254]; 
    assign layer_0[1015] = in[14] | in[77]; 
    assign layer_0[1016] = in[73] | in[65]; 
    assign layer_0[1017] = in[90] | in[173]; 
    assign layer_0[1018] = ~(in[121] | in[129]); 
    assign layer_0[1019] = in[244] & in[222]; 
    assign layer_0[1020] = ~in[233]; 
    assign layer_0[1021] = ~in[130]; 
    assign layer_0[1022] = in[200] ^ in[175]; 
    assign layer_0[1023] = ~(in[193] | in[179]); 
    assign layer_0[1024] = ~(in[161] ^ in[121]); 
    assign layer_0[1025] = in[117]; 
    assign layer_0[1026] = ~in[98]; 
    assign layer_0[1027] = in[51] & in[0]; 
    assign layer_0[1028] = ~(in[165] | in[229]); 
    assign layer_0[1029] = in[88] & ~in[212]; 
    assign layer_0[1030] = in[27]; 
    assign layer_0[1031] = in[35]; 
    assign layer_0[1032] = ~in[134] | (in[210] & in[134]); 
    assign layer_0[1033] = ~(in[167] ^ in[113]); 
    assign layer_0[1034] = in[41] ^ in[143]; 
    assign layer_0[1035] = ~in[127] | (in[64] & in[127]); 
    assign layer_0[1036] = in[169] & ~in[162]; 
    assign layer_0[1037] = in[88]; 
    assign layer_0[1038] = in[76] ^ in[127]; 
    assign layer_0[1039] = ~in[149]; 
    assign layer_0[1040] = in[51] ^ in[92]; 
    assign layer_0[1041] = ~(in[179] & in[235]); 
    assign layer_0[1042] = ~in[59] | (in[59] & in[45]); 
    assign layer_0[1043] = ~(in[155] | in[29]); 
    assign layer_0[1044] = in[42] ^ in[126]; 
    assign layer_0[1045] = in[119] & in[210]; 
    assign layer_0[1046] = in[170] & ~in[94]; 
    assign layer_0[1047] = ~in[85]; 
    assign layer_0[1048] = ~(in[68] | in[148]); 
    assign layer_0[1049] = in[161] & ~in[221]; 
    assign layer_0[1050] = ~in[185] | (in[207] & in[185]); 
    assign layer_0[1051] = in[82]; 
    assign layer_0[1052] = in[108]; 
    assign layer_0[1053] = in[136] ^ in[242]; 
    assign layer_0[1054] = in[42]; 
    assign layer_0[1055] = in[41] & in[113]; 
    assign layer_0[1056] = ~(in[112] | in[9]); 
    assign layer_0[1057] = ~in[224]; 
    assign layer_0[1058] = in[234] | in[248]; 
    assign layer_0[1059] = in[153] | in[52]; 
    assign layer_0[1060] = ~in[99]; 
    assign layer_0[1061] = ~(in[87] & in[147]); 
    assign layer_0[1062] = ~in[123] | (in[123] & in[164]); 
    assign layer_0[1063] = in[190] | in[249]; 
    assign layer_0[1064] = in[121] | in[226]; 
    assign layer_0[1065] = ~in[163] | (in[163] & in[204]); 
    assign layer_0[1066] = ~in[84]; 
    assign layer_0[1067] = ~(in[23] ^ in[14]); 
    assign layer_0[1068] = in[230]; 
    assign layer_0[1069] = in[65] & ~in[0]; 
    assign layer_0[1070] = in[107] & ~in[63]; 
    assign layer_0[1071] = ~in[189] | (in[189] & in[73]); 
    assign layer_0[1072] = ~in[151]; 
    assign layer_0[1073] = in[200] & ~in[100]; 
    assign layer_0[1074] = ~in[60] | (in[93] & in[60]); 
    assign layer_0[1075] = ~in[102] | (in[102] & in[165]); 
    assign layer_0[1076] = in[217] & ~in[254]; 
    assign layer_0[1077] = ~in[176]; 
    assign layer_0[1078] = ~in[86]; 
    assign layer_0[1079] = ~(in[180] ^ in[228]); 
    assign layer_0[1080] = in[154]; 
    assign layer_0[1081] = in[160] & in[137]; 
    assign layer_0[1082] = ~in[88] | (in[126] & in[88]); 
    assign layer_0[1083] = ~in[60] | (in[60] & in[84]); 
    assign layer_0[1084] = ~(in[84] ^ in[58]); 
    assign layer_0[1085] = in[51] | in[27]; 
    assign layer_0[1086] = in[96] ^ in[176]; 
    assign layer_0[1087] = ~in[71] | (in[147] & in[71]); 
    assign layer_0[1088] = ~(in[107] ^ in[139]); 
    assign layer_0[1089] = in[135]; 
    assign layer_0[1090] = in[128] | in[138]; 
    assign layer_0[1091] = ~(in[203] | in[172]); 
    assign layer_0[1092] = in[201]; 
    assign layer_0[1093] = in[171]; 
    assign layer_0[1094] = ~(in[126] | in[182]); 
    assign layer_0[1095] = ~(in[111] ^ in[84]); 
    assign layer_0[1096] = in[223] & ~in[228]; 
    assign layer_0[1097] = in[165] & ~in[111]; 
    assign layer_0[1098] = in[172] | in[250]; 
    assign layer_0[1099] = in[185] ^ in[147]; 
    assign layer_0[1100] = ~in[100] | (in[211] & in[100]); 
    assign layer_0[1101] = in[87] & ~in[209]; 
    assign layer_0[1102] = ~in[65] | (in[178] & in[65]); 
    assign layer_0[1103] = in[187] ^ in[250]; 
    assign layer_0[1104] = ~in[144] | (in[205] & in[144]); 
    assign layer_0[1105] = ~in[93]; 
    assign layer_0[1106] = ~in[223] | (in[223] & in[247]); 
    assign layer_0[1107] = in[227] | in[148]; 
    assign layer_0[1108] = in[7]; 
    assign layer_0[1109] = ~in[168] | (in[239] & in[168]); 
    assign layer_0[1110] = in[230] & ~in[181]; 
    assign layer_0[1111] = in[233] & in[134]; 
    assign layer_0[1112] = in[235] ^ in[125]; 
    assign layer_0[1113] = ~in[124]; 
    assign layer_0[1114] = in[92] & in[58]; 
    assign layer_0[1115] = in[209] | in[138]; 
    assign layer_0[1116] = in[211]; 
    assign layer_0[1117] = in[35]; 
    assign layer_0[1118] = ~in[230]; 
    assign layer_0[1119] = ~in[94] | (in[25] & in[94]); 
    assign layer_0[1120] = ~in[254] | (in[254] & in[176]); 
    assign layer_0[1121] = ~in[216] | (in[159] & in[216]); 
    assign layer_0[1122] = ~in[229]; 
    assign layer_0[1123] = in[72] & ~in[45]; 
    assign layer_0[1124] = ~in[57]; 
    assign layer_0[1125] = ~in[103]; 
    assign layer_0[1126] = ~(in[248] | in[228]); 
    assign layer_0[1127] = ~in[188]; 
    assign layer_0[1128] = in[105] & ~in[54]; 
    assign layer_0[1129] = ~(in[176] | in[235]); 
    assign layer_0[1130] = in[99]; 
    assign layer_0[1131] = ~(in[58] ^ in[49]); 
    assign layer_0[1132] = ~(in[96] | in[224]); 
    assign layer_0[1133] = in[131] & in[147]; 
    assign layer_0[1134] = ~in[87]; 
    assign layer_0[1135] = in[155] & in[129]; 
    assign layer_0[1136] = in[83]; 
    assign layer_0[1137] = in[107]; 
    assign layer_0[1138] = in[225] ^ in[163]; 
    assign layer_0[1139] = in[243] ^ in[186]; 
    assign layer_0[1140] = ~in[104] | (in[104] & in[10]); 
    assign layer_0[1141] = in[34] & ~in[40]; 
    assign layer_0[1142] = ~in[68]; 
    assign layer_0[1143] = ~in[168]; 
    assign layer_0[1144] = ~in[115] | (in[45] & in[115]); 
    assign layer_0[1145] = in[250] & in[242]; 
    assign layer_0[1146] = in[172] | in[106]; 
    assign layer_0[1147] = ~in[232]; 
    assign layer_0[1148] = ~(in[169] | in[42]); 
    assign layer_0[1149] = in[78]; 
    assign layer_0[1150] = ~in[75] | (in[20] & in[75]); 
    assign layer_0[1151] = in[136] & ~in[179]; 
    assign layer_0[1152] = in[174] ^ in[92]; 
    assign layer_0[1153] = in[178] | in[162]; 
    assign layer_0[1154] = ~in[168]; 
    assign layer_0[1155] = in[216]; 
    assign layer_0[1156] = ~in[230] | (in[149] & in[230]); 
    assign layer_0[1157] = ~in[159] | (in[159] & in[31]); 
    assign layer_0[1158] = in[117] & in[111]; 
    assign layer_0[1159] = in[160] & in[32]; 
    assign layer_0[1160] = in[115]; 
    assign layer_0[1161] = in[220] & in[161]; 
    assign layer_0[1162] = ~(in[140] | in[97]); 
    assign layer_0[1163] = ~(in[114] ^ in[200]); 
    assign layer_0[1164] = in[214] & in[233]; 
    assign layer_0[1165] = ~in[164] | (in[164] & in[227]); 
    assign layer_0[1166] = in[124] & ~in[80]; 
    assign layer_0[1167] = ~(in[140] & in[58]); 
    assign layer_0[1168] = in[250] ^ in[239]; 
    assign layer_0[1169] = ~(in[251] ^ in[241]); 
    assign layer_0[1170] = in[214] & ~in[236]; 
    assign layer_0[1171] = ~in[89]; 
    assign layer_0[1172] = ~(in[234] | in[138]); 
    assign layer_0[1173] = in[26]; 
    assign layer_0[1174] = ~(in[175] | in[235]); 
    assign layer_0[1175] = in[85] & ~in[115]; 
    assign layer_0[1176] = ~(in[17] & in[30]); 
    assign layer_0[1177] = in[123] & ~in[227]; 
    assign layer_0[1178] = ~(in[70] & in[121]); 
    assign layer_0[1179] = in[96] | in[165]; 
    assign layer_0[1180] = ~in[94]; 
    assign layer_0[1181] = in[159] ^ in[165]; 
    assign layer_0[1182] = ~in[26]; 
    assign layer_0[1183] = ~in[148] | (in[195] & in[148]); 
    assign layer_0[1184] = ~in[178] | (in[178] & in[149]); 
    assign layer_0[1185] = in[185] & ~in[235]; 
    assign layer_0[1186] = in[100]; 
    assign layer_0[1187] = ~in[90]; 
    assign layer_0[1188] = ~in[8]; 
    assign layer_0[1189] = ~(in[202] | in[232]); 
    assign layer_0[1190] = in[80]; 
    assign layer_0[1191] = ~(in[4] ^ in[0]); 
    assign layer_0[1192] = ~(in[173] | in[157]); 
    assign layer_0[1193] = ~in[157]; 
    assign layer_0[1194] = ~in[106]; 
    assign layer_0[1195] = ~(in[36] & in[37]); 
    assign layer_0[1196] = ~(in[254] ^ in[189]); 
    assign layer_0[1197] = in[142] | in[63]; 
    assign layer_0[1198] = ~(in[26] ^ in[37]); 
    assign layer_0[1199] = ~(in[201] | in[253]); 
    assign layer_0[1200] = in[215]; 
    assign layer_0[1201] = in[112]; 
    assign layer_0[1202] = ~in[100] | (in[219] & in[100]); 
    assign layer_0[1203] = ~in[150]; 
    assign layer_0[1204] = in[178]; 
    assign layer_0[1205] = in[189]; 
    assign layer_0[1206] = ~in[70] | (in[112] & in[70]); 
    assign layer_0[1207] = in[160] & ~in[153]; 
    assign layer_0[1208] = ~in[61] | (in[11] & in[61]); 
    assign layer_0[1209] = in[34] & in[94]; 
    assign layer_0[1210] = in[107] | in[82]; 
    assign layer_0[1211] = ~in[228] | (in[228] & in[241]); 
    assign layer_0[1212] = in[156] & ~in[142]; 
    assign layer_0[1213] = ~in[18] | (in[18] & in[29]); 
    assign layer_0[1214] = ~in[71]; 
    assign layer_0[1215] = in[212] | in[98]; 
    assign layer_0[1216] = ~in[182] | (in[178] & in[182]); 
    assign layer_0[1217] = ~in[219]; 
    assign layer_0[1218] = ~in[105]; 
    assign layer_0[1219] = ~in[59] | (in[101] & in[59]); 
    assign layer_0[1220] = ~in[7]; 
    assign layer_0[1221] = in[139] | in[86]; 
    assign layer_0[1222] = in[56] & ~in[15]; 
    assign layer_0[1223] = ~in[58] | (in[40] & in[58]); 
    assign layer_0[1224] = ~in[119]; 
    assign layer_0[1225] = ~(in[209] | in[255]); 
    assign layer_0[1226] = ~in[47] | (in[47] & in[136]); 
    assign layer_0[1227] = ~in[121] | (in[27] & in[121]); 
    assign layer_0[1228] = ~(in[3] ^ in[50]); 
    assign layer_0[1229] = ~in[153] | (in[204] & in[153]); 
    assign layer_0[1230] = in[151] & in[198]; 
    assign layer_0[1231] = in[214] | in[203]; 
    assign layer_0[1232] = ~in[107] | (in[107] & in[178]); 
    assign layer_0[1233] = in[43] & in[48]; 
    assign layer_0[1234] = in[85] & in[46]; 
    assign layer_0[1235] = ~in[175] | (in[223] & in[175]); 
    assign layer_0[1236] = in[88] ^ in[142]; 
    assign layer_0[1237] = in[165] & ~in[189]; 
    assign layer_0[1238] = ~in[123] | (in[166] & in[123]); 
    assign layer_0[1239] = ~in[75]; 
    assign layer_0[1240] = in[38] | in[55]; 
    assign layer_0[1241] = ~(in[173] | in[115]); 
    assign layer_0[1242] = in[11] & ~in[56]; 
    assign layer_0[1243] = ~in[99] | (in[99] & in[78]); 
    assign layer_0[1244] = in[203] ^ in[172]; 
    assign layer_0[1245] = in[92] ^ in[45]; 
    assign layer_0[1246] = in[221] & in[250]; 
    assign layer_0[1247] = in[81]; 
    assign layer_0[1248] = ~(in[225] ^ in[109]); 
    assign layer_0[1249] = in[98] & ~in[2]; 
    assign layer_0[1250] = ~in[153] | (in[209] & in[153]); 
    assign layer_0[1251] = ~(in[149] & in[64]); 
    assign layer_0[1252] = in[151]; 
    assign layer_0[1253] = in[197] ^ in[75]; 
    assign layer_0[1254] = ~in[138]; 
    assign layer_0[1255] = in[216] & in[107]; 
    assign layer_0[1256] = in[122] & ~in[143]; 
    assign layer_0[1257] = in[247] ^ in[191]; 
    assign layer_0[1258] = in[109] ^ in[145]; 
    assign layer_0[1259] = in[124]; 
    assign layer_0[1260] = ~in[253]; 
    assign layer_0[1261] = ~in[0]; 
    assign layer_0[1262] = in[3] & ~in[96]; 
    assign layer_0[1263] = in[229] ^ in[174]; 
    assign layer_0[1264] = ~(in[132] & in[33]); 
    assign layer_0[1265] = in[136] & ~in[241]; 
    assign layer_0[1266] = ~in[30] | (in[30] & in[28]); 
    assign layer_0[1267] = ~in[207]; 
    assign layer_0[1268] = in[60] & in[99]; 
    assign layer_0[1269] = ~(in[25] | in[146]); 
    assign layer_0[1270] = ~in[182] | (in[91] & in[182]); 
    assign layer_0[1271] = ~in[103] | (in[103] & in[87]); 
    assign layer_0[1272] = in[115]; 
    assign layer_0[1273] = ~in[56] | (in[56] & in[10]); 
    assign layer_0[1274] = in[116]; 
    assign layer_0[1275] = in[189] | in[210]; 
    assign layer_0[1276] = in[61]; 
    assign layer_0[1277] = ~in[199]; 
    assign layer_0[1278] = ~(in[233] ^ in[214]); 
    assign layer_0[1279] = in[184] & ~in[220]; 
    assign layer_0[1280] = ~in[211]; 
    assign layer_0[1281] = ~in[100] | (in[100] & in[95]); 
    assign layer_0[1282] = in[177] & ~in[241]; 
    assign layer_0[1283] = in[228] & ~in[254]; 
    assign layer_0[1284] = in[183] & ~in[70]; 
    assign layer_0[1285] = ~(in[95] ^ in[8]); 
    assign layer_0[1286] = in[101]; 
    assign layer_0[1287] = in[132] & ~in[22]; 
    assign layer_0[1288] = in[98] & ~in[96]; 
    assign layer_0[1289] = ~(in[143] ^ in[202]); 
    assign layer_0[1290] = in[75] | in[42]; 
    assign layer_0[1291] = in[197] | in[93]; 
    assign layer_0[1292] = in[220]; 
    assign layer_0[1293] = ~in[164]; 
    assign layer_0[1294] = ~in[71]; 
    assign layer_0[1295] = ~(in[254] | in[196]); 
    assign layer_0[1296] = ~(in[209] ^ in[180]); 
    assign layer_0[1297] = in[134] ^ in[177]; 
    assign layer_0[1298] = in[184] & in[189]; 
    assign layer_0[1299] = in[216]; 
    assign layer_0[1300] = in[162] | in[218]; 
    assign layer_0[1301] = in[174] | in[61]; 
    assign layer_0[1302] = ~(in[111] ^ in[182]); 
    assign layer_0[1303] = in[135]; 
    assign layer_0[1304] = in[201] & in[238]; 
    assign layer_0[1305] = ~in[251] | (in[201] & in[251]); 
    assign layer_0[1306] = ~(in[13] | in[77]); 
    assign layer_0[1307] = ~in[30] | (in[64] & in[30]); 
    assign layer_0[1308] = in[86] | in[85]; 
    assign layer_0[1309] = ~in[236] | (in[236] & in[196]); 
    assign layer_0[1310] = ~(in[101] | in[124]); 
    assign layer_0[1311] = ~in[170] | (in[170] & in[230]); 
    assign layer_0[1312] = ~in[147]; 
    assign layer_0[1313] = ~(in[74] & in[97]); 
    assign layer_0[1314] = ~in[107]; 
    assign layer_0[1315] = ~in[62]; 
    assign layer_0[1316] = ~in[202]; 
    assign layer_0[1317] = in[172] ^ in[62]; 
    assign layer_0[1318] = in[19] | in[22]; 
    assign layer_0[1319] = ~in[81] | (in[81] & in[113]); 
    assign layer_0[1320] = ~(in[194] | in[156]); 
    assign layer_0[1321] = ~in[95]; 
    assign layer_0[1322] = in[154] & ~in[224]; 
    assign layer_0[1323] = ~(in[117] ^ in[96]); 
    assign layer_0[1324] = in[111] | in[88]; 
    assign layer_0[1325] = ~(in[42] | in[141]); 
    assign layer_0[1326] = ~in[103]; 
    assign layer_0[1327] = ~(in[109] | in[107]); 
    assign layer_0[1328] = in[7] | in[128]; 
    assign layer_0[1329] = ~(in[24] | in[69]); 
    assign layer_0[1330] = ~in[181]; 
    assign layer_0[1331] = ~in[170] | (in[170] & in[131]); 
    assign layer_0[1332] = ~in[63]; 
    assign layer_0[1333] = ~(in[201] | in[81]); 
    assign layer_0[1334] = in[74]; 
    assign layer_0[1335] = in[122]; 
    assign layer_0[1336] = ~(in[185] ^ in[230]); 
    assign layer_0[1337] = in[83]; 
    assign layer_0[1338] = in[4] ^ in[53]; 
    assign layer_0[1339] = ~(in[53] & in[133]); 
    assign layer_0[1340] = in[19]; 
    assign layer_0[1341] = in[62] & ~in[72]; 
    assign layer_0[1342] = ~(in[73] ^ in[53]); 
    assign layer_0[1343] = in[122] & ~in[222]; 
    assign layer_0[1344] = in[164] ^ in[182]; 
    assign layer_0[1345] = in[196] ^ in[226]; 
    assign layer_0[1346] = in[0] & ~in[60]; 
    assign layer_0[1347] = in[134]; 
    assign layer_0[1348] = ~(in[174] | in[203]); 
    assign layer_0[1349] = ~in[150] | (in[150] & in[34]); 
    assign layer_0[1350] = ~in[215]; 
    assign layer_0[1351] = ~in[225] | (in[225] & in[237]); 
    assign layer_0[1352] = ~in[194]; 
    assign layer_0[1353] = ~in[125]; 
    assign layer_0[1354] = ~in[71]; 
    assign layer_0[1355] = in[164] & ~in[134]; 
    assign layer_0[1356] = in[109]; 
    assign layer_0[1357] = ~in[43] | (in[43] & in[22]); 
    assign layer_0[1358] = in[155]; 
    assign layer_0[1359] = in[52] | in[149]; 
    assign layer_0[1360] = in[141] & ~in[206]; 
    assign layer_0[1361] = ~(in[9] ^ in[73]); 
    assign layer_0[1362] = in[100] & ~in[163]; 
    assign layer_0[1363] = ~in[86] | (in[147] & in[86]); 
    assign layer_0[1364] = in[99] ^ in[171]; 
    assign layer_0[1365] = in[17] | in[45]; 
    assign layer_0[1366] = in[86] & ~in[161]; 
    assign layer_0[1367] = ~in[196]; 
    assign layer_0[1368] = ~(in[60] ^ in[157]); 
    assign layer_0[1369] = in[1] ^ in[43]; 
    assign layer_0[1370] = ~in[56]; 
    assign layer_0[1371] = ~(in[216] | in[98]); 
    assign layer_0[1372] = in[80] | in[201]; 
    assign layer_0[1373] = in[14]; 
    assign layer_0[1374] = in[85]; 
    assign layer_0[1375] = ~in[160] | (in[247] & in[160]); 
    assign layer_0[1376] = ~in[212]; 
    assign layer_0[1377] = in[208]; 
    assign layer_0[1378] = ~(in[70] & in[92]); 
    assign layer_0[1379] = ~in[21]; 
    assign layer_0[1380] = in[130] ^ in[73]; 
    assign layer_0[1381] = in[82] ^ in[160]; 
    assign layer_0[1382] = in[91]; 
    assign layer_0[1383] = ~(in[223] ^ in[252]); 
    assign layer_0[1384] = in[74] & in[11]; 
    assign layer_0[1385] = ~in[255] | (in[206] & in[255]); 
    assign layer_0[1386] = ~(in[45] | in[140]); 
    assign layer_0[1387] = ~in[141]; 
    assign layer_0[1388] = in[147] & ~in[65]; 
    assign layer_0[1389] = in[195] | in[232]; 
    assign layer_0[1390] = ~in[120]; 
    assign layer_0[1391] = ~in[72] | (in[72] & in[134]); 
    assign layer_0[1392] = ~(in[12] | in[86]); 
    assign layer_0[1393] = in[151]; 
    assign layer_0[1394] = in[87]; 
    assign layer_0[1395] = in[167] & in[77]; 
    assign layer_0[1396] = in[106] & ~in[53]; 
    assign layer_0[1397] = ~in[119] | (in[119] & in[24]); 
    assign layer_0[1398] = in[105] | in[96]; 
    assign layer_0[1399] = ~(in[72] | in[41]); 
    assign layer_0[1400] = ~in[186]; 
    assign layer_0[1401] = in[218] & ~in[220]; 
    assign layer_0[1402] = ~in[85] | (in[172] & in[85]); 
    assign layer_0[1403] = in[11] | in[21]; 
    assign layer_0[1404] = ~in[94]; 
    assign layer_0[1405] = in[56] & ~in[148]; 
    assign layer_0[1406] = in[245] ^ in[200]; 
    assign layer_0[1407] = ~in[102] | (in[39] & in[102]); 
    assign layer_0[1408] = in[93] & in[210]; 
    assign layer_0[1409] = ~in[136] | (in[136] & in[8]); 
    assign layer_0[1410] = ~in[86] | (in[86] & in[111]); 
    assign layer_0[1411] = in[54]; 
    assign layer_0[1412] = in[205] | in[124]; 
    assign layer_0[1413] = in[23]; 
    assign layer_0[1414] = ~in[170]; 
    assign layer_0[1415] = in[15] | in[133]; 
    assign layer_0[1416] = ~(in[165] | in[208]); 
    assign layer_0[1417] = ~(in[203] | in[165]); 
    assign layer_0[1418] = in[155] & ~in[177]; 
    assign layer_0[1419] = ~in[213] | (in[213] & in[129]); 
    assign layer_0[1420] = in[6]; 
    assign layer_0[1421] = in[65] & in[151]; 
    assign layer_0[1422] = in[45] & ~in[5]; 
    assign layer_0[1423] = in[142] | in[120]; 
    assign layer_0[1424] = ~in[172]; 
    assign layer_0[1425] = in[30] & ~in[2]; 
    assign layer_0[1426] = ~in[178] | (in[104] & in[178]); 
    assign layer_0[1427] = ~(in[105] ^ in[224]); 
    assign layer_0[1428] = ~(in[60] | in[3]); 
    assign layer_0[1429] = in[76] ^ in[74]; 
    assign layer_0[1430] = ~(in[139] ^ in[181]); 
    assign layer_0[1431] = ~(in[77] ^ in[23]); 
    assign layer_0[1432] = in[23]; 
    assign layer_0[1433] = ~(in[66] | in[53]); 
    assign layer_0[1434] = in[12] ^ in[70]; 
    assign layer_0[1435] = in[185] & ~in[206]; 
    assign layer_0[1436] = ~in[43]; 
    assign layer_0[1437] = in[163]; 
    assign layer_0[1438] = in[40] & ~in[155]; 
    assign layer_0[1439] = in[47] | in[0]; 
    assign layer_0[1440] = ~in[106] | (in[106] & in[111]); 
    assign layer_0[1441] = ~in[239] | (in[197] & in[239]); 
    assign layer_0[1442] = in[190]; 
    assign layer_0[1443] = in[239] & ~in[179]; 
    assign layer_0[1444] = in[27]; 
    assign layer_0[1445] = in[99] ^ in[29]; 
    assign layer_0[1446] = in[83] & ~in[87]; 
    assign layer_0[1447] = in[24] | in[39]; 
    assign layer_0[1448] = ~(in[157] & in[220]); 
    assign layer_0[1449] = in[119] & ~in[149]; 
    assign layer_0[1450] = ~in[126] | (in[173] & in[126]); 
    assign layer_0[1451] = in[143]; 
    assign layer_0[1452] = in[105]; 
    assign layer_0[1453] = in[118] & ~in[160]; 
    assign layer_0[1454] = in[200]; 
    assign layer_0[1455] = in[121] & ~in[65]; 
    assign layer_0[1456] = in[77] | in[189]; 
    assign layer_0[1457] = in[89]; 
    assign layer_0[1458] = ~(in[159] ^ in[57]); 
    assign layer_0[1459] = ~(in[40] & in[94]); 
    assign layer_0[1460] = ~(in[228] & in[114]); 
    assign layer_0[1461] = in[44] | in[64]; 
    assign layer_0[1462] = in[217] & in[250]; 
    assign layer_0[1463] = in[252] ^ in[211]; 
    assign layer_0[1464] = ~(in[208] & in[93]); 
    assign layer_0[1465] = in[197] & ~in[87]; 
    assign layer_0[1466] = in[252] & ~in[148]; 
    assign layer_0[1467] = in[161] & ~in[39]; 
    assign layer_0[1468] = in[95] | in[27]; 
    assign layer_0[1469] = ~in[38] | (in[38] & in[56]); 
    assign layer_0[1470] = ~in[86]; 
    assign layer_0[1471] = in[118]; 
    assign layer_0[1472] = in[91] & in[130]; 
    assign layer_0[1473] = in[201] & ~in[189]; 
    assign layer_0[1474] = in[104]; 
    assign layer_0[1475] = in[159] | in[139]; 
    assign layer_0[1476] = in[89]; 
    assign layer_0[1477] = in[202]; 
    assign layer_0[1478] = ~(in[125] ^ in[139]); 
    assign layer_0[1479] = ~(in[121] | in[202]); 
    assign layer_0[1480] = in[140] & ~in[97]; 
    assign layer_0[1481] = ~in[187] | (in[223] & in[187]); 
    assign layer_0[1482] = in[135] & ~in[243]; 
    assign layer_0[1483] = in[99] ^ in[37]; 
    assign layer_0[1484] = in[104] & ~in[3]; 
    assign layer_0[1485] = ~in[202]; 
    assign layer_0[1486] = ~in[108]; 
    assign layer_0[1487] = in[228] & ~in[174]; 
    assign layer_0[1488] = in[183]; 
    assign layer_0[1489] = ~(in[48] | in[134]); 
    assign layer_0[1490] = ~in[121] | (in[65] & in[121]); 
    assign layer_0[1491] = in[21] | in[13]; 
    assign layer_0[1492] = ~(in[84] & in[181]); 
    assign layer_0[1493] = in[231] & ~in[138]; 
    assign layer_0[1494] = in[162] & ~in[208]; 
    assign layer_0[1495] = in[147]; 
    assign layer_0[1496] = in[42]; 
    assign layer_0[1497] = ~(in[166] ^ in[118]); 
    assign layer_0[1498] = in[187]; 
    assign layer_0[1499] = in[142] ^ in[52]; 
    assign layer_0[1500] = in[172] & in[138]; 
    assign layer_0[1501] = in[158] | in[133]; 
    assign layer_0[1502] = in[74] ^ in[43]; 
    assign layer_0[1503] = in[214] ^ in[241]; 
    assign layer_0[1504] = in[66] ^ in[110]; 
    assign layer_0[1505] = in[30] ^ in[104]; 
    assign layer_0[1506] = ~in[232]; 
    assign layer_0[1507] = ~in[153]; 
    assign layer_0[1508] = ~in[215] | (in[215] & in[160]); 
    assign layer_0[1509] = ~in[53]; 
    assign layer_0[1510] = ~in[119] | (in[119] & in[81]); 
    assign layer_0[1511] = in[244] ^ in[227]; 
    assign layer_0[1512] = in[41] | in[117]; 
    assign layer_0[1513] = in[52] & in[139]; 
    assign layer_0[1514] = ~(in[23] & in[3]); 
    assign layer_0[1515] = ~in[47]; 
    assign layer_0[1516] = in[231]; 
    assign layer_0[1517] = in[28]; 
    assign layer_0[1518] = ~(in[158] ^ in[155]); 
    assign layer_0[1519] = ~in[40] | (in[12] & in[40]); 
    assign layer_0[1520] = in[211] & ~in[85]; 
    assign layer_0[1521] = ~in[172]; 
    assign layer_0[1522] = in[53]; 
    assign layer_0[1523] = ~(in[81] & in[48]); 
    assign layer_0[1524] = in[19]; 
    assign layer_0[1525] = in[201] | in[163]; 
    assign layer_0[1526] = in[103]; 
    assign layer_0[1527] = ~in[117]; 
    assign layer_0[1528] = ~in[132]; 
    assign layer_0[1529] = ~in[147] | (in[199] & in[147]); 
    assign layer_0[1530] = ~(in[90] & in[177]); 
    assign layer_0[1531] = ~in[248]; 
    assign layer_0[1532] = ~(in[170] ^ in[59]); 
    assign layer_0[1533] = in[152] & ~in[113]; 
    assign layer_0[1534] = ~in[75] | (in[21] & in[75]); 
    assign layer_0[1535] = ~in[77] | (in[77] & in[49]); 
    assign layer_0[1536] = ~in[91]; 
    assign layer_0[1537] = ~(in[5] ^ in[18]); 
    assign layer_0[1538] = in[73] ^ in[12]; 
    assign layer_0[1539] = ~(in[142] | in[65]); 
    assign layer_0[1540] = in[169] | in[138]; 
    assign layer_0[1541] = ~in[136] | (in[136] & in[208]); 
    assign layer_0[1542] = in[216] & ~in[111]; 
    assign layer_0[1543] = ~in[69]; 
    assign layer_0[1544] = in[119]; 
    assign layer_0[1545] = in[8] & ~in[125]; 
    assign layer_0[1546] = ~in[252]; 
    assign layer_0[1547] = in[64] | in[115]; 
    assign layer_0[1548] = ~in[81]; 
    assign layer_0[1549] = in[86] | in[122]; 
    assign layer_0[1550] = in[11] ^ in[67]; 
    assign layer_0[1551] = ~in[172]; 
    assign layer_0[1552] = in[39] ^ in[74]; 
    assign layer_0[1553] = ~(in[29] | in[46]); 
    assign layer_0[1554] = in[171] & ~in[144]; 
    assign layer_0[1555] = in[94]; 
    assign layer_0[1556] = ~in[186]; 
    assign layer_0[1557] = in[89] & ~in[31]; 
    assign layer_0[1558] = in[160] | in[249]; 
    assign layer_0[1559] = in[242] | in[205]; 
    assign layer_0[1560] = ~in[182] | (in[182] & in[176]); 
    assign layer_0[1561] = in[188] | in[181]; 
    assign layer_0[1562] = in[132] & ~in[37]; 
    assign layer_0[1563] = in[124] | in[100]; 
    assign layer_0[1564] = in[54]; 
    assign layer_0[1565] = in[49] ^ in[36]; 
    assign layer_0[1566] = in[94] & ~in[8]; 
    assign layer_0[1567] = ~(in[249] ^ in[223]); 
    assign layer_0[1568] = ~in[122]; 
    assign layer_0[1569] = in[125]; 
    assign layer_0[1570] = in[129]; 
    assign layer_0[1571] = in[121]; 
    assign layer_0[1572] = in[202] | in[174]; 
    assign layer_0[1573] = in[121] & in[185]; 
    assign layer_0[1574] = ~(in[90] | in[72]); 
    assign layer_0[1575] = in[110]; 
    assign layer_0[1576] = ~in[184] | (in[184] & in[166]); 
    assign layer_0[1577] = in[108]; 
    assign layer_0[1578] = in[240]; 
    assign layer_0[1579] = in[70]; 
    assign layer_0[1580] = in[220] ^ in[159]; 
    assign layer_0[1581] = ~in[92]; 
    assign layer_0[1582] = in[219] & ~in[162]; 
    assign layer_0[1583] = ~(in[188] | in[255]); 
    assign layer_0[1584] = ~(in[169] & in[122]); 
    assign layer_0[1585] = in[141] & ~in[170]; 
    assign layer_0[1586] = in[140] & in[148]; 
    assign layer_0[1587] = ~in[137]; 
    assign layer_0[1588] = ~in[174] | (in[222] & in[174]); 
    assign layer_0[1589] = ~(in[18] | in[121]); 
    assign layer_0[1590] = in[70] & ~in[143]; 
    assign layer_0[1591] = in[211] ^ in[115]; 
    assign layer_0[1592] = in[245] | in[250]; 
    assign layer_0[1593] = ~in[211]; 
    assign layer_0[1594] = in[142] & ~in[211]; 
    assign layer_0[1595] = in[39]; 
    assign layer_0[1596] = ~(in[125] | in[160]); 
    assign layer_0[1597] = in[168]; 
    assign layer_0[1598] = ~(in[104] ^ in[6]); 
    assign layer_0[1599] = ~in[137] | (in[137] & in[96]); 
    assign layer_0[1600] = in[133] & ~in[121]; 
    assign layer_0[1601] = ~(in[61] & in[142]); 
    assign layer_0[1602] = in[36] ^ in[90]; 
    assign layer_0[1603] = ~(in[56] & in[50]); 
    assign layer_0[1604] = ~in[62] | (in[160] & in[62]); 
    assign layer_0[1605] = ~in[242]; 
    assign layer_0[1606] = in[138]; 
    assign layer_0[1607] = in[121] & ~in[31]; 
    assign layer_0[1608] = ~(in[80] & in[38]); 
    assign layer_0[1609] = in[51]; 
    assign layer_0[1610] = in[25] ^ in[30]; 
    assign layer_0[1611] = ~in[56]; 
    assign layer_0[1612] = ~in[81]; 
    assign layer_0[1613] = ~(in[241] & in[160]); 
    assign layer_0[1614] = ~in[240] | (in[240] & in[139]); 
    assign layer_0[1615] = in[137] & ~in[246]; 
    assign layer_0[1616] = ~(in[152] | in[235]); 
    assign layer_0[1617] = ~in[95]; 
    assign layer_0[1618] = in[132] ^ in[162]; 
    assign layer_0[1619] = in[244] | in[247]; 
    assign layer_0[1620] = ~in[24] | (in[113] & in[24]); 
    assign layer_0[1621] = in[231]; 
    assign layer_0[1622] = ~in[44] | (in[44] & in[162]); 
    assign layer_0[1623] = ~(in[37] ^ in[87]); 
    assign layer_0[1624] = ~in[21]; 
    assign layer_0[1625] = in[191] & ~in[172]; 
    assign layer_0[1626] = in[138]; 
    assign layer_0[1627] = in[97] ^ in[101]; 
    assign layer_0[1628] = in[102] & ~in[50]; 
    assign layer_0[1629] = ~in[105] | (in[223] & in[105]); 
    assign layer_0[1630] = ~(in[248] & in[253]); 
    assign layer_0[1631] = in[213] ^ in[233]; 
    assign layer_0[1632] = in[195] | in[194]; 
    assign layer_0[1633] = in[198] & ~in[178]; 
    assign layer_0[1634] = ~in[247]; 
    assign layer_0[1635] = in[74] ^ in[117]; 
    assign layer_0[1636] = ~(in[251] ^ in[218]); 
    assign layer_0[1637] = in[116] & ~in[120]; 
    assign layer_0[1638] = in[189]; 
    assign layer_0[1639] = in[153] ^ in[173]; 
    assign layer_0[1640] = in[187]; 
    assign layer_0[1641] = in[136] & ~in[231]; 
    assign layer_0[1642] = ~in[217]; 
    assign layer_0[1643] = in[134]; 
    assign layer_0[1644] = in[254] ^ in[248]; 
    assign layer_0[1645] = ~in[174] | (in[189] & in[174]); 
    assign layer_0[1646] = in[105]; 
    assign layer_0[1647] = ~(in[18] | in[23]); 
    assign layer_0[1648] = ~in[141] | (in[60] & in[141]); 
    assign layer_0[1649] = in[214] & in[186]; 
    assign layer_0[1650] = ~in[233]; 
    assign layer_0[1651] = in[185] | in[182]; 
    assign layer_0[1652] = ~in[25] | (in[25] & in[128]); 
    assign layer_0[1653] = ~in[91]; 
    assign layer_0[1654] = ~(in[61] | in[84]); 
    assign layer_0[1655] = in[121] & ~in[16]; 
    assign layer_0[1656] = ~in[182]; 
    assign layer_0[1657] = ~in[169]; 
    assign layer_0[1658] = in[234] & ~in[136]; 
    assign layer_0[1659] = in[71] & ~in[52]; 
    assign layer_0[1660] = ~in[147]; 
    assign layer_0[1661] = in[14] & ~in[89]; 
    assign layer_0[1662] = ~(in[68] | in[58]); 
    assign layer_0[1663] = in[163] | in[222]; 
    assign layer_0[1664] = in[219] ^ in[215]; 
    assign layer_0[1665] = in[157] | in[197]; 
    assign layer_0[1666] = in[19] | in[64]; 
    assign layer_0[1667] = in[27] ^ in[85]; 
    assign layer_0[1668] = in[98] ^ in[37]; 
    assign layer_0[1669] = ~(in[28] & in[87]); 
    assign layer_0[1670] = ~in[217] | (in[217] & in[116]); 
    assign layer_0[1671] = ~in[245] | (in[245] & in[191]); 
    assign layer_0[1672] = ~(in[135] & in[106]); 
    assign layer_0[1673] = ~in[164]; 
    assign layer_0[1674] = in[120] & ~in[205]; 
    assign layer_0[1675] = in[16] ^ in[131]; 
    assign layer_0[1676] = in[49] & in[162]; 
    assign layer_0[1677] = in[115] & ~in[143]; 
    assign layer_0[1678] = in[236] | in[165]; 
    assign layer_0[1679] = in[211] | in[228]; 
    assign layer_0[1680] = in[201] & ~in[81]; 
    assign layer_0[1681] = in[13]; 
    assign layer_0[1682] = ~(in[64] & in[114]); 
    assign layer_0[1683] = in[140]; 
    assign layer_0[1684] = in[180] & ~in[164]; 
    assign layer_0[1685] = in[194]; 
    assign layer_0[1686] = in[4] | in[110]; 
    assign layer_0[1687] = ~(in[20] ^ in[42]); 
    assign layer_0[1688] = in[64] | in[41]; 
    assign layer_0[1689] = ~(in[202] | in[225]); 
    assign layer_0[1690] = ~(in[34] ^ in[141]); 
    assign layer_0[1691] = ~(in[93] ^ in[11]); 
    assign layer_0[1692] = in[235]; 
    assign layer_0[1693] = in[99]; 
    assign layer_0[1694] = ~(in[0] ^ in[64]); 
    assign layer_0[1695] = in[100]; 
    assign layer_0[1696] = ~in[38]; 
    assign layer_0[1697] = ~in[43] | (in[21] & in[43]); 
    assign layer_0[1698] = in[227] | in[234]; 
    assign layer_0[1699] = ~in[168]; 
    assign layer_0[1700] = ~in[225] | (in[183] & in[225]); 
    assign layer_0[1701] = in[148] & ~in[38]; 
    assign layer_0[1702] = in[219] ^ in[180]; 
    assign layer_0[1703] = ~in[155]; 
    assign layer_0[1704] = ~(in[5] ^ in[33]); 
    assign layer_0[1705] = in[54]; 
    assign layer_0[1706] = ~(in[86] | in[104]); 
    assign layer_0[1707] = in[48] & ~in[170]; 
    assign layer_0[1708] = ~(in[27] | in[114]); 
    assign layer_0[1709] = ~in[137]; 
    assign layer_0[1710] = ~in[64] | (in[174] & in[64]); 
    assign layer_0[1711] = in[85] | in[212]; 
    assign layer_0[1712] = ~(in[202] ^ in[117]); 
    assign layer_0[1713] = in[52] & ~in[22]; 
    assign layer_0[1714] = in[54] & ~in[40]; 
    assign layer_0[1715] = in[192]; 
    assign layer_0[1716] = in[21] ^ in[121]; 
    assign layer_0[1717] = ~in[83] | (in[83] & in[180]); 
    assign layer_0[1718] = ~(in[26] & in[94]); 
    assign layer_0[1719] = in[207]; 
    assign layer_0[1720] = in[136] & ~in[226]; 
    assign layer_0[1721] = ~in[92] | (in[92] & in[80]); 
    assign layer_0[1722] = ~(in[193] & in[228]); 
    assign layer_0[1723] = in[180]; 
    assign layer_0[1724] = ~(in[105] | in[146]); 
    assign layer_0[1725] = in[117]; 
    assign layer_0[1726] = ~(in[85] ^ in[0]); 
    assign layer_0[1727] = in[218] & in[165]; 
    assign layer_0[1728] = ~(in[4] & in[67]); 
    assign layer_0[1729] = in[172] | in[82]; 
    assign layer_0[1730] = in[216]; 
    assign layer_0[1731] = ~in[151] | (in[232] & in[151]); 
    assign layer_0[1732] = ~(in[12] | in[67]); 
    assign layer_0[1733] = in[127] & in[219]; 
    assign layer_0[1734] = in[122]; 
    assign layer_0[1735] = in[109] | in[6]; 
    assign layer_0[1736] = ~in[90] | (in[12] & in[90]); 
    assign layer_0[1737] = in[204] & ~in[84]; 
    assign layer_0[1738] = ~in[84] | (in[84] & in[202]); 
    assign layer_0[1739] = in[251] & ~in[208]; 
    assign layer_0[1740] = ~in[141]; 
    assign layer_0[1741] = in[31] & in[59]; 
    assign layer_0[1742] = in[169] & ~in[196]; 
    assign layer_0[1743] = ~in[177] | (in[177] & in[54]); 
    assign layer_0[1744] = ~(in[126] ^ in[89]); 
    assign layer_0[1745] = in[167] & in[40]; 
    assign layer_0[1746] = in[214] ^ in[146]; 
    assign layer_0[1747] = ~in[149] | (in[78] & in[149]); 
    assign layer_0[1748] = ~in[171] | (in[81] & in[171]); 
    assign layer_0[1749] = in[25]; 
    assign layer_0[1750] = in[254]; 
    assign layer_0[1751] = in[120] ^ in[165]; 
    assign layer_0[1752] = ~(in[223] ^ in[162]); 
    assign layer_0[1753] = in[70] & ~in[34]; 
    assign layer_0[1754] = in[72]; 
    assign layer_0[1755] = ~in[187]; 
    assign layer_0[1756] = in[36] ^ in[55]; 
    assign layer_0[1757] = ~in[236]; 
    assign layer_0[1758] = ~(in[84] & in[153]); 
    assign layer_0[1759] = ~in[236]; 
    assign layer_0[1760] = in[238] | in[203]; 
    assign layer_0[1761] = ~(in[140] ^ in[216]); 
    assign layer_0[1762] = in[45] | in[100]; 
    assign layer_0[1763] = in[239] | in[197]; 
    assign layer_0[1764] = in[91] ^ in[3]; 
    assign layer_0[1765] = in[211] ^ in[142]; 
    assign layer_0[1766] = ~(in[214] | in[194]); 
    assign layer_0[1767] = in[24] ^ in[138]; 
    assign layer_0[1768] = ~(in[176] ^ in[225]); 
    assign layer_0[1769] = ~in[123]; 
    assign layer_0[1770] = in[6] & in[79]; 
    assign layer_0[1771] = in[54] & in[112]; 
    assign layer_0[1772] = in[201] | in[79]; 
    assign layer_0[1773] = in[70] & ~in[108]; 
    assign layer_0[1774] = ~(in[170] ^ in[150]); 
    assign layer_0[1775] = in[69]; 
    assign layer_0[1776] = ~in[175] | (in[222] & in[175]); 
    assign layer_0[1777] = in[154]; 
    assign layer_0[1778] = in[241] | in[126]; 
    assign layer_0[1779] = ~(in[152] | in[51]); 
    assign layer_0[1780] = ~in[136]; 
    assign layer_0[1781] = ~in[124]; 
    assign layer_0[1782] = ~in[127] | (in[127] & in[192]); 
    assign layer_0[1783] = ~(in[43] | in[171]); 
    assign layer_0[1784] = ~in[159]; 
    assign layer_0[1785] = ~in[121]; 
    assign layer_0[1786] = ~in[45] | (in[45] & in[144]); 
    assign layer_0[1787] = in[254]; 
    assign layer_0[1788] = ~in[190] | (in[94] & in[190]); 
    assign layer_0[1789] = ~in[110] | (in[8] & in[110]); 
    assign layer_0[1790] = ~in[239] | (in[223] & in[239]); 
    assign layer_0[1791] = in[180] & ~in[62]; 
    assign layer_0[1792] = ~in[124]; 
    assign layer_0[1793] = ~in[85] | (in[85] & in[107]); 
    assign layer_0[1794] = ~in[88] | (in[33] & in[88]); 
    assign layer_0[1795] = ~(in[240] ^ in[144]); 
    assign layer_0[1796] = in[168]; 
    assign layer_0[1797] = in[8]; 
    assign layer_0[1798] = in[174]; 
    assign layer_0[1799] = in[176] & in[81]; 
    assign layer_0[1800] = ~(in[154] ^ in[209]); 
    assign layer_0[1801] = in[229]; 
    assign layer_0[1802] = in[118]; 
    assign layer_0[1803] = ~(in[133] | in[221]); 
    assign layer_0[1804] = ~(in[10] & in[73]); 
    assign layer_0[1805] = in[124] & ~in[19]; 
    assign layer_0[1806] = in[178] & in[59]; 
    assign layer_0[1807] = ~(in[12] ^ in[46]); 
    assign layer_0[1808] = in[106] | in[196]; 
    assign layer_0[1809] = ~(in[4] ^ in[80]); 
    assign layer_0[1810] = ~in[126]; 
    assign layer_0[1811] = ~(in[168] ^ in[202]); 
    assign layer_0[1812] = ~in[129] | (in[129] & in[234]); 
    assign layer_0[1813] = ~in[133]; 
    assign layer_0[1814] = ~(in[48] | in[170]); 
    assign layer_0[1815] = in[202] ^ in[75]; 
    assign layer_0[1816] = ~in[166]; 
    assign layer_0[1817] = ~in[218] | (in[250] & in[218]); 
    assign layer_0[1818] = in[219] | in[161]; 
    assign layer_0[1819] = ~in[238] | (in[223] & in[238]); 
    assign layer_0[1820] = ~in[152] | (in[249] & in[152]); 
    assign layer_0[1821] = ~in[181] | (in[240] & in[181]); 
    assign layer_0[1822] = ~(in[225] | in[184]); 
    assign layer_0[1823] = ~in[161]; 
    assign layer_0[1824] = ~in[42] | (in[42] & in[162]); 
    assign layer_0[1825] = ~in[221]; 
    assign layer_0[1826] = ~(in[67] | in[24]); 
    assign layer_0[1827] = ~in[132]; 
    assign layer_0[1828] = ~in[70] | (in[60] & in[70]); 
    assign layer_0[1829] = in[46] & in[92]; 
    assign layer_0[1830] = in[39]; 
    assign layer_0[1831] = ~(in[91] & in[71]); 
    assign layer_0[1832] = ~(in[199] & in[123]); 
    assign layer_0[1833] = in[189] ^ in[93]; 
    assign layer_0[1834] = ~in[27] | (in[8] & in[27]); 
    assign layer_0[1835] = in[36] | in[104]; 
    assign layer_0[1836] = ~in[108]; 
    assign layer_0[1837] = in[107] & ~in[223]; 
    assign layer_0[1838] = ~(in[248] ^ in[242]); 
    assign layer_0[1839] = in[174] ^ in[82]; 
    assign layer_0[1840] = in[157] | in[122]; 
    assign layer_0[1841] = ~(in[122] & in[61]); 
    assign layer_0[1842] = ~in[214] | (in[214] & in[242]); 
    assign layer_0[1843] = ~(in[59] ^ in[138]); 
    assign layer_0[1844] = ~in[170]; 
    assign layer_0[1845] = in[101] & ~in[45]; 
    assign layer_0[1846] = in[128] & ~in[117]; 
    assign layer_0[1847] = in[119]; 
    assign layer_0[1848] = ~(in[56] | in[100]); 
    assign layer_0[1849] = in[189]; 
    assign layer_0[1850] = in[82]; 
    assign layer_0[1851] = in[74] & ~in[35]; 
    assign layer_0[1852] = ~(in[224] | in[168]); 
    assign layer_0[1853] = ~(in[70] ^ in[114]); 
    assign layer_0[1854] = in[171] & in[223]; 
    assign layer_0[1855] = in[252] | in[229]; 
    assign layer_0[1856] = ~in[149] | (in[198] & in[149]); 
    assign layer_0[1857] = in[235] ^ in[122]; 
    assign layer_0[1858] = in[99] & ~in[14]; 
    assign layer_0[1859] = ~in[131] | (in[176] & in[131]); 
    assign layer_0[1860] = ~(in[252] | in[154]); 
    assign layer_0[1861] = in[198] & ~in[248]; 
    assign layer_0[1862] = in[104] & ~in[101]; 
    assign layer_0[1863] = in[49] ^ in[80]; 
    assign layer_0[1864] = in[18] & in[62]; 
    assign layer_0[1865] = ~in[85]; 
    assign layer_0[1866] = ~(in[97] ^ in[94]); 
    assign layer_0[1867] = ~in[114]; 
    assign layer_0[1868] = in[196] ^ in[173]; 
    assign layer_0[1869] = ~(in[92] | in[75]); 
    assign layer_0[1870] = ~(in[239] ^ in[202]); 
    assign layer_0[1871] = in[43] & ~in[4]; 
    assign layer_0[1872] = in[137]; 
    assign layer_0[1873] = in[254] | in[172]; 
    assign layer_0[1874] = in[53] | in[16]; 
    assign layer_0[1875] = in[5] & ~in[84]; 
    assign layer_0[1876] = ~in[186] | (in[186] & in[175]); 
    assign layer_0[1877] = ~in[170]; 
    assign layer_0[1878] = in[123]; 
    assign layer_0[1879] = in[68]; 
    assign layer_0[1880] = ~in[36]; 
    assign layer_0[1881] = in[44]; 
    assign layer_0[1882] = ~in[49]; 
    assign layer_0[1883] = in[155] & in[38]; 
    assign layer_0[1884] = ~in[249]; 
    assign layer_0[1885] = ~in[42] | (in[42] & in[49]); 
    assign layer_0[1886] = in[213] & in[254]; 
    assign layer_0[1887] = ~(in[86] & in[185]); 
    assign layer_0[1888] = in[204] | in[239]; 
    assign layer_0[1889] = ~in[197] | (in[197] & in[229]); 
    assign layer_0[1890] = in[52] | in[1]; 
    assign layer_0[1891] = ~in[74] | (in[74] & in[48]); 
    assign layer_0[1892] = in[247] | in[248]; 
    assign layer_0[1893] = in[56] & in[160]; 
    assign layer_0[1894] = in[65] | in[105]; 
    assign layer_0[1895] = in[134] & ~in[37]; 
    assign layer_0[1896] = in[28] & in[51]; 
    assign layer_0[1897] = ~(in[65] & in[85]); 
    assign layer_0[1898] = in[243] | in[246]; 
    assign layer_0[1899] = in[213] & ~in[236]; 
    assign layer_0[1900] = ~(in[231] ^ in[228]); 
    assign layer_0[1901] = in[148] | in[44]; 
    assign layer_0[1902] = in[194]; 
    assign layer_0[1903] = in[195] ^ in[111]; 
    assign layer_0[1904] = in[151] ^ in[167]; 
    assign layer_0[1905] = ~in[171]; 
    assign layer_0[1906] = in[211] ^ in[169]; 
    assign layer_0[1907] = in[162] & ~in[237]; 
    assign layer_0[1908] = ~(in[12] | in[131]); 
    assign layer_0[1909] = in[170] | in[201]; 
    assign layer_0[1910] = ~in[140] | (in[195] & in[140]); 
    assign layer_0[1911] = ~in[244] | (in[223] & in[244]); 
    assign layer_0[1912] = ~in[61] | (in[31] & in[61]); 
    assign layer_0[1913] = ~in[43] | (in[43] & in[93]); 
    assign layer_0[1914] = ~(in[9] | in[27]); 
    assign layer_0[1915] = ~in[154]; 
    assign layer_0[1916] = ~in[6]; 
    assign layer_0[1917] = in[29]; 
    assign layer_0[1918] = in[225] | in[249]; 
    assign layer_0[1919] = ~in[107]; 
    assign layer_0[1920] = ~in[165]; 
    assign layer_0[1921] = ~in[107] | (in[43] & in[107]); 
    assign layer_0[1922] = in[252] | in[231]; 
    assign layer_0[1923] = in[4] ^ in[63]; 
    assign layer_0[1924] = ~in[122]; 
    assign layer_0[1925] = in[88] | in[97]; 
    assign layer_0[1926] = ~in[168]; 
    assign layer_0[1927] = ~(in[145] & in[144]); 
    assign layer_0[1928] = in[100] | in[120]; 
    assign layer_0[1929] = in[248] ^ in[237]; 
    assign layer_0[1930] = ~in[201]; 
    assign layer_0[1931] = ~in[166]; 
    assign layer_0[1932] = in[8] | in[134]; 
    assign layer_0[1933] = ~(in[192] & in[81]); 
    assign layer_0[1934] = in[85]; 
    assign layer_0[1935] = in[50] & ~in[79]; 
    assign layer_0[1936] = ~(in[214] ^ in[216]); 
    assign layer_0[1937] = in[42] ^ in[142]; 
    assign layer_0[1938] = ~in[59]; 
    assign layer_0[1939] = in[108]; 
    assign layer_0[1940] = ~in[104] | (in[36] & in[104]); 
    assign layer_0[1941] = ~in[104] | (in[104] & in[96]); 
    assign layer_0[1942] = ~in[173]; 
    assign layer_0[1943] = ~in[150] | (in[208] & in[150]); 
    assign layer_0[1944] = ~(in[149] ^ in[201]); 
    assign layer_0[1945] = in[237] ^ in[239]; 
    assign layer_0[1946] = ~(in[226] | in[250]); 
    assign layer_0[1947] = ~(in[57] & in[168]); 
    assign layer_0[1948] = ~(in[232] ^ in[226]); 
    assign layer_0[1949] = ~in[151] | (in[151] & in[127]); 
    assign layer_0[1950] = in[218] ^ in[246]; 
    assign layer_0[1951] = in[75] & ~in[191]; 
    assign layer_0[1952] = ~(in[139] & in[62]); 
    assign layer_0[1953] = ~(in[242] & in[224]); 
    assign layer_0[1954] = ~(in[130] & in[141]); 
    assign layer_0[1955] = in[210]; 
    assign layer_0[1956] = ~in[119]; 
    assign layer_0[1957] = ~in[64] | (in[64] & in[173]); 
    assign layer_0[1958] = in[161] | in[255]; 
    assign layer_0[1959] = in[149]; 
    assign layer_0[1960] = in[243]; 
    assign layer_0[1961] = in[102] & ~in[230]; 
    assign layer_0[1962] = ~in[70] | (in[70] & in[62]); 
    assign layer_0[1963] = in[20] | in[83]; 
    assign layer_0[1964] = ~in[201] | (in[159] & in[201]); 
    assign layer_0[1965] = ~in[239] | (in[239] & in[243]); 
    assign layer_0[1966] = in[146]; 
    assign layer_0[1967] = in[239] | in[198]; 
    assign layer_0[1968] = in[231] | in[251]; 
    assign layer_0[1969] = ~(in[188] | in[102]); 
    assign layer_0[1970] = ~in[196]; 
    assign layer_0[1971] = ~(in[170] | in[177]); 
    assign layer_0[1972] = in[4]; 
    assign layer_0[1973] = in[171]; 
    assign layer_0[1974] = ~in[175] | (in[175] & in[159]); 
    assign layer_0[1975] = ~in[136]; 
    assign layer_0[1976] = ~in[176]; 
    assign layer_0[1977] = in[153] | in[50]; 
    assign layer_0[1978] = in[125] & ~in[15]; 
    assign layer_0[1979] = in[154] & in[74]; 
    assign layer_0[1980] = in[93] | in[200]; 
    assign layer_0[1981] = in[164] & ~in[250]; 
    assign layer_0[1982] = in[235] | in[183]; 
    assign layer_0[1983] = in[116]; 
    assign layer_0[1984] = ~in[40]; 
    assign layer_0[1985] = ~(in[239] | in[185]); 
    assign layer_0[1986] = ~(in[195] & in[109]); 
    assign layer_0[1987] = in[131] & ~in[85]; 
    assign layer_0[1988] = in[103] & ~in[9]; 
    assign layer_0[1989] = ~in[159] | (in[50] & in[159]); 
    assign layer_0[1990] = ~in[107]; 
    assign layer_0[1991] = in[11] ^ in[68]; 
    assign layer_0[1992] = in[137] & in[40]; 
    assign layer_0[1993] = ~(in[198] & in[171]); 
    assign layer_0[1994] = in[221] & in[209]; 
    assign layer_0[1995] = in[3] & in[48]; 
    assign layer_0[1996] = ~in[151]; 
    assign layer_0[1997] = ~(in[26] & in[51]); 
    assign layer_0[1998] = ~in[86] | (in[86] & in[23]); 
    assign layer_0[1999] = in[103] & ~in[19]; 
    assign layer_0[2000] = ~in[40]; 
    assign layer_0[2001] = in[112] | in[193]; 
    assign layer_0[2002] = in[156]; 
    assign layer_0[2003] = in[85]; 
    assign layer_0[2004] = in[229]; 
    assign layer_0[2005] = in[185] | in[68]; 
    assign layer_0[2006] = ~(in[101] ^ in[214]); 
    assign layer_0[2007] = in[23] ^ in[18]; 
    assign layer_0[2008] = ~(in[24] ^ in[142]); 
    assign layer_0[2009] = in[141] & ~in[225]; 
    assign layer_0[2010] = ~(in[47] ^ in[30]); 
    assign layer_0[2011] = ~(in[118] & in[91]); 
    assign layer_0[2012] = in[25] ^ in[8]; 
    assign layer_0[2013] = in[197] | in[208]; 
    assign layer_0[2014] = ~(in[55] & in[120]); 
    assign layer_0[2015] = in[90] & ~in[76]; 
    assign layer_0[2016] = ~(in[242] ^ in[210]); 
    assign layer_0[2017] = in[211]; 
    assign layer_0[2018] = ~(in[110] | in[155]); 
    assign layer_0[2019] = ~(in[137] & in[29]); 
    assign layer_0[2020] = ~(in[65] ^ in[169]); 
    assign layer_0[2021] = in[9] & ~in[82]; 
    assign layer_0[2022] = ~(in[243] | in[245]); 
    assign layer_0[2023] = ~in[39] | (in[39] & in[26]); 
    assign layer_0[2024] = in[87]; 
    assign layer_0[2025] = in[3] & ~in[27]; 
    assign layer_0[2026] = in[135] | in[61]; 
    assign layer_0[2027] = ~in[168]; 
    assign layer_0[2028] = ~(in[93] | in[40]); 
    assign layer_0[2029] = in[147]; 
    assign layer_0[2030] = ~in[220] | (in[220] & in[224]); 
    assign layer_0[2031] = in[4] ^ in[90]; 
    assign layer_0[2032] = in[195] & ~in[143]; 
    assign layer_0[2033] = ~in[35]; 
    assign layer_0[2034] = ~in[74]; 
    assign layer_0[2035] = in[0]; 
    assign layer_0[2036] = ~in[201] | (in[134] & in[201]); 
    assign layer_0[2037] = ~(in[61] | in[167]); 
    assign layer_0[2038] = ~in[142] | (in[228] & in[142]); 
    assign layer_0[2039] = ~(in[73] | in[109]); 
    assign layer_0[2040] = in[26] | in[62]; 
    assign layer_0[2041] = ~(in[106] ^ in[160]); 
    assign layer_0[2042] = ~in[170] | (in[76] & in[170]); 
    assign layer_0[2043] = ~(in[177] ^ in[57]); 
    assign layer_0[2044] = in[139]; 
    assign layer_0[2045] = ~(in[238] ^ in[111]); 
    assign layer_0[2046] = in[177] ^ in[107]; 
    assign layer_0[2047] = ~(in[214] ^ in[203]); 
    assign layer_0[2048] = in[254]; 
    assign layer_0[2049] = ~in[152] | (in[152] & in[172]); 
    assign layer_0[2050] = ~(in[17] & in[65]); 
    assign layer_0[2051] = ~in[172] | (in[191] & in[172]); 
    assign layer_0[2052] = ~in[127]; 
    assign layer_0[2053] = in[247] & ~in[235]; 
    assign layer_0[2054] = in[221]; 
    assign layer_0[2055] = ~(in[85] | in[90]); 
    assign layer_0[2056] = ~in[101]; 
    assign layer_0[2057] = ~(in[16] ^ in[138]); 
    assign layer_0[2058] = ~(in[90] | in[96]); 
    assign layer_0[2059] = in[202] & ~in[123]; 
    assign layer_0[2060] = ~in[165]; 
    assign layer_0[2061] = in[188] | in[62]; 
    assign layer_0[2062] = ~in[242]; 
    assign layer_0[2063] = in[100] | in[183]; 
    assign layer_0[2064] = ~in[135] | (in[28] & in[135]); 
    assign layer_0[2065] = ~(in[171] & in[172]); 
    assign layer_0[2066] = ~(in[218] & in[151]); 
    assign layer_0[2067] = ~(in[185] | in[201]); 
    assign layer_0[2068] = ~in[124]; 
    assign layer_0[2069] = in[237] & ~in[189]; 
    assign layer_0[2070] = in[43]; 
    assign layer_0[2071] = in[36] | in[25]; 
    assign layer_0[2072] = in[62] | in[84]; 
    assign layer_0[2073] = ~in[146]; 
    assign layer_0[2074] = in[22]; 
    assign layer_0[2075] = ~(in[91] | in[159]); 
    assign layer_0[2076] = ~in[39]; 
    assign layer_0[2077] = in[166]; 
    assign layer_0[2078] = in[28] & in[0]; 
    assign layer_0[2079] = in[125]; 
    assign layer_0[2080] = ~in[114]; 
    assign layer_0[2081] = ~in[121]; 
    assign layer_0[2082] = in[164] ^ in[166]; 
    assign layer_0[2083] = ~in[244] | (in[129] & in[244]); 
    assign layer_0[2084] = in[19] & ~in[23]; 
    assign layer_0[2085] = ~(in[199] | in[231]); 
    assign layer_0[2086] = in[61] ^ in[159]; 
    assign layer_0[2087] = in[154] ^ in[108]; 
    assign layer_0[2088] = ~in[109]; 
    assign layer_0[2089] = ~(in[241] ^ in[175]); 
    assign layer_0[2090] = ~(in[123] ^ in[17]); 
    assign layer_0[2091] = in[100] | in[225]; 
    assign layer_0[2092] = ~in[100]; 
    assign layer_0[2093] = ~in[129]; 
    assign layer_0[2094] = ~in[100]; 
    assign layer_0[2095] = ~(in[105] ^ in[150]); 
    assign layer_0[2096] = in[11] & ~in[68]; 
    assign layer_0[2097] = ~(in[104] | in[145]); 
    assign layer_0[2098] = ~(in[170] | in[168]); 
    assign layer_0[2099] = in[183] & ~in[118]; 
    assign layer_0[2100] = ~in[137]; 
    assign layer_0[2101] = in[30] | in[57]; 
    assign layer_0[2102] = in[153] & ~in[163]; 
    assign layer_0[2103] = in[197] ^ in[201]; 
    assign layer_0[2104] = in[183]; 
    assign layer_0[2105] = in[203] | in[131]; 
    assign layer_0[2106] = ~in[4] | (in[12] & in[4]); 
    assign layer_0[2107] = ~(in[191] ^ in[246]); 
    assign layer_0[2108] = ~(in[227] ^ in[144]); 
    assign layer_0[2109] = ~(in[15] & in[47]); 
    assign layer_0[2110] = ~in[70]; 
    assign layer_0[2111] = ~in[243]; 
    assign layer_0[2112] = ~(in[21] | in[121]); 
    assign layer_0[2113] = in[149] & ~in[58]; 
    assign layer_0[2114] = ~(in[171] | in[76]); 
    assign layer_0[2115] = ~(in[208] ^ in[159]); 
    assign layer_0[2116] = in[251] ^ in[186]; 
    assign layer_0[2117] = ~in[85] | (in[30] & in[85]); 
    assign layer_0[2118] = in[21]; 
    assign layer_0[2119] = ~(in[196] & in[121]); 
    assign layer_0[2120] = ~(in[140] ^ in[135]); 
    assign layer_0[2121] = ~in[39]; 
    assign layer_0[2122] = ~(in[19] | in[97]); 
    assign layer_0[2123] = ~in[22] | (in[41] & in[22]); 
    assign layer_0[2124] = ~in[30] | (in[52] & in[30]); 
    assign layer_0[2125] = in[14] & ~in[0]; 
    assign layer_0[2126] = ~(in[73] | in[14]); 
    assign layer_0[2127] = ~in[6] | (in[69] & in[6]); 
    assign layer_0[2128] = in[28] & ~in[83]; 
    assign layer_0[2129] = ~in[11] | (in[11] & in[55]); 
    assign layer_0[2130] = in[224]; 
    assign layer_0[2131] = ~in[161] | (in[62] & in[161]); 
    assign layer_0[2132] = in[230] | in[116]; 
    assign layer_0[2133] = in[0] ^ in[86]; 
    assign layer_0[2134] = ~(in[249] | in[155]); 
    assign layer_0[2135] = in[25] ^ in[17]; 
    assign layer_0[2136] = in[154] & ~in[49]; 
    assign layer_0[2137] = ~(in[28] ^ in[82]); 
    assign layer_0[2138] = in[219]; 
    assign layer_0[2139] = ~(in[37] ^ in[48]); 
    assign layer_0[2140] = ~in[178] | (in[244] & in[178]); 
    assign layer_0[2141] = in[218] ^ in[234]; 
    assign layer_0[2142] = in[10] | in[72]; 
    assign layer_0[2143] = ~(in[243] | in[159]); 
    assign layer_0[2144] = in[25] & ~in[72]; 
    assign layer_0[2145] = in[17] ^ in[136]; 
    assign layer_0[2146] = in[185]; 
    assign layer_0[2147] = ~(in[90] | in[21]); 
    assign layer_0[2148] = ~in[215]; 
    assign layer_0[2149] = ~in[136] | (in[8] & in[136]); 
    assign layer_0[2150] = ~in[135]; 
    assign layer_0[2151] = in[59]; 
    assign layer_0[2152] = ~(in[110] ^ in[202]); 
    assign layer_0[2153] = in[117]; 
    assign layer_0[2154] = in[238] & in[210]; 
    assign layer_0[2155] = in[205] | in[147]; 
    assign layer_0[2156] = in[11] ^ in[69]; 
    assign layer_0[2157] = ~in[139]; 
    assign layer_0[2158] = ~in[177] | (in[177] & in[192]); 
    assign layer_0[2159] = in[155] | in[28]; 
    assign layer_0[2160] = in[124] & ~in[232]; 
    assign layer_0[2161] = in[221] & ~in[195]; 
    assign layer_0[2162] = in[63] & in[160]; 
    assign layer_0[2163] = in[47]; 
    assign layer_0[2164] = ~(in[178] & in[174]); 
    assign layer_0[2165] = ~(in[134] | in[9]); 
    assign layer_0[2166] = ~(in[139] | in[66]); 
    assign layer_0[2167] = in[53]; 
    assign layer_0[2168] = in[43]; 
    assign layer_0[2169] = ~in[133] | (in[63] & in[133]); 
    assign layer_0[2170] = in[103]; 
    assign layer_0[2171] = in[109]; 
    assign layer_0[2172] = ~in[105] | (in[205] & in[105]); 
    assign layer_0[2173] = ~in[50] | (in[50] & in[176]); 
    assign layer_0[2174] = ~in[158]; 
    assign layer_0[2175] = ~(in[235] | in[213]); 
    assign layer_0[2176] = ~(in[219] | in[152]); 
    assign layer_0[2177] = in[105] & ~in[212]; 
    assign layer_0[2178] = in[85] ^ in[87]; 
    assign layer_0[2179] = ~in[68] | (in[68] & in[37]); 
    assign layer_0[2180] = ~in[187]; 
    assign layer_0[2181] = in[197] | in[205]; 
    assign layer_0[2182] = ~in[169]; 
    assign layer_0[2183] = ~(in[95] & in[152]); 
    assign layer_0[2184] = ~in[99]; 
    assign layer_0[2185] = ~in[186] | (in[186] & in[210]); 
    assign layer_0[2186] = in[104] & ~in[188]; 
    assign layer_0[2187] = in[226] | in[114]; 
    assign layer_0[2188] = ~(in[183] ^ in[215]); 
    assign layer_0[2189] = in[200] ^ in[141]; 
    assign layer_0[2190] = in[230] & in[193]; 
    assign layer_0[2191] = ~in[167] | (in[175] & in[167]); 
    assign layer_0[2192] = in[198]; 
    assign layer_0[2193] = in[46] | in[129]; 
    assign layer_0[2194] = ~(in[119] | in[34]); 
    assign layer_0[2195] = ~in[124]; 
    assign layer_0[2196] = in[170] & in[91]; 
    assign layer_0[2197] = in[134]; 
    assign layer_0[2198] = in[58] | in[77]; 
    assign layer_0[2199] = in[138] & ~in[111]; 
    assign layer_0[2200] = in[123] & ~in[184]; 
    assign layer_0[2201] = ~in[42] | (in[42] & in[104]); 
    assign layer_0[2202] = in[176] | in[180]; 
    assign layer_0[2203] = ~in[80]; 
    assign layer_0[2204] = ~in[139] | (in[253] & in[139]); 
    assign layer_0[2205] = ~in[90] | (in[112] & in[90]); 
    assign layer_0[2206] = ~in[66]; 
    assign layer_0[2207] = in[114]; 
    assign layer_0[2208] = ~in[154] | (in[154] & in[165]); 
    assign layer_0[2209] = in[133] & ~in[234]; 
    assign layer_0[2210] = in[3] | in[123]; 
    assign layer_0[2211] = in[218] & ~in[134]; 
    assign layer_0[2212] = ~in[216]; 
    assign layer_0[2213] = ~in[175] | (in[110] & in[175]); 
    assign layer_0[2214] = in[188] & ~in[242]; 
    assign layer_0[2215] = ~(in[36] ^ in[7]); 
    assign layer_0[2216] = in[136]; 
    assign layer_0[2217] = in[141] & ~in[143]; 
    assign layer_0[2218] = in[40] ^ in[122]; 
    assign layer_0[2219] = ~(in[106] | in[127]); 
    assign layer_0[2220] = in[53] ^ in[12]; 
    assign layer_0[2221] = ~(in[231] | in[161]); 
    assign layer_0[2222] = in[200] & ~in[127]; 
    assign layer_0[2223] = ~(in[176] | in[153]); 
    assign layer_0[2224] = ~in[55]; 
    assign layer_0[2225] = ~(in[187] & in[68]); 
    assign layer_0[2226] = in[140]; 
    assign layer_0[2227] = in[150] | in[58]; 
    assign layer_0[2228] = ~in[123]; 
    assign layer_0[2229] = in[8]; 
    assign layer_0[2230] = ~(in[171] | in[196]); 
    assign layer_0[2231] = in[92] | in[138]; 
    assign layer_0[2232] = ~(in[45] ^ in[133]); 
    assign layer_0[2233] = in[4]; 
    assign layer_0[2234] = ~(in[32] & in[59]); 
    assign layer_0[2235] = ~in[168] | (in[246] & in[168]); 
    assign layer_0[2236] = ~in[35] | (in[109] & in[35]); 
    assign layer_0[2237] = ~in[143]; 
    assign layer_0[2238] = ~in[197]; 
    assign layer_0[2239] = in[155]; 
    assign layer_0[2240] = ~in[1]; 
    assign layer_0[2241] = ~in[154] | (in[154] & in[28]); 
    assign layer_0[2242] = ~in[16] | (in[2] & in[16]); 
    assign layer_0[2243] = ~in[49] | (in[124] & in[49]); 
    assign layer_0[2244] = ~in[160] | (in[254] & in[160]); 
    assign layer_0[2245] = ~in[111]; 
    assign layer_0[2246] = ~(in[193] ^ in[123]); 
    assign layer_0[2247] = ~in[54] | (in[54] & in[64]); 
    assign layer_0[2248] = in[96] | in[25]; 
    assign layer_0[2249] = ~(in[27] ^ in[73]); 
    assign layer_0[2250] = ~(in[175] ^ in[197]); 
    assign layer_0[2251] = ~(in[74] & in[57]); 
    assign layer_0[2252] = ~in[36]; 
    assign layer_0[2253] = ~(in[168] & in[85]); 
    assign layer_0[2254] = ~(in[83] ^ in[86]); 
    assign layer_0[2255] = in[13] | in[107]; 
    assign layer_0[2256] = ~(in[138] ^ in[193]); 
    assign layer_0[2257] = in[224] & in[148]; 
    assign layer_0[2258] = ~in[76] | (in[76] & in[111]); 
    assign layer_0[2259] = ~in[209]; 
    assign layer_0[2260] = in[221]; 
    assign layer_0[2261] = ~in[57] | (in[57] & in[23]); 
    assign layer_0[2262] = ~in[251] | (in[141] & in[251]); 
    assign layer_0[2263] = ~in[114]; 
    assign layer_0[2264] = in[37]; 
    assign layer_0[2265] = ~(in[180] ^ in[103]); 
    assign layer_0[2266] = ~(in[208] ^ in[90]); 
    assign layer_0[2267] = in[43] | in[146]; 
    assign layer_0[2268] = ~in[219] | (in[130] & in[219]); 
    assign layer_0[2269] = ~in[131]; 
    assign layer_0[2270] = ~in[150] | (in[189] & in[150]); 
    assign layer_0[2271] = in[57] ^ in[140]; 
    assign layer_0[2272] = ~in[80]; 
    assign layer_0[2273] = in[101] & ~in[191]; 
    assign layer_0[2274] = in[78] ^ in[127]; 
    assign layer_0[2275] = ~in[246]; 
    assign layer_0[2276] = ~in[158]; 
    assign layer_0[2277] = ~in[39] | (in[54] & in[39]); 
    assign layer_0[2278] = in[120] | in[159]; 
    assign layer_0[2279] = in[83] & ~in[137]; 
    assign layer_0[2280] = in[164] ^ in[224]; 
    assign layer_0[2281] = ~in[255] | (in[139] & in[255]); 
    assign layer_0[2282] = in[109] | in[7]; 
    assign layer_0[2283] = in[208] & in[143]; 
    assign layer_0[2284] = in[1]; 
    assign layer_0[2285] = ~in[101]; 
    assign layer_0[2286] = in[134] | in[221]; 
    assign layer_0[2287] = ~(in[72] ^ in[113]); 
    assign layer_0[2288] = ~in[43]; 
    assign layer_0[2289] = ~in[105]; 
    assign layer_0[2290] = in[152] & in[57]; 
    assign layer_0[2291] = in[21] ^ in[127]; 
    assign layer_0[2292] = ~(in[178] | in[195]); 
    assign layer_0[2293] = in[90] & ~in[207]; 
    assign layer_0[2294] = in[101] & in[71]; 
    assign layer_0[2295] = in[16] | in[67]; 
    assign layer_0[2296] = in[96] | in[87]; 
    assign layer_0[2297] = in[184] ^ in[95]; 
    assign layer_0[2298] = ~(in[157] | in[237]); 
    assign layer_0[2299] = ~in[74]; 
    assign layer_0[2300] = in[161]; 
    assign layer_0[2301] = ~in[240]; 
    assign layer_0[2302] = in[242] & ~in[169]; 
    assign layer_0[2303] = in[129] ^ in[24]; 
    assign layer_0[2304] = in[123] & in[211]; 
    assign layer_0[2305] = ~(in[141] | in[110]); 
    assign layer_0[2306] = ~(in[76] ^ in[43]); 
    assign layer_0[2307] = in[110] | in[112]; 
    assign layer_0[2308] = in[92]; 
    assign layer_0[2309] = in[77] & ~in[3]; 
    assign layer_0[2310] = in[75] | in[94]; 
    assign layer_0[2311] = in[18]; 
    assign layer_0[2312] = ~(in[112] & in[48]); 
    assign layer_0[2313] = ~in[136] | (in[136] & in[101]); 
    assign layer_0[2314] = ~in[214] | (in[214] & in[94]); 
    assign layer_0[2315] = ~in[147]; 
    assign layer_0[2316] = ~(in[46] | in[41]); 
    assign layer_0[2317] = in[216] & ~in[237]; 
    assign layer_0[2318] = ~(in[172] ^ in[45]); 
    assign layer_0[2319] = in[56]; 
    assign layer_0[2320] = ~(in[211] | in[178]); 
    assign layer_0[2321] = in[167] | in[48]; 
    assign layer_0[2322] = ~(in[170] ^ in[157]); 
    assign layer_0[2323] = in[87] | in[131]; 
    assign layer_0[2324] = ~(in[2] | in[61]); 
    assign layer_0[2325] = in[204] & in[182]; 
    assign layer_0[2326] = in[218]; 
    assign layer_0[2327] = in[20]; 
    assign layer_0[2328] = ~(in[44] & in[146]); 
    assign layer_0[2329] = ~in[150] | (in[22] & in[150]); 
    assign layer_0[2330] = ~(in[251] | in[234]); 
    assign layer_0[2331] = in[108] & ~in[193]; 
    assign layer_0[2332] = in[121] & ~in[228]; 
    assign layer_0[2333] = in[126]; 
    assign layer_0[2334] = in[149]; 
    assign layer_0[2335] = ~in[22]; 
    assign layer_0[2336] = ~(in[107] | in[47]); 
    assign layer_0[2337] = ~in[149] | (in[149] & in[82]); 
    assign layer_0[2338] = ~in[55] | (in[55] & in[96]); 
    assign layer_0[2339] = ~in[168] | (in[168] & in[228]); 
    assign layer_0[2340] = in[47] ^ in[126]; 
    assign layer_0[2341] = ~in[131]; 
    assign layer_0[2342] = ~in[105]; 
    assign layer_0[2343] = in[78] & ~in[36]; 
    assign layer_0[2344] = in[107]; 
    assign layer_0[2345] = in[73]; 
    assign layer_0[2346] = ~(in[213] ^ in[96]); 
    assign layer_0[2347] = ~in[128]; 
    assign layer_0[2348] = in[81] ^ in[140]; 
    assign layer_0[2349] = in[90] & ~in[124]; 
    assign layer_0[2350] = ~in[55]; 
    assign layer_0[2351] = in[108] | in[145]; 
    assign layer_0[2352] = ~in[94]; 
    assign layer_0[2353] = ~in[194] | (in[194] & in[240]); 
    assign layer_0[2354] = ~(in[171] | in[45]); 
    assign layer_0[2355] = ~in[195] | (in[195] & in[235]); 
    assign layer_0[2356] = in[19]; 
    assign layer_0[2357] = in[101] ^ in[98]; 
    assign layer_0[2358] = in[208] & in[238]; 
    assign layer_0[2359] = ~in[157]; 
    assign layer_0[2360] = ~in[38] | (in[69] & in[38]); 
    assign layer_0[2361] = in[223] | in[147]; 
    assign layer_0[2362] = ~in[212] | (in[212] & in[255]); 
    assign layer_0[2363] = in[136] & ~in[246]; 
    assign layer_0[2364] = in[86] | in[47]; 
    assign layer_0[2365] = ~(in[74] | in[163]); 
    assign layer_0[2366] = ~in[213]; 
    assign layer_0[2367] = in[41] & ~in[71]; 
    assign layer_0[2368] = in[214]; 
    assign layer_0[2369] = in[163] ^ in[185]; 
    assign layer_0[2370] = ~(in[7] ^ in[102]); 
    assign layer_0[2371] = in[27] | in[138]; 
    assign layer_0[2372] = ~in[99] | (in[206] & in[99]); 
    assign layer_0[2373] = in[244] & ~in[128]; 
    assign layer_0[2374] = ~in[157]; 
    assign layer_0[2375] = in[42]; 
    assign layer_0[2376] = ~in[248] | (in[146] & in[248]); 
    assign layer_0[2377] = ~in[141]; 
    assign layer_0[2378] = in[27] ^ in[129]; 
    assign layer_0[2379] = ~in[74]; 
    assign layer_0[2380] = in[44] | in[66]; 
    assign layer_0[2381] = in[151] & ~in[48]; 
    assign layer_0[2382] = ~in[168] | (in[73] & in[168]); 
    assign layer_0[2383] = in[211] & in[207]; 
    assign layer_0[2384] = in[81] & ~in[74]; 
    assign layer_0[2385] = in[89]; 
    assign layer_0[2386] = ~in[180]; 
    assign layer_0[2387] = in[27] ^ in[30]; 
    assign layer_0[2388] = in[172] ^ in[239]; 
    assign layer_0[2389] = ~(in[117] & in[202]); 
    assign layer_0[2390] = in[102] & ~in[222]; 
    assign layer_0[2391] = ~in[70]; 
    assign layer_0[2392] = in[23] ^ in[49]; 
    assign layer_0[2393] = in[232] ^ in[188]; 
    assign layer_0[2394] = ~in[77]; 
    assign layer_0[2395] = in[131] & ~in[47]; 
    assign layer_0[2396] = ~in[143]; 
    assign layer_0[2397] = in[196]; 
    assign layer_0[2398] = in[231] & ~in[217]; 
    assign layer_0[2399] = ~in[243]; 
    assign layer_0[2400] = in[159] & in[142]; 
    assign layer_0[2401] = ~(in[234] | in[165]); 
    assign layer_0[2402] = in[200] & in[108]; 
    assign layer_0[2403] = ~(in[131] | in[214]); 
    assign layer_0[2404] = ~(in[98] | in[62]); 
    assign layer_0[2405] = in[81]; 
    assign layer_0[2406] = in[2] & ~in[90]; 
    assign layer_0[2407] = ~in[179]; 
    assign layer_0[2408] = in[44] ^ in[76]; 
    assign layer_0[2409] = ~in[228]; 
    assign layer_0[2410] = in[28] & in[129]; 
    assign layer_0[2411] = ~(in[179] | in[187]); 
    assign layer_0[2412] = in[233]; 
    assign layer_0[2413] = 1'b0; 
    assign layer_0[2414] = ~in[125]; 
    assign layer_0[2415] = ~in[168] | (in[164] & in[168]); 
    assign layer_0[2416] = ~in[32] | (in[32] & in[131]); 
    assign layer_0[2417] = ~in[119] | (in[237] & in[119]); 
    assign layer_0[2418] = ~in[73]; 
    assign layer_0[2419] = ~in[109]; 
    assign layer_0[2420] = in[242] & in[227]; 
    assign layer_0[2421] = ~in[212] | (in[185] & in[212]); 
    assign layer_0[2422] = in[126] | in[69]; 
    assign layer_0[2423] = in[238] & in[145]; 
    assign layer_0[2424] = in[27]; 
    assign layer_0[2425] = in[238] & in[209]; 
    assign layer_0[2426] = ~in[26]; 
    assign layer_0[2427] = ~in[234]; 
    assign layer_0[2428] = ~(in[63] & in[53]); 
    assign layer_0[2429] = in[137] & ~in[158]; 
    assign layer_0[2430] = in[132] ^ in[163]; 
    assign layer_0[2431] = in[150] & ~in[202]; 
    assign layer_0[2432] = in[81] ^ in[110]; 
    assign layer_0[2433] = ~(in[146] | in[62]); 
    assign layer_0[2434] = ~in[122] | (in[122] & in[208]); 
    assign layer_0[2435] = ~in[34] | (in[34] & in[92]); 
    assign layer_0[2436] = ~(in[161] ^ in[58]); 
    assign layer_0[2437] = ~(in[96] ^ in[51]); 
    assign layer_0[2438] = in[155]; 
    assign layer_0[2439] = in[35] | in[52]; 
    assign layer_0[2440] = ~in[171] | (in[171] & in[143]); 
    assign layer_0[2441] = ~in[120] | (in[120] & in[191]); 
    assign layer_0[2442] = ~in[25] | (in[32] & in[25]); 
    assign layer_0[2443] = in[218]; 
    assign layer_0[2444] = ~(in[95] & in[141]); 
    assign layer_0[2445] = in[6]; 
    assign layer_0[2446] = in[111] & ~in[177]; 
    assign layer_0[2447] = in[64] & ~in[60]; 
    assign layer_0[2448] = ~(in[132] | in[224]); 
    assign layer_0[2449] = ~(in[48] | in[173]); 
    assign layer_0[2450] = in[7] | in[18]; 
    assign layer_0[2451] = ~(in[39] ^ in[17]); 
    assign layer_0[2452] = ~(in[16] | in[122]); 
    assign layer_0[2453] = in[228] | in[220]; 
    assign layer_0[2454] = in[99] & ~in[192]; 
    assign layer_0[2455] = in[120] & ~in[37]; 
    assign layer_0[2456] = in[244] & ~in[251]; 
    assign layer_0[2457] = in[195]; 
    assign layer_0[2458] = ~(in[186] | in[80]); 
    assign layer_0[2459] = in[191] ^ in[158]; 
    assign layer_0[2460] = in[135] & ~in[129]; 
    assign layer_0[2461] = ~(in[142] ^ in[14]); 
    assign layer_0[2462] = ~in[197]; 
    assign layer_0[2463] = in[179] | in[95]; 
    assign layer_0[2464] = ~in[239]; 
    assign layer_0[2465] = ~(in[118] ^ in[149]); 
    assign layer_0[2466] = in[228]; 
    assign layer_0[2467] = ~in[198]; 
    assign layer_0[2468] = in[75] & ~in[88]; 
    assign layer_0[2469] = in[161] | in[160]; 
    assign layer_0[2470] = in[136]; 
    assign layer_0[2471] = in[70] & in[90]; 
    assign layer_0[2472] = in[248] & ~in[222]; 
    assign layer_0[2473] = in[215]; 
    assign layer_0[2474] = in[168] & ~in[148]; 
    assign layer_0[2475] = ~in[70] | (in[70] & in[144]); 
    assign layer_0[2476] = ~in[65] | (in[92] & in[65]); 
    assign layer_0[2477] = in[58] | in[98]; 
    assign layer_0[2478] = ~(in[138] | in[80]); 
    assign layer_0[2479] = ~in[202]; 
    assign layer_0[2480] = ~(in[65] | in[110]); 
    assign layer_0[2481] = in[181]; 
    assign layer_0[2482] = in[182] ^ in[159]; 
    assign layer_0[2483] = ~(in[194] | in[147]); 
    assign layer_0[2484] = ~(in[176] & in[134]); 
    assign layer_0[2485] = in[204] & in[104]; 
    assign layer_0[2486] = in[249] | in[138]; 
    assign layer_0[2487] = in[66]; 
    assign layer_0[2488] = ~(in[22] | in[33]); 
    assign layer_0[2489] = ~(in[49] ^ in[117]); 
    assign layer_0[2490] = in[233] & in[182]; 
    assign layer_0[2491] = ~(in[207] ^ in[243]); 
    assign layer_0[2492] = ~in[220]; 
    assign layer_0[2493] = in[56]; 
    assign layer_0[2494] = in[97] & ~in[145]; 
    assign layer_0[2495] = in[234] & ~in[175]; 
    assign layer_0[2496] = ~(in[34] ^ in[84]); 
    assign layer_0[2497] = in[69] | in[51]; 
    assign layer_0[2498] = in[65] & in[98]; 
    assign layer_0[2499] = in[167] & ~in[246]; 
    assign layer_0[2500] = in[89] & ~in[13]; 
    assign layer_0[2501] = ~in[215] | (in[226] & in[215]); 
    assign layer_0[2502] = ~(in[76] ^ in[190]); 
    assign layer_0[2503] = in[57]; 
    assign layer_0[2504] = ~(in[53] ^ in[125]); 
    assign layer_0[2505] = in[70]; 
    assign layer_0[2506] = in[153] | in[79]; 
    assign layer_0[2507] = ~(in[232] ^ in[240]); 
    assign layer_0[2508] = ~in[203]; 
    assign layer_0[2509] = in[105] | in[0]; 
    assign layer_0[2510] = in[120] & ~in[114]; 
    assign layer_0[2511] = ~(in[70] ^ in[102]); 
    assign layer_0[2512] = in[83]; 
    assign layer_0[2513] = ~(in[108] ^ in[64]); 
    assign layer_0[2514] = ~in[168] | (in[203] & in[168]); 
    assign layer_0[2515] = in[184]; 
    assign layer_0[2516] = in[80] | in[187]; 
    assign layer_0[2517] = in[114] | in[63]; 
    assign layer_0[2518] = in[65] & ~in[57]; 
    assign layer_0[2519] = ~(in[78] | in[77]); 
    assign layer_0[2520] = in[86]; 
    assign layer_0[2521] = in[69] ^ in[21]; 
    assign layer_0[2522] = in[98] ^ in[85]; 
    assign layer_0[2523] = ~(in[27] | in[2]); 
    assign layer_0[2524] = in[218] & ~in[157]; 
    assign layer_0[2525] = ~in[216]; 
    assign layer_0[2526] = ~in[213] | (in[229] & in[213]); 
    assign layer_0[2527] = in[11] ^ in[3]; 
    assign layer_0[2528] = ~(in[55] | in[47]); 
    assign layer_0[2529] = ~in[127] | (in[127] & in[185]); 
    assign layer_0[2530] = ~(in[157] ^ in[30]); 
    assign layer_0[2531] = ~in[57]; 
    assign layer_0[2532] = ~(in[203] | in[200]); 
    assign layer_0[2533] = ~in[146]; 
    assign layer_0[2534] = ~(in[74] & in[186]); 
    assign layer_0[2535] = ~in[202]; 
    assign layer_0[2536] = ~in[88]; 
    assign layer_0[2537] = in[104]; 
    assign layer_0[2538] = ~in[229] | (in[222] & in[229]); 
    assign layer_0[2539] = in[94] & ~in[1]; 
    assign layer_0[2540] = ~in[65] | (in[192] & in[65]); 
    assign layer_0[2541] = in[190] | in[146]; 
    assign layer_0[2542] = in[99] & ~in[75]; 
    assign layer_0[2543] = ~(in[85] ^ in[80]); 
    assign layer_0[2544] = in[78] & ~in[129]; 
    assign layer_0[2545] = ~in[115]; 
    assign layer_0[2546] = ~(in[80] ^ in[70]); 
    assign layer_0[2547] = in[14] | in[141]; 
    assign layer_0[2548] = in[153] & ~in[190]; 
    assign layer_0[2549] = in[196]; 
    assign layer_0[2550] = in[175] | in[233]; 
    assign layer_0[2551] = in[73] & ~in[80]; 
    assign layer_0[2552] = in[6] | in[46]; 
    assign layer_0[2553] = ~(in[55] | in[177]); 
    assign layer_0[2554] = ~(in[244] ^ in[202]); 
    assign layer_0[2555] = in[35] & ~in[69]; 
    assign layer_0[2556] = ~(in[105] | in[181]); 
    assign layer_0[2557] = ~in[9] | (in[55] & in[9]); 
    assign layer_0[2558] = ~in[40] | (in[40] & in[33]); 
    assign layer_0[2559] = ~in[78] | (in[12] & in[78]); 
    assign layer_0[2560] = ~(in[224] | in[198]); 
    assign layer_0[2561] = in[65]; 
    assign layer_0[2562] = ~(in[144] & in[104]); 
    assign layer_0[2563] = ~(in[221] | in[195]); 
    assign layer_0[2564] = in[79] & ~in[77]; 
    assign layer_0[2565] = ~(in[64] ^ in[179]); 
    assign layer_0[2566] = ~in[166]; 
    assign layer_0[2567] = in[46] ^ in[48]; 
    assign layer_0[2568] = in[121]; 
    assign layer_0[2569] = in[242]; 
    assign layer_0[2570] = in[89]; 
    assign layer_0[2571] = in[129] ^ in[33]; 
    assign layer_0[2572] = in[66] ^ in[1]; 
    assign layer_0[2573] = ~in[168] | (in[124] & in[168]); 
    assign layer_0[2574] = in[66] | in[44]; 
    assign layer_0[2575] = ~in[99] | (in[99] & in[175]); 
    assign layer_0[2576] = in[184]; 
    assign layer_0[2577] = in[62] & ~in[186]; 
    assign layer_0[2578] = ~(in[110] | in[117]); 
    assign layer_0[2579] = in[95] & in[99]; 
    assign layer_0[2580] = in[73]; 
    assign layer_0[2581] = in[80] ^ in[162]; 
    assign layer_0[2582] = ~(in[216] | in[130]); 
    assign layer_0[2583] = in[31]; 
    assign layer_0[2584] = ~in[198]; 
    assign layer_0[2585] = ~(in[211] ^ in[99]); 
    assign layer_0[2586] = in[184]; 
    assign layer_0[2587] = ~in[121]; 
    assign layer_0[2588] = ~in[70] | (in[17] & in[70]); 
    assign layer_0[2589] = in[216] ^ in[234]; 
    assign layer_0[2590] = ~in[200] | (in[200] & in[236]); 
    assign layer_0[2591] = ~in[64]; 
    assign layer_0[2592] = ~in[119] | (in[56] & in[119]); 
    assign layer_0[2593] = ~in[141]; 
    assign layer_0[2594] = in[251] & ~in[235]; 
    assign layer_0[2595] = in[107] & in[166]; 
    assign layer_0[2596] = ~in[104] | (in[104] & in[210]); 
    assign layer_0[2597] = ~in[56]; 
    assign layer_0[2598] = ~in[88] | (in[95] & in[88]); 
    assign layer_0[2599] = ~(in[240] & in[123]); 
    assign layer_0[2600] = in[106] & ~in[182]; 
    assign layer_0[2601] = ~in[102]; 
    assign layer_0[2602] = in[9] & in[23]; 
    assign layer_0[2603] = ~in[111]; 
    assign layer_0[2604] = ~in[149] | (in[149] & in[94]); 
    assign layer_0[2605] = ~in[134] | (in[134] & in[132]); 
    assign layer_0[2606] = ~in[166] | (in[54] & in[166]); 
    assign layer_0[2607] = ~(in[20] | in[123]); 
    assign layer_0[2608] = ~in[88] | (in[88] & in[9]); 
    assign layer_0[2609] = ~(in[55] ^ in[104]); 
    assign layer_0[2610] = in[254]; 
    assign layer_0[2611] = ~in[93] | (in[12] & in[93]); 
    assign layer_0[2612] = ~in[225] | (in[164] & in[225]); 
    assign layer_0[2613] = in[98]; 
    assign layer_0[2614] = ~(in[196] | in[68]); 
    assign layer_0[2615] = in[149]; 
    assign layer_0[2616] = in[33] | in[85]; 
    assign layer_0[2617] = ~in[4] | (in[4] & in[98]); 
    assign layer_0[2618] = ~in[165] | (in[47] & in[165]); 
    assign layer_0[2619] = in[87] | in[94]; 
    assign layer_0[2620] = ~(in[252] | in[222]); 
    assign layer_0[2621] = ~in[7] | (in[7] & in[128]); 
    assign layer_0[2622] = ~(in[28] | in[26]); 
    assign layer_0[2623] = in[173] ^ in[47]; 
    assign layer_0[2624] = ~(in[72] | in[63]); 
    assign layer_0[2625] = in[166]; 
    assign layer_0[2626] = in[0] | in[21]; 
    assign layer_0[2627] = in[63] & ~in[36]; 
    assign layer_0[2628] = in[83] & ~in[142]; 
    assign layer_0[2629] = in[26] | in[141]; 
    assign layer_0[2630] = ~in[154] | (in[154] & in[142]); 
    assign layer_0[2631] = ~(in[0] & in[10]); 
    assign layer_0[2632] = in[238] & ~in[163]; 
    assign layer_0[2633] = ~in[74] | (in[33] & in[74]); 
    assign layer_0[2634] = in[214]; 
    assign layer_0[2635] = in[132] & ~in[90]; 
    assign layer_0[2636] = ~in[204]; 
    assign layer_0[2637] = in[95] | in[2]; 
    assign layer_0[2638] = in[27] & ~in[71]; 
    assign layer_0[2639] = in[57] ^ in[177]; 
    assign layer_0[2640] = in[213] | in[176]; 
    assign layer_0[2641] = in[127] & in[16]; 
    assign layer_0[2642] = in[49]; 
    assign layer_0[2643] = in[198] | in[86]; 
    assign layer_0[2644] = ~(in[102] | in[31]); 
    assign layer_0[2645] = in[217]; 
    assign layer_0[2646] = ~(in[12] | in[24]); 
    assign layer_0[2647] = ~in[152] | (in[160] & in[152]); 
    assign layer_0[2648] = in[191] & ~in[80]; 
    assign layer_0[2649] = in[251] ^ in[168]; 
    assign layer_0[2650] = in[56] & in[120]; 
    assign layer_0[2651] = ~in[233]; 
    assign layer_0[2652] = ~(in[4] | in[87]); 
    assign layer_0[2653] = ~in[168] | (in[238] & in[168]); 
    assign layer_0[2654] = ~(in[205] ^ in[224]); 
    assign layer_0[2655] = ~(in[41] ^ in[0]); 
    assign layer_0[2656] = in[218]; 
    assign layer_0[2657] = in[211]; 
    assign layer_0[2658] = in[226]; 
    assign layer_0[2659] = ~(in[158] ^ in[157]); 
    assign layer_0[2660] = ~(in[15] | in[109]); 
    assign layer_0[2661] = in[11] & ~in[6]; 
    assign layer_0[2662] = ~in[19]; 
    assign layer_0[2663] = ~(in[158] ^ in[68]); 
    assign layer_0[2664] = in[181]; 
    assign layer_0[2665] = ~in[222]; 
    assign layer_0[2666] = ~in[156]; 
    assign layer_0[2667] = ~in[178]; 
    assign layer_0[2668] = in[61] | in[35]; 
    assign layer_0[2669] = in[35] & ~in[39]; 
    assign layer_0[2670] = in[124] | in[123]; 
    assign layer_0[2671] = ~(in[49] | in[147]); 
    assign layer_0[2672] = ~in[133] | (in[133] & in[82]); 
    assign layer_0[2673] = in[237] | in[247]; 
    assign layer_0[2674] = ~in[65]; 
    assign layer_0[2675] = ~in[244] | (in[255] & in[244]); 
    assign layer_0[2676] = in[132] ^ in[110]; 
    assign layer_0[2677] = in[190] | in[99]; 
    assign layer_0[2678] = ~(in[96] | in[74]); 
    assign layer_0[2679] = ~(in[222] & in[176]); 
    assign layer_0[2680] = in[242] & ~in[169]; 
    assign layer_0[2681] = in[213] & in[131]; 
    assign layer_0[2682] = in[176] ^ in[240]; 
    assign layer_0[2683] = in[5]; 
    assign layer_0[2684] = ~(in[110] | in[111]); 
    assign layer_0[2685] = in[84] ^ in[30]; 
    assign layer_0[2686] = in[144]; 
    assign layer_0[2687] = in[192] & in[159]; 
    assign layer_0[2688] = in[84] & ~in[34]; 
    assign layer_0[2689] = in[174]; 
    assign layer_0[2690] = ~in[126]; 
    assign layer_0[2691] = ~(in[75] | in[38]); 
    assign layer_0[2692] = in[197] & in[164]; 
    assign layer_0[2693] = ~in[223]; 
    assign layer_0[2694] = ~(in[201] ^ in[234]); 
    assign layer_0[2695] = ~in[213]; 
    assign layer_0[2696] = ~(in[200] | in[202]); 
    assign layer_0[2697] = in[62]; 
    assign layer_0[2698] = ~in[117]; 
    assign layer_0[2699] = in[35] | in[163]; 
    assign layer_0[2700] = ~(in[171] ^ in[209]); 
    assign layer_0[2701] = in[113] | in[215]; 
    assign layer_0[2702] = in[19] | in[6]; 
    assign layer_0[2703] = in[39] & ~in[152]; 
    assign layer_0[2704] = ~(in[82] ^ in[22]); 
    assign layer_0[2705] = ~in[122] | (in[122] & in[181]); 
    assign layer_0[2706] = ~(in[105] | in[128]); 
    assign layer_0[2707] = ~(in[55] & in[14]); 
    assign layer_0[2708] = ~in[198]; 
    assign layer_0[2709] = in[43] & ~in[171]; 
    assign layer_0[2710] = in[0]; 
    assign layer_0[2711] = in[251] | in[253]; 
    assign layer_0[2712] = ~(in[117] | in[21]); 
    assign layer_0[2713] = ~(in[0] | in[8]); 
    assign layer_0[2714] = in[159]; 
    assign layer_0[2715] = in[173]; 
    assign layer_0[2716] = ~in[45]; 
    assign layer_0[2717] = ~(in[181] ^ in[95]); 
    assign layer_0[2718] = ~(in[5] & in[125]); 
    assign layer_0[2719] = ~in[150] | (in[56] & in[150]); 
    assign layer_0[2720] = ~(in[241] & in[199]); 
    assign layer_0[2721] = in[108] & ~in[49]; 
    assign layer_0[2722] = in[156]; 
    assign layer_0[2723] = in[67] | in[159]; 
    assign layer_0[2724] = in[57]; 
    assign layer_0[2725] = ~(in[172] | in[119]); 
    assign layer_0[2726] = ~in[167]; 
    assign layer_0[2727] = ~(in[161] | in[255]); 
    assign layer_0[2728] = in[152] & in[196]; 
    assign layer_0[2729] = ~in[240]; 
    assign layer_0[2730] = ~(in[133] | in[141]); 
    assign layer_0[2731] = in[168]; 
    assign layer_0[2732] = ~(in[144] & in[47]); 
    assign layer_0[2733] = in[102] & in[201]; 
    assign layer_0[2734] = in[217]; 
    assign layer_0[2735] = ~(in[238] ^ in[239]); 
    assign layer_0[2736] = ~(in[82] | in[121]); 
    assign layer_0[2737] = ~in[135] | (in[117] & in[135]); 
    assign layer_0[2738] = in[182] | in[161]; 
    assign layer_0[2739] = in[114]; 
    assign layer_0[2740] = in[161] & ~in[181]; 
    assign layer_0[2741] = ~(in[195] | in[75]); 
    assign layer_0[2742] = in[244]; 
    assign layer_0[2743] = in[131] & ~in[21]; 
    assign layer_0[2744] = ~in[119] | (in[239] & in[119]); 
    assign layer_0[2745] = ~in[31] | (in[31] & in[143]); 
    assign layer_0[2746] = in[103] & ~in[200]; 
    assign layer_0[2747] = in[142] & ~in[211]; 
    assign layer_0[2748] = in[88] & ~in[182]; 
    assign layer_0[2749] = ~in[102] | (in[64] & in[102]); 
    assign layer_0[2750] = ~(in[60] | in[84]); 
    assign layer_0[2751] = ~(in[62] | in[41]); 
    assign layer_0[2752] = ~(in[247] | in[248]); 
    assign layer_0[2753] = in[213] & ~in[222]; 
    assign layer_0[2754] = ~in[230]; 
    assign layer_0[2755] = in[225] & in[246]; 
    assign layer_0[2756] = ~in[26]; 
    assign layer_0[2757] = in[223] & in[112]; 
    assign layer_0[2758] = ~in[215] | (in[215] & in[159]); 
    assign layer_0[2759] = in[31] & in[56]; 
    assign layer_0[2760] = in[184] | in[112]; 
    assign layer_0[2761] = ~in[247] | (in[247] & in[159]); 
    assign layer_0[2762] = ~(in[209] ^ in[123]); 
    assign layer_0[2763] = in[24]; 
    assign layer_0[2764] = in[168] & ~in[83]; 
    assign layer_0[2765] = ~in[89] | (in[53] & in[89]); 
    assign layer_0[2766] = in[219]; 
    assign layer_0[2767] = ~(in[134] & in[162]); 
    assign layer_0[2768] = ~in[226] | (in[226] & in[138]); 
    assign layer_0[2769] = ~in[167]; 
    assign layer_0[2770] = in[88]; 
    assign layer_0[2771] = ~in[140] | (in[83] & in[140]); 
    assign layer_0[2772] = ~in[206]; 
    assign layer_0[2773] = ~in[148] | (in[148] & in[60]); 
    assign layer_0[2774] = in[163] ^ in[52]; 
    assign layer_0[2775] = ~in[239] | (in[239] & in[111]); 
    assign layer_0[2776] = ~(in[8] ^ in[95]); 
    assign layer_0[2777] = ~in[195]; 
    assign layer_0[2778] = ~in[89]; 
    assign layer_0[2779] = in[71]; 
    assign layer_0[2780] = in[11]; 
    assign layer_0[2781] = ~(in[156] ^ in[98]); 
    assign layer_0[2782] = ~in[75]; 
    assign layer_0[2783] = in[110] | in[177]; 
    assign layer_0[2784] = ~in[29]; 
    assign layer_0[2785] = ~(in[164] ^ in[205]); 
    assign layer_0[2786] = ~(in[219] & in[218]); 
    assign layer_0[2787] = in[170] & ~in[156]; 
    assign layer_0[2788] = ~(in[94] | in[217]); 
    assign layer_0[2789] = ~in[168] | (in[168] & in[176]); 
    assign layer_0[2790] = ~in[0] | (in[34] & in[0]); 
    assign layer_0[2791] = ~(in[233] ^ in[169]); 
    assign layer_0[2792] = ~(in[111] | in[230]); 
    assign layer_0[2793] = ~(in[230] | in[242]); 
    assign layer_0[2794] = in[12] & in[116]; 
    assign layer_0[2795] = in[87] ^ in[84]; 
    assign layer_0[2796] = ~(in[136] & in[134]); 
    assign layer_0[2797] = in[71] & ~in[124]; 
    assign layer_0[2798] = ~in[49]; 
    assign layer_0[2799] = ~in[58] | (in[23] & in[58]); 
    assign layer_0[2800] = in[104]; 
    assign layer_0[2801] = ~in[123]; 
    assign layer_0[2802] = ~in[20]; 
    assign layer_0[2803] = in[165]; 
    assign layer_0[2804] = ~(in[56] ^ in[168]); 
    assign layer_0[2805] = ~in[20] | (in[20] & in[111]); 
    assign layer_0[2806] = in[110] | in[79]; 
    assign layer_0[2807] = in[224] & in[197]; 
    assign layer_0[2808] = ~(in[132] | in[245]); 
    assign layer_0[2809] = in[102] & ~in[134]; 
    assign layer_0[2810] = ~in[73] | (in[73] & in[35]); 
    assign layer_0[2811] = ~(in[244] | in[161]); 
    assign layer_0[2812] = ~(in[40] & in[3]); 
    assign layer_0[2813] = in[144]; 
    assign layer_0[2814] = ~(in[78] | in[132]); 
    assign layer_0[2815] = ~in[68] | (in[159] & in[68]); 
    assign layer_0[2816] = in[185] & ~in[206]; 
    assign layer_0[2817] = ~(in[222] & in[233]); 
    assign layer_0[2818] = in[55] ^ in[91]; 
    assign layer_0[2819] = in[246]; 
    assign layer_0[2820] = in[110]; 
    assign layer_0[2821] = in[46] ^ in[2]; 
    assign layer_0[2822] = in[82]; 
    assign layer_0[2823] = ~in[109]; 
    assign layer_0[2824] = in[3] & ~in[81]; 
    assign layer_0[2825] = ~in[163]; 
    assign layer_0[2826] = ~in[49] | (in[19] & in[49]); 
    assign layer_0[2827] = in[190]; 
    assign layer_0[2828] = ~in[80] | (in[80] & in[11]); 
    assign layer_0[2829] = ~(in[66] | in[38]); 
    assign layer_0[2830] = in[71] & ~in[66]; 
    assign layer_0[2831] = ~in[246]; 
    assign layer_0[2832] = in[38]; 
    assign layer_0[2833] = ~in[148] | (in[64] & in[148]); 
    assign layer_0[2834] = in[151]; 
    assign layer_0[2835] = in[213] & ~in[95]; 
    assign layer_0[2836] = in[183]; 
    assign layer_0[2837] = ~(in[33] & in[37]); 
    assign layer_0[2838] = in[162] & ~in[133]; 
    assign layer_0[2839] = in[72]; 
    assign layer_0[2840] = ~(in[163] ^ in[222]); 
    assign layer_0[2841] = ~in[208]; 
    assign layer_0[2842] = in[133] & ~in[21]; 
    assign layer_0[2843] = ~(in[36] ^ in[83]); 
    assign layer_0[2844] = in[74]; 
    assign layer_0[2845] = in[169]; 
    assign layer_0[2846] = ~in[92] | (in[92] & in[28]); 
    assign layer_0[2847] = ~in[156]; 
    assign layer_0[2848] = in[157]; 
    assign layer_0[2849] = ~(in[90] & in[204]); 
    assign layer_0[2850] = in[42] & ~in[32]; 
    assign layer_0[2851] = in[231] | in[229]; 
    assign layer_0[2852] = ~in[71] | (in[71] & in[186]); 
    assign layer_0[2853] = in[218]; 
    assign layer_0[2854] = in[215] & ~in[147]; 
    assign layer_0[2855] = in[90]; 
    assign layer_0[2856] = ~(in[182] ^ in[118]); 
    assign layer_0[2857] = in[125]; 
    assign layer_0[2858] = ~in[123]; 
    assign layer_0[2859] = ~(in[226] & in[230]); 
    assign layer_0[2860] = ~(in[66] ^ in[84]); 
    assign layer_0[2861] = ~in[238] | (in[114] & in[238]); 
    assign layer_0[2862] = in[90] & ~in[15]; 
    assign layer_0[2863] = in[250]; 
    assign layer_0[2864] = in[105]; 
    assign layer_0[2865] = ~(in[239] | in[151]); 
    assign layer_0[2866] = in[89] & ~in[132]; 
    assign layer_0[2867] = in[93] ^ in[83]; 
    assign layer_0[2868] = ~in[143]; 
    assign layer_0[2869] = ~(in[113] | in[180]); 
    assign layer_0[2870] = in[164] & in[180]; 
    assign layer_0[2871] = ~(in[188] ^ in[220]); 
    assign layer_0[2872] = ~in[70]; 
    assign layer_0[2873] = in[157]; 
    assign layer_0[2874] = ~(in[228] ^ in[251]); 
    assign layer_0[2875] = ~in[168] | (in[168] & in[170]); 
    assign layer_0[2876] = ~in[13] | (in[13] & in[80]); 
    assign layer_0[2877] = ~(in[1] ^ in[102]); 
    assign layer_0[2878] = ~in[197]; 
    assign layer_0[2879] = in[193] | in[72]; 
    assign layer_0[2880] = ~in[105]; 
    assign layer_0[2881] = ~in[113] | (in[18] & in[113]); 
    assign layer_0[2882] = in[90] & in[106]; 
    assign layer_0[2883] = ~in[61]; 
    assign layer_0[2884] = in[85] & ~in[66]; 
    assign layer_0[2885] = ~in[244] | (in[244] & in[129]); 
    assign layer_0[2886] = ~in[1] | (in[1] & in[87]); 
    assign layer_0[2887] = in[247]; 
    assign layer_0[2888] = in[64] | in[53]; 
    assign layer_0[2889] = ~in[228] | (in[228] & in[222]); 
    assign layer_0[2890] = in[90] ^ in[91]; 
    assign layer_0[2891] = in[243] ^ in[127]; 
    assign layer_0[2892] = ~in[45] | (in[109] & in[45]); 
    assign layer_0[2893] = ~(in[164] ^ in[212]); 
    assign layer_0[2894] = ~in[165] | (in[244] & in[165]); 
    assign layer_0[2895] = ~in[29] | (in[29] & in[30]); 
    assign layer_0[2896] = in[200] | in[255]; 
    assign layer_0[2897] = ~in[178] | (in[244] & in[178]); 
    assign layer_0[2898] = in[76] & ~in[144]; 
    assign layer_0[2899] = in[126]; 
    assign layer_0[2900] = ~(in[143] ^ in[224]); 
    assign layer_0[2901] = in[0] & ~in[106]; 
    assign layer_0[2902] = in[9] ^ in[22]; 
    assign layer_0[2903] = in[117]; 
    assign layer_0[2904] = in[248]; 
    assign layer_0[2905] = in[162]; 
    assign layer_0[2906] = in[198] & ~in[224]; 
    assign layer_0[2907] = ~(in[225] & in[176]); 
    assign layer_0[2908] = in[116] | in[124]; 
    assign layer_0[2909] = in[252] & ~in[185]; 
    assign layer_0[2910] = in[91] & ~in[65]; 
    assign layer_0[2911] = ~in[201]; 
    assign layer_0[2912] = ~(in[203] | in[212]); 
    assign layer_0[2913] = ~in[152] | (in[152] & in[40]); 
    assign layer_0[2914] = ~(in[241] ^ in[136]); 
    assign layer_0[2915] = in[15] & ~in[142]; 
    assign layer_0[2916] = in[104] & ~in[219]; 
    assign layer_0[2917] = ~(in[169] ^ in[110]); 
    assign layer_0[2918] = in[139] & ~in[38]; 
    assign layer_0[2919] = in[53] & ~in[111]; 
    assign layer_0[2920] = in[199] | in[213]; 
    assign layer_0[2921] = in[164]; 
    assign layer_0[2922] = in[126]; 
    assign layer_0[2923] = in[107]; 
    assign layer_0[2924] = in[251] | in[233]; 
    assign layer_0[2925] = in[149]; 
    assign layer_0[2926] = in[235] & ~in[125]; 
    assign layer_0[2927] = in[150]; 
    assign layer_0[2928] = ~(in[44] & in[147]); 
    assign layer_0[2929] = in[246] & ~in[143]; 
    assign layer_0[2930] = in[119]; 
    assign layer_0[2931] = ~(in[83] ^ in[147]); 
    assign layer_0[2932] = ~in[78] | (in[77] & in[78]); 
    assign layer_0[2933] = ~(in[208] | in[167]); 
    assign layer_0[2934] = in[173] & ~in[232]; 
    assign layer_0[2935] = in[39]; 
    assign layer_0[2936] = in[19]; 
    assign layer_0[2937] = ~(in[145] | in[25]); 
    assign layer_0[2938] = in[149] & ~in[247]; 
    assign layer_0[2939] = in[36] ^ in[60]; 
    assign layer_0[2940] = ~(in[109] | in[51]); 
    assign layer_0[2941] = in[52] ^ in[134]; 
    assign layer_0[2942] = ~in[87] | (in[87] & in[29]); 
    assign layer_0[2943] = in[204]; 
    assign layer_0[2944] = in[252] ^ in[193]; 
    assign layer_0[2945] = in[48] & in[129]; 
    assign layer_0[2946] = in[133] ^ in[230]; 
    assign layer_0[2947] = in[82]; 
    assign layer_0[2948] = in[88]; 
    assign layer_0[2949] = ~in[237]; 
    assign layer_0[2950] = ~(in[57] & in[173]); 
    assign layer_0[2951] = in[82]; 
    assign layer_0[2952] = ~in[22] | (in[37] & in[22]); 
    assign layer_0[2953] = in[124] ^ in[84]; 
    assign layer_0[2954] = in[27]; 
    assign layer_0[2955] = ~(in[43] ^ in[14]); 
    assign layer_0[2956] = in[118]; 
    assign layer_0[2957] = ~in[182] | (in[157] & in[182]); 
    assign layer_0[2958] = ~in[45]; 
    assign layer_0[2959] = in[181]; 
    assign layer_0[2960] = ~in[146]; 
    assign layer_0[2961] = in[184] & ~in[183]; 
    assign layer_0[2962] = in[165]; 
    assign layer_0[2963] = ~(in[97] ^ in[150]); 
    assign layer_0[2964] = ~(in[95] ^ in[201]); 
    assign layer_0[2965] = in[19]; 
    assign layer_0[2966] = ~in[95]; 
    assign layer_0[2967] = in[241] | in[124]; 
    assign layer_0[2968] = in[107]; 
    assign layer_0[2969] = ~(in[50] | in[101]); 
    assign layer_0[2970] = ~in[163] | (in[93] & in[163]); 
    assign layer_0[2971] = in[154]; 
    assign layer_0[2972] = in[86]; 
    assign layer_0[2973] = ~in[72] | (in[72] & in[137]); 
    assign layer_0[2974] = ~in[181]; 
    assign layer_0[2975] = ~in[196] | (in[236] & in[196]); 
    assign layer_0[2976] = in[131]; 
    assign layer_0[2977] = in[207] & ~in[179]; 
    assign layer_0[2978] = in[100] ^ in[147]; 
    assign layer_0[2979] = ~(in[83] & in[13]); 
    assign layer_0[2980] = in[51] | in[34]; 
    assign layer_0[2981] = ~in[58]; 
    assign layer_0[2982] = in[199] | in[225]; 
    assign layer_0[2983] = ~in[106]; 
    assign layer_0[2984] = ~in[72] | (in[72] & in[192]); 
    assign layer_0[2985] = in[221] ^ in[172]; 
    assign layer_0[2986] = ~in[77]; 
    assign layer_0[2987] = in[131] ^ in[197]; 
    assign layer_0[2988] = ~in[24] | (in[24] & in[93]); 
    assign layer_0[2989] = ~in[82]; 
    assign layer_0[2990] = ~in[202] | (in[159] & in[202]); 
    assign layer_0[2991] = ~(in[253] ^ in[209]); 
    assign layer_0[2992] = ~(in[11] & in[115]); 
    assign layer_0[2993] = ~(in[34] & in[33]); 
    assign layer_0[2994] = in[41]; 
    assign layer_0[2995] = in[133] & ~in[107]; 
    assign layer_0[2996] = in[132] & ~in[89]; 
    assign layer_0[2997] = in[169] | in[195]; 
    assign layer_0[2998] = ~in[39]; 
    assign layer_0[2999] = ~(in[1] | in[54]); 
    assign layer_0[3000] = in[57]; 
    assign layer_0[3001] = in[157] & ~in[145]; 
    assign layer_0[3002] = in[110]; 
    assign layer_0[3003] = ~(in[54] | in[160]); 
    assign layer_0[3004] = in[159] | in[245]; 
    assign layer_0[3005] = in[20] | in[98]; 
    assign layer_0[3006] = ~in[152]; 
    assign layer_0[3007] = in[60] & ~in[181]; 
    assign layer_0[3008] = in[210] | in[111]; 
    assign layer_0[3009] = ~(in[11] ^ in[40]); 
    assign layer_0[3010] = in[178] | in[85]; 
    assign layer_0[3011] = in[126] ^ in[170]; 
    assign layer_0[3012] = ~in[150]; 
    assign layer_0[3013] = ~(in[40] | in[30]); 
    assign layer_0[3014] = ~(in[245] ^ in[147]); 
    assign layer_0[3015] = ~in[149]; 
    assign layer_0[3016] = in[54] & in[90]; 
    assign layer_0[3017] = ~in[95] | (in[95] & in[145]); 
    assign layer_0[3018] = in[113] ^ in[15]; 
    assign layer_0[3019] = ~in[121] | (in[20] & in[121]); 
    assign layer_0[3020] = in[126]; 
    assign layer_0[3021] = in[112] & ~in[240]; 
    assign layer_0[3022] = in[125] | in[60]; 
    assign layer_0[3023] = in[206] & ~in[228]; 
    assign layer_0[3024] = ~in[177]; 
    assign layer_0[3025] = ~(in[183] ^ in[85]); 
    assign layer_0[3026] = ~(in[223] & in[174]); 
    assign layer_0[3027] = ~in[160] | (in[129] & in[160]); 
    assign layer_0[3028] = in[228] & ~in[157]; 
    assign layer_0[3029] = in[89] & in[199]; 
    assign layer_0[3030] = in[175]; 
    assign layer_0[3031] = ~(in[121] | in[84]); 
    assign layer_0[3032] = ~(in[150] ^ in[112]); 
    assign layer_0[3033] = in[242]; 
    assign layer_0[3034] = in[151] & ~in[229]; 
    assign layer_0[3035] = in[186] | in[125]; 
    assign layer_0[3036] = ~in[157]; 
    assign layer_0[3037] = ~(in[73] & in[122]); 
    assign layer_0[3038] = in[152]; 
    assign layer_0[3039] = ~in[108]; 
    assign layer_0[3040] = in[232] & ~in[171]; 
    assign layer_0[3041] = in[79] | in[176]; 
    assign layer_0[3042] = in[79] & in[115]; 
    assign layer_0[3043] = ~in[166]; 
    assign layer_0[3044] = in[83] & ~in[200]; 
    assign layer_0[3045] = ~(in[63] ^ in[53]); 
    assign layer_0[3046] = in[129] | in[232]; 
    assign layer_0[3047] = ~in[160]; 
    assign layer_0[3048] = ~in[86] | (in[155] & in[86]); 
    assign layer_0[3049] = in[242] & ~in[241]; 
    assign layer_0[3050] = in[178]; 
    assign layer_0[3051] = in[229]; 
    assign layer_0[3052] = in[17] | in[9]; 
    assign layer_0[3053] = in[32] | in[112]; 
    assign layer_0[3054] = ~in[165] | (in[129] & in[165]); 
    assign layer_0[3055] = ~(in[54] & in[180]); 
    assign layer_0[3056] = ~(in[82] | in[179]); 
    assign layer_0[3057] = in[254] & in[129]; 
    assign layer_0[3058] = in[61]; 
    assign layer_0[3059] = ~in[139]; 
    assign layer_0[3060] = ~in[225] | (in[217] & in[225]); 
    assign layer_0[3061] = ~(in[145] ^ in[130]); 
    assign layer_0[3062] = ~(in[158] ^ in[40]); 
    assign layer_0[3063] = ~(in[175] | in[171]); 
    assign layer_0[3064] = in[238] | in[166]; 
    assign layer_0[3065] = in[163]; 
    assign layer_0[3066] = ~(in[157] ^ in[208]); 
    assign layer_0[3067] = in[182] & in[106]; 
    assign layer_0[3068] = in[101]; 
    assign layer_0[3069] = in[34] & in[69]; 
    assign layer_0[3070] = ~in[216] | (in[164] & in[216]); 
    assign layer_0[3071] = ~in[182] | (in[182] & in[235]); 
    assign layer_0[3072] = ~(in[55] ^ in[84]); 
    assign layer_0[3073] = in[132] ^ in[16]; 
    assign layer_0[3074] = in[201] & ~in[85]; 
    assign layer_0[3075] = ~in[128] | (in[128] & in[192]); 
    assign layer_0[3076] = ~(in[100] ^ in[17]); 
    assign layer_0[3077] = ~(in[40] | in[81]); 
    assign layer_0[3078] = in[217] & ~in[208]; 
    assign layer_0[3079] = in[109] ^ in[147]; 
    assign layer_0[3080] = in[164] | in[203]; 
    assign layer_0[3081] = ~(in[139] & in[152]); 
    assign layer_0[3082] = ~(in[126] & in[238]); 
    assign layer_0[3083] = ~(in[101] ^ in[87]); 
    assign layer_0[3084] = in[219] & ~in[229]; 
    assign layer_0[3085] = in[81] & ~in[3]; 
    assign layer_0[3086] = ~(in[242] | in[160]); 
    assign layer_0[3087] = ~in[211] | (in[211] & in[235]); 
    assign layer_0[3088] = ~in[147]; 
    assign layer_0[3089] = ~in[89] | (in[151] & in[89]); 
    assign layer_0[3090] = ~in[232] | (in[144] & in[232]); 
    assign layer_0[3091] = in[213] & ~in[125]; 
    assign layer_0[3092] = ~(in[152] ^ in[247]); 
    assign layer_0[3093] = ~in[106]; 
    assign layer_0[3094] = in[38] & ~in[96]; 
    assign layer_0[3095] = ~in[244] | (in[246] & in[244]); 
    assign layer_0[3096] = ~in[74]; 
    assign layer_0[3097] = ~(in[248] | in[232]); 
    assign layer_0[3098] = in[10] | in[69]; 
    assign layer_0[3099] = ~(in[180] ^ in[121]); 
    assign layer_0[3100] = ~in[90]; 
    assign layer_0[3101] = ~in[140]; 
    assign layer_0[3102] = in[137] & ~in[252]; 
    assign layer_0[3103] = ~(in[140] & in[61]); 
    assign layer_0[3104] = ~(in[14] & in[96]); 
    assign layer_0[3105] = ~in[49]; 
    assign layer_0[3106] = in[54] & ~in[133]; 
    assign layer_0[3107] = in[165]; 
    assign layer_0[3108] = ~in[196]; 
    assign layer_0[3109] = in[79] & ~in[128]; 
    assign layer_0[3110] = in[57] & in[177]; 
    assign layer_0[3111] = ~in[89]; 
    assign layer_0[3112] = in[70]; 
    assign layer_0[3113] = ~in[142]; 
    assign layer_0[3114] = ~(in[180] & in[226]); 
    assign layer_0[3115] = in[192] & in[145]; 
    assign layer_0[3116] = ~in[77]; 
    assign layer_0[3117] = ~in[181]; 
    assign layer_0[3118] = in[254]; 
    assign layer_0[3119] = in[3] | in[89]; 
    assign layer_0[3120] = in[108] | in[174]; 
    assign layer_0[3121] = in[73]; 
    assign layer_0[3122] = in[253] & ~in[168]; 
    assign layer_0[3123] = in[21] | in[53]; 
    assign layer_0[3124] = ~(in[51] ^ in[134]); 
    assign layer_0[3125] = ~in[17] | (in[40] & in[17]); 
    assign layer_0[3126] = ~in[38] | (in[38] & in[64]); 
    assign layer_0[3127] = in[31] & in[157]; 
    assign layer_0[3128] = ~in[134]; 
    assign layer_0[3129] = in[81] | in[46]; 
    assign layer_0[3130] = ~in[46] | (in[7] & in[46]); 
    assign layer_0[3131] = in[60] ^ in[13]; 
    assign layer_0[3132] = in[2] & in[58]; 
    assign layer_0[3133] = ~(in[143] | in[193]); 
    assign layer_0[3134] = in[97] | in[42]; 
    assign layer_0[3135] = in[194]; 
    assign layer_0[3136] = ~(in[30] & in[21]); 
    assign layer_0[3137] = ~in[243]; 
    assign layer_0[3138] = ~(in[248] | in[183]); 
    assign layer_0[3139] = in[92]; 
    assign layer_0[3140] = in[165]; 
    assign layer_0[3141] = in[190] ^ in[98]; 
    assign layer_0[3142] = in[24] | in[60]; 
    assign layer_0[3143] = ~(in[204] ^ in[111]); 
    assign layer_0[3144] = in[172] | in[190]; 
    assign layer_0[3145] = in[198]; 
    assign layer_0[3146] = in[117]; 
    assign layer_0[3147] = in[77]; 
    assign layer_0[3148] = in[30] | in[122]; 
    assign layer_0[3149] = ~in[40] | (in[26] & in[40]); 
    assign layer_0[3150] = ~(in[116] ^ in[176]); 
    assign layer_0[3151] = in[120] | in[74]; 
    assign layer_0[3152] = ~in[227]; 
    assign layer_0[3153] = in[215] & in[90]; 
    assign layer_0[3154] = in[195] | in[163]; 
    assign layer_0[3155] = ~in[249]; 
    assign layer_0[3156] = in[71]; 
    assign layer_0[3157] = in[199] & in[101]; 
    assign layer_0[3158] = in[76]; 
    assign layer_0[3159] = in[149]; 
    assign layer_0[3160] = in[28]; 
    assign layer_0[3161] = ~(in[227] | in[226]); 
    assign layer_0[3162] = ~(in[152] & in[81]); 
    assign layer_0[3163] = in[67] & ~in[100]; 
    assign layer_0[3164] = in[238] ^ in[111]; 
    assign layer_0[3165] = ~(in[156] ^ in[159]); 
    assign layer_0[3166] = in[158]; 
    assign layer_0[3167] = in[215]; 
    assign layer_0[3168] = in[227]; 
    assign layer_0[3169] = ~(in[47] & in[72]); 
    assign layer_0[3170] = ~in[132] | (in[132] & in[25]); 
    assign layer_0[3171] = ~(in[12] ^ in[13]); 
    assign layer_0[3172] = in[50] & ~in[16]; 
    assign layer_0[3173] = in[109] | in[125]; 
    assign layer_0[3174] = in[220] ^ in[241]; 
    assign layer_0[3175] = ~(in[39] | in[131]); 
    assign layer_0[3176] = in[137] & ~in[158]; 
    assign layer_0[3177] = ~(in[160] ^ in[109]); 
    assign layer_0[3178] = ~(in[8] ^ in[109]); 
    assign layer_0[3179] = in[133]; 
    assign layer_0[3180] = in[114]; 
    assign layer_0[3181] = ~(in[135] | in[225]); 
    assign layer_0[3182] = in[105] & ~in[150]; 
    assign layer_0[3183] = ~in[229]; 
    assign layer_0[3184] = in[15]; 
    assign layer_0[3185] = ~in[190]; 
    assign layer_0[3186] = ~in[68]; 
    assign layer_0[3187] = ~in[117]; 
    assign layer_0[3188] = in[102] & ~in[206]; 
    assign layer_0[3189] = in[120] & ~in[220]; 
    assign layer_0[3190] = in[77]; 
    assign layer_0[3191] = ~(in[69] | in[18]); 
    assign layer_0[3192] = in[65] & in[62]; 
    assign layer_0[3193] = ~in[57] | (in[165] & in[57]); 
    assign layer_0[3194] = ~in[57]; 
    assign layer_0[3195] = ~(in[246] | in[244]); 
    assign layer_0[3196] = in[138] & ~in[38]; 
    assign layer_0[3197] = ~(in[113] & in[104]); 
    assign layer_0[3198] = in[40] & ~in[111]; 
    assign layer_0[3199] = in[102]; 
    assign layer_0[3200] = ~in[90] | (in[90] & in[147]); 
    assign layer_0[3201] = in[181] | in[167]; 
    assign layer_0[3202] = in[69]; 
    assign layer_0[3203] = ~in[91] | (in[91] & in[156]); 
    assign layer_0[3204] = in[140] ^ in[143]; 
    assign layer_0[3205] = ~(in[145] | in[118]); 
    assign layer_0[3206] = ~(in[225] | in[166]); 
    assign layer_0[3207] = ~in[187] | (in[187] & in[160]); 
    assign layer_0[3208] = in[137]; 
    assign layer_0[3209] = in[169]; 
    assign layer_0[3210] = in[254] | in[148]; 
    assign layer_0[3211] = ~in[152] | (in[84] & in[152]); 
    assign layer_0[3212] = in[112] | in[190]; 
    assign layer_0[3213] = in[100] | in[220]; 
    assign layer_0[3214] = in[98] ^ in[76]; 
    assign layer_0[3215] = in[133] | in[248]; 
    assign layer_0[3216] = ~in[40] | (in[40] & in[32]); 
    assign layer_0[3217] = ~in[37] | (in[4] & in[37]); 
    assign layer_0[3218] = ~(in[247] | in[226]); 
    assign layer_0[3219] = ~in[250]; 
    assign layer_0[3220] = in[212]; 
    assign layer_0[3221] = ~in[104]; 
    assign layer_0[3222] = ~(in[71] ^ in[172]); 
    assign layer_0[3223] = in[127] & ~in[36]; 
    assign layer_0[3224] = ~(in[119] | in[175]); 
    assign layer_0[3225] = in[138]; 
    assign layer_0[3226] = in[29] & in[119]; 
    assign layer_0[3227] = in[10] | in[89]; 
    assign layer_0[3228] = ~in[163] | (in[163] & in[46]); 
    assign layer_0[3229] = in[216] & in[252]; 
    assign layer_0[3230] = in[163] & ~in[99]; 
    assign layer_0[3231] = in[187] & ~in[62]; 
    assign layer_0[3232] = in[91] & ~in[15]; 
    assign layer_0[3233] = in[254] ^ in[206]; 
    assign layer_0[3234] = in[221] | in[212]; 
    assign layer_0[3235] = ~in[245]; 
    assign layer_0[3236] = ~in[67]; 
    assign layer_0[3237] = in[43] ^ in[137]; 
    assign layer_0[3238] = ~in[34]; 
    assign layer_0[3239] = ~(in[133] & in[118]); 
    assign layer_0[3240] = ~in[115]; 
    assign layer_0[3241] = in[22] | in[27]; 
    assign layer_0[3242] = in[150]; 
    assign layer_0[3243] = ~in[187] | (in[216] & in[187]); 
    assign layer_0[3244] = ~in[224] | (in[224] & in[166]); 
    assign layer_0[3245] = ~in[56] | (in[56] & in[20]); 
    assign layer_0[3246] = in[152] & ~in[227]; 
    assign layer_0[3247] = ~in[135]; 
    assign layer_0[3248] = in[249] ^ in[219]; 
    assign layer_0[3249] = ~(in[18] ^ in[139]); 
    assign layer_0[3250] = in[39]; 
    assign layer_0[3251] = in[190] & ~in[251]; 
    assign layer_0[3252] = ~(in[177] | in[152]); 
    assign layer_0[3253] = in[9] ^ in[50]; 
    assign layer_0[3254] = ~in[91] | (in[38] & in[91]); 
    assign layer_0[3255] = in[99]; 
    assign layer_0[3256] = ~in[197] | (in[248] & in[197]); 
    assign layer_0[3257] = in[186] ^ in[101]; 
    assign layer_0[3258] = in[212]; 
    assign layer_0[3259] = ~in[82] | (in[82] & in[78]); 
    assign layer_0[3260] = ~(in[236] | in[247]); 
    assign layer_0[3261] = ~in[152] | (in[39] & in[152]); 
    assign layer_0[3262] = ~(in[69] ^ in[171]); 
    assign layer_0[3263] = ~(in[198] | in[213]); 
    assign layer_0[3264] = in[180] & ~in[246]; 
    assign layer_0[3265] = ~(in[146] | in[192]); 
    assign layer_0[3266] = ~in[113]; 
    assign layer_0[3267] = ~(in[60] | in[79]); 
    assign layer_0[3268] = ~(in[81] & in[128]); 
    assign layer_0[3269] = in[203]; 
    assign layer_0[3270] = in[76] | in[60]; 
    assign layer_0[3271] = ~(in[205] & in[140]); 
    assign layer_0[3272] = ~in[160]; 
    assign layer_0[3273] = ~in[96]; 
    assign layer_0[3274] = in[70]; 
    assign layer_0[3275] = in[113] | in[146]; 
    assign layer_0[3276] = ~in[91] | (in[91] & in[43]); 
    assign layer_0[3277] = ~in[123]; 
    assign layer_0[3278] = in[237] & in[155]; 
    assign layer_0[3279] = ~(in[106] | in[135]); 
    assign layer_0[3280] = ~(in[248] & in[222]); 
    assign layer_0[3281] = ~(in[199] | in[97]); 
    assign layer_0[3282] = in[53] ^ in[71]; 
    assign layer_0[3283] = in[99] | in[160]; 
    assign layer_0[3284] = in[97]; 
    assign layer_0[3285] = ~(in[143] & in[179]); 
    assign layer_0[3286] = ~in[132] | (in[132] & in[20]); 
    assign layer_0[3287] = ~(in[155] ^ in[239]); 
    assign layer_0[3288] = in[111] & in[21]; 
    assign layer_0[3289] = in[121] & ~in[175]; 
    assign layer_0[3290] = ~in[116]; 
    assign layer_0[3291] = ~(in[28] | in[37]); 
    assign layer_0[3292] = in[142] | in[143]; 
    assign layer_0[3293] = in[25] ^ in[87]; 
    assign layer_0[3294] = in[198] ^ in[201]; 
    assign layer_0[3295] = in[142] | in[88]; 
    assign layer_0[3296] = in[173] | in[57]; 
    assign layer_0[3297] = in[154] & ~in[234]; 
    assign layer_0[3298] = ~(in[221] ^ in[112]); 
    assign layer_0[3299] = in[27] & ~in[3]; 
    assign layer_0[3300] = ~(in[164] | in[69]); 
    assign layer_0[3301] = ~(in[89] & in[201]); 
    assign layer_0[3302] = in[4] ^ in[27]; 
    assign layer_0[3303] = in[104] & in[155]; 
    assign layer_0[3304] = in[198]; 
    assign layer_0[3305] = in[72] & ~in[103]; 
    assign layer_0[3306] = ~(in[18] ^ in[78]); 
    assign layer_0[3307] = ~in[214]; 
    assign layer_0[3308] = in[79] ^ in[21]; 
    assign layer_0[3309] = ~(in[142] & in[60]); 
    assign layer_0[3310] = in[64] | in[159]; 
    assign layer_0[3311] = ~(in[104] | in[127]); 
    assign layer_0[3312] = ~(in[135] & in[121]); 
    assign layer_0[3313] = ~in[5] | (in[5] & in[11]); 
    assign layer_0[3314] = in[119] | in[27]; 
    assign layer_0[3315] = in[82] ^ in[8]; 
    assign layer_0[3316] = in[170] | in[192]; 
    assign layer_0[3317] = ~(in[18] | in[37]); 
    assign layer_0[3318] = ~(in[6] & in[58]); 
    assign layer_0[3319] = in[242] ^ in[245]; 
    assign layer_0[3320] = ~in[78]; 
    assign layer_0[3321] = in[209] | in[228]; 
    assign layer_0[3322] = in[186] & ~in[97]; 
    assign layer_0[3323] = ~in[214]; 
    assign layer_0[3324] = in[101] & in[58]; 
    assign layer_0[3325] = in[100] & ~in[79]; 
    assign layer_0[3326] = ~(in[69] | in[108]); 
    assign layer_0[3327] = in[251] ^ in[159]; 
    assign layer_0[3328] = ~(in[127] & in[221]); 
    assign layer_0[3329] = in[126] | in[157]; 
    assign layer_0[3330] = in[109] & in[47]; 
    assign layer_0[3331] = ~(in[21] | in[3]); 
    assign layer_0[3332] = in[197] & ~in[138]; 
    assign layer_0[3333] = in[133]; 
    assign layer_0[3334] = ~(in[210] ^ in[143]); 
    assign layer_0[3335] = in[155] & ~in[50]; 
    assign layer_0[3336] = ~in[212] | (in[212] & in[176]); 
    assign layer_0[3337] = ~in[153]; 
    assign layer_0[3338] = ~in[52] | (in[52] & in[153]); 
    assign layer_0[3339] = ~(in[182] | in[82]); 
    assign layer_0[3340] = in[202]; 
    assign layer_0[3341] = in[82] | in[18]; 
    assign layer_0[3342] = ~in[92]; 
    assign layer_0[3343] = ~in[182]; 
    assign layer_0[3344] = in[3] & ~in[54]; 
    assign layer_0[3345] = ~in[139] | (in[139] & in[146]); 
    assign layer_0[3346] = ~in[141] | (in[224] & in[141]); 
    assign layer_0[3347] = ~in[147]; 
    assign layer_0[3348] = in[37] | in[40]; 
    assign layer_0[3349] = ~(in[215] | in[159]); 
    assign layer_0[3350] = in[31]; 
    assign layer_0[3351] = ~(in[148] & in[200]); 
    assign layer_0[3352] = in[124] ^ in[43]; 
    assign layer_0[3353] = in[4] ^ in[119]; 
    assign layer_0[3354] = ~in[186] | (in[140] & in[186]); 
    assign layer_0[3355] = in[149] & ~in[193]; 
    assign layer_0[3356] = in[122] ^ in[229]; 
    assign layer_0[3357] = ~in[253]; 
    assign layer_0[3358] = in[158]; 
    assign layer_0[3359] = in[171] & ~in[201]; 
    assign layer_0[3360] = ~in[46] | (in[46] & in[99]); 
    assign layer_0[3361] = ~in[180]; 
    assign layer_0[3362] = ~in[88] | (in[88] & in[94]); 
    assign layer_0[3363] = in[61] & ~in[11]; 
    assign layer_0[3364] = in[196] | in[210]; 
    assign layer_0[3365] = ~(in[204] | in[164]); 
    assign layer_0[3366] = in[138]; 
    assign layer_0[3367] = ~in[100]; 
    assign layer_0[3368] = in[174] ^ in[170]; 
    assign layer_0[3369] = ~(in[90] ^ in[197]); 
    assign layer_0[3370] = in[2]; 
    assign layer_0[3371] = ~in[107] | (in[68] & in[107]); 
    assign layer_0[3372] = ~(in[245] | in[213]); 
    assign layer_0[3373] = in[171] & ~in[163]; 
    assign layer_0[3374] = ~(in[241] | in[250]); 
    assign layer_0[3375] = in[97]; 
    assign layer_0[3376] = ~(in[85] & in[91]); 
    assign layer_0[3377] = in[187] & in[207]; 
    assign layer_0[3378] = ~(in[173] ^ in[163]); 
    assign layer_0[3379] = ~(in[30] | in[25]); 
    assign layer_0[3380] = ~in[163] | (in[163] & in[225]); 
    assign layer_0[3381] = in[209] ^ in[218]; 
    assign layer_0[3382] = ~in[39]; 
    assign layer_0[3383] = in[94] | in[108]; 
    assign layer_0[3384] = ~(in[145] & in[18]); 
    assign layer_0[3385] = in[31] | in[126]; 
    assign layer_0[3386] = ~in[51] | (in[1] & in[51]); 
    assign layer_0[3387] = ~in[148]; 
    assign layer_0[3388] = ~(in[73] & in[108]); 
    assign layer_0[3389] = ~in[27]; 
    assign layer_0[3390] = ~in[184] | (in[75] & in[184]); 
    assign layer_0[3391] = ~in[51]; 
    assign layer_0[3392] = ~(in[219] & in[235]); 
    assign layer_0[3393] = in[118] & ~in[210]; 
    assign layer_0[3394] = in[138] | in[254]; 
    assign layer_0[3395] = in[204] | in[148]; 
    assign layer_0[3396] = in[171]; 
    assign layer_0[3397] = in[72]; 
    assign layer_0[3398] = ~in[152] | (in[229] & in[152]); 
    assign layer_0[3399] = ~in[132]; 
    assign layer_0[3400] = ~in[38] | (in[38] & in[40]); 
    assign layer_0[3401] = in[90]; 
    assign layer_0[3402] = ~in[123]; 
    assign layer_0[3403] = in[66] ^ in[59]; 
    assign layer_0[3404] = ~in[129]; 
    assign layer_0[3405] = ~in[88]; 
    assign layer_0[3406] = in[218] & ~in[233]; 
    assign layer_0[3407] = in[79] ^ in[38]; 
    assign layer_0[3408] = in[45]; 
    assign layer_0[3409] = ~(in[139] ^ in[15]); 
    assign layer_0[3410] = ~(in[200] | in[147]); 
    assign layer_0[3411] = in[76] ^ in[145]; 
    assign layer_0[3412] = in[154] & ~in[186]; 
    assign layer_0[3413] = in[229] & in[188]; 
    assign layer_0[3414] = in[227] | in[137]; 
    assign layer_0[3415] = in[46] | in[5]; 
    assign layer_0[3416] = ~in[118]; 
    assign layer_0[3417] = in[26] ^ in[57]; 
    assign layer_0[3418] = in[248]; 
    assign layer_0[3419] = in[224] ^ in[228]; 
    assign layer_0[3420] = in[67] | in[143]; 
    assign layer_0[3421] = ~(in[74] & in[52]); 
    assign layer_0[3422] = ~in[118] | (in[201] & in[118]); 
    assign layer_0[3423] = in[179]; 
    assign layer_0[3424] = ~in[219] | (in[219] & in[96]); 
    assign layer_0[3425] = in[40] & in[118]; 
    assign layer_0[3426] = in[25] ^ in[86]; 
    assign layer_0[3427] = ~in[120]; 
    assign layer_0[3428] = ~in[104] | (in[30] & in[104]); 
    assign layer_0[3429] = in[95] | in[190]; 
    assign layer_0[3430] = in[40]; 
    assign layer_0[3431] = in[230] & ~in[222]; 
    assign layer_0[3432] = in[38] & in[30]; 
    assign layer_0[3433] = ~in[110] | (in[36] & in[110]); 
    assign layer_0[3434] = in[86] & ~in[113]; 
    assign layer_0[3435] = ~(in[21] | in[60]); 
    assign layer_0[3436] = in[48] ^ in[60]; 
    assign layer_0[3437] = ~(in[86] & in[140]); 
    assign layer_0[3438] = in[76] & ~in[49]; 
    assign layer_0[3439] = ~in[121] | (in[121] & in[109]); 
    assign layer_0[3440] = in[60] | in[106]; 
    assign layer_0[3441] = ~(in[95] ^ in[220]); 
    assign layer_0[3442] = ~in[71]; 
    assign layer_0[3443] = ~in[36]; 
    assign layer_0[3444] = ~in[170]; 
    assign layer_0[3445] = in[163] | in[171]; 
    assign layer_0[3446] = in[103] & ~in[1]; 
    assign layer_0[3447] = ~in[212] | (in[212] & in[200]); 
    assign layer_0[3448] = in[63]; 
    assign layer_0[3449] = in[89]; 
    assign layer_0[3450] = in[18] ^ in[63]; 
    assign layer_0[3451] = in[54] & ~in[99]; 
    assign layer_0[3452] = in[185]; 
    assign layer_0[3453] = in[91]; 
    assign layer_0[3454] = ~in[60]; 
    assign layer_0[3455] = ~(in[148] | in[140]); 
    assign layer_0[3456] = in[87] ^ in[38]; 
    assign layer_0[3457] = in[119] & in[155]; 
    assign layer_0[3458] = in[152] & ~in[28]; 
    assign layer_0[3459] = ~(in[72] & in[166]); 
    assign layer_0[3460] = in[96] & in[20]; 
    assign layer_0[3461] = ~in[222] | (in[222] & in[99]); 
    assign layer_0[3462] = ~(in[214] & in[121]); 
    assign layer_0[3463] = ~in[159]; 
    assign layer_0[3464] = in[192] | in[182]; 
    assign layer_0[3465] = ~(in[248] | in[182]); 
    assign layer_0[3466] = in[248] ^ in[140]; 
    assign layer_0[3467] = ~(in[64] ^ in[144]); 
    assign layer_0[3468] = ~in[55]; 
    assign layer_0[3469] = in[175]; 
    assign layer_0[3470] = in[59] & ~in[176]; 
    assign layer_0[3471] = ~in[178]; 
    assign layer_0[3472] = in[230]; 
    assign layer_0[3473] = in[157]; 
    assign layer_0[3474] = ~in[54] | (in[29] & in[54]); 
    assign layer_0[3475] = ~(in[85] | in[47]); 
    assign layer_0[3476] = ~in[40]; 
    assign layer_0[3477] = in[108]; 
    assign layer_0[3478] = in[136]; 
    assign layer_0[3479] = ~in[49]; 
    assign layer_0[3480] = in[33] ^ in[95]; 
    assign layer_0[3481] = ~in[65]; 
    assign layer_0[3482] = ~(in[232] ^ in[194]); 
    assign layer_0[3483] = ~in[100]; 
    assign layer_0[3484] = ~(in[83] | in[123]); 
    assign layer_0[3485] = ~(in[221] | in[229]); 
    assign layer_0[3486] = in[62]; 
    assign layer_0[3487] = in[200] ^ in[97]; 
    assign layer_0[3488] = in[9] & ~in[47]; 
    assign layer_0[3489] = in[63] ^ in[52]; 
    assign layer_0[3490] = ~(in[104] & in[165]); 
    assign layer_0[3491] = ~(in[211] ^ in[160]); 
    assign layer_0[3492] = ~in[38] | (in[38] & in[27]); 
    assign layer_0[3493] = ~(in[119] | in[97]); 
    assign layer_0[3494] = in[40]; 
    assign layer_0[3495] = in[198] | in[79]; 
    assign layer_0[3496] = ~(in[254] | in[171]); 
    assign layer_0[3497] = ~(in[170] & in[95]); 
    assign layer_0[3498] = in[160] | in[218]; 
    assign layer_0[3499] = in[192]; 
    assign layer_0[3500] = ~in[142] | (in[142] & in[96]); 
    assign layer_0[3501] = in[149]; 
    assign layer_0[3502] = in[254] ^ in[193]; 
    assign layer_0[3503] = ~(in[44] | in[146]); 
    assign layer_0[3504] = ~(in[17] & in[118]); 
    assign layer_0[3505] = ~(in[150] | in[161]); 
    assign layer_0[3506] = ~(in[13] ^ in[7]); 
    assign layer_0[3507] = in[69] | in[175]; 
    assign layer_0[3508] = in[192] & ~in[223]; 
    assign layer_0[3509] = in[196]; 
    assign layer_0[3510] = in[85]; 
    assign layer_0[3511] = in[193] | in[173]; 
    assign layer_0[3512] = in[90] & ~in[43]; 
    assign layer_0[3513] = ~in[90] | (in[53] & in[90]); 
    assign layer_0[3514] = ~in[44] | (in[44] & in[108]); 
    assign layer_0[3515] = ~(in[57] & in[116]); 
    assign layer_0[3516] = in[180]; 
    assign layer_0[3517] = ~(in[107] & in[119]); 
    assign layer_0[3518] = ~(in[62] & in[74]); 
    assign layer_0[3519] = in[117] & ~in[52]; 
    assign layer_0[3520] = ~in[171] | (in[171] & in[168]); 
    assign layer_0[3521] = in[149] ^ in[210]; 
    assign layer_0[3522] = ~(in[233] & in[114]); 
    assign layer_0[3523] = in[208] | in[247]; 
    assign layer_0[3524] = ~in[231]; 
    assign layer_0[3525] = ~in[2]; 
    assign layer_0[3526] = in[119] & ~in[69]; 
    assign layer_0[3527] = ~in[88] | (in[88] & in[115]); 
    assign layer_0[3528] = ~in[172] | (in[50] & in[172]); 
    assign layer_0[3529] = ~in[110] | (in[110] & in[222]); 
    assign layer_0[3530] = ~in[227] | (in[227] & in[163]); 
    assign layer_0[3531] = in[182] | in[223]; 
    assign layer_0[3532] = ~(in[234] ^ in[244]); 
    assign layer_0[3533] = ~(in[134] & in[105]); 
    assign layer_0[3534] = in[233] & in[117]; 
    assign layer_0[3535] = ~(in[52] | in[156]); 
    assign layer_0[3536] = in[66] | in[128]; 
    assign layer_0[3537] = ~in[8]; 
    assign layer_0[3538] = in[108] & in[188]; 
    assign layer_0[3539] = ~(in[240] | in[122]); 
    assign layer_0[3540] = ~in[86]; 
    assign layer_0[3541] = ~in[127]; 
    assign layer_0[3542] = in[137] & ~in[54]; 
    assign layer_0[3543] = in[133]; 
    assign layer_0[3544] = ~(in[214] ^ in[219]); 
    assign layer_0[3545] = ~(in[218] ^ in[121]); 
    assign layer_0[3546] = ~(in[37] ^ in[86]); 
    assign layer_0[3547] = ~in[70]; 
    assign layer_0[3548] = in[152] & ~in[211]; 
    assign layer_0[3549] = in[65] ^ in[145]; 
    assign layer_0[3550] = in[95] | in[54]; 
    assign layer_0[3551] = ~(in[194] ^ in[233]); 
    assign layer_0[3552] = ~in[224] | (in[224] & in[201]); 
    assign layer_0[3553] = ~in[216]; 
    assign layer_0[3554] = in[189] & in[165]; 
    assign layer_0[3555] = ~in[243]; 
    assign layer_0[3556] = in[232]; 
    assign layer_0[3557] = in[113] & ~in[73]; 
    assign layer_0[3558] = in[29] | in[138]; 
    assign layer_0[3559] = in[229] | in[223]; 
    assign layer_0[3560] = in[180] & ~in[150]; 
    assign layer_0[3561] = in[71] & ~in[154]; 
    assign layer_0[3562] = ~(in[207] ^ in[98]); 
    assign layer_0[3563] = ~in[110] | (in[235] & in[110]); 
    assign layer_0[3564] = in[244] & ~in[208]; 
    assign layer_0[3565] = in[66] ^ in[142]; 
    assign layer_0[3566] = ~in[176]; 
    assign layer_0[3567] = in[5]; 
    assign layer_0[3568] = in[120] | in[69]; 
    assign layer_0[3569] = ~(in[37] & in[5]); 
    assign layer_0[3570] = in[59] & ~in[46]; 
    assign layer_0[3571] = ~in[96]; 
    assign layer_0[3572] = ~in[57] | (in[160] & in[57]); 
    assign layer_0[3573] = ~in[155]; 
    assign layer_0[3574] = in[16] ^ in[38]; 
    assign layer_0[3575] = ~in[87] | (in[159] & in[87]); 
    assign layer_0[3576] = in[59] ^ in[44]; 
    assign layer_0[3577] = in[33] & ~in[63]; 
    assign layer_0[3578] = in[89] & in[106]; 
    assign layer_0[3579] = ~in[39] | (in[39] & in[117]); 
    assign layer_0[3580] = in[246] | in[126]; 
    assign layer_0[3581] = ~in[186] | (in[206] & in[186]); 
    assign layer_0[3582] = in[159] ^ in[87]; 
    assign layer_0[3583] = in[188] & ~in[114]; 
    assign layer_0[3584] = ~in[133] | (in[157] & in[133]); 
    assign layer_0[3585] = in[108] & ~in[41]; 
    assign layer_0[3586] = in[128] & ~in[251]; 
    assign layer_0[3587] = in[134]; 
    assign layer_0[3588] = ~in[133]; 
    assign layer_0[3589] = ~in[132]; 
    assign layer_0[3590] = in[183] | in[255]; 
    assign layer_0[3591] = in[153]; 
    assign layer_0[3592] = in[38] ^ in[3]; 
    assign layer_0[3593] = ~(in[183] ^ in[240]); 
    assign layer_0[3594] = ~in[84] | (in[21] & in[84]); 
    assign layer_0[3595] = ~(in[139] ^ in[153]); 
    assign layer_0[3596] = in[119] & ~in[70]; 
    assign layer_0[3597] = ~in[210] | (in[210] & in[121]); 
    assign layer_0[3598] = in[14] | in[61]; 
    assign layer_0[3599] = in[163] ^ in[121]; 
    assign layer_0[3600] = in[156] & ~in[139]; 
    assign layer_0[3601] = ~(in[173] ^ in[53]); 
    assign layer_0[3602] = in[222] ^ in[103]; 
    assign layer_0[3603] = in[152] & ~in[144]; 
    assign layer_0[3604] = ~in[89]; 
    assign layer_0[3605] = in[58] & ~in[79]; 
    assign layer_0[3606] = in[225] | in[207]; 
    assign layer_0[3607] = in[53]; 
    assign layer_0[3608] = ~in[197]; 
    assign layer_0[3609] = in[27] ^ in[60]; 
    assign layer_0[3610] = in[186]; 
    assign layer_0[3611] = ~in[182]; 
    assign layer_0[3612] = ~(in[226] | in[239]); 
    assign layer_0[3613] = in[201]; 
    assign layer_0[3614] = ~in[42]; 
    assign layer_0[3615] = ~in[150] | (in[150] & in[210]); 
    assign layer_0[3616] = in[34]; 
    assign layer_0[3617] = in[98]; 
    assign layer_0[3618] = ~in[125] | (in[125] & in[127]); 
    assign layer_0[3619] = ~in[172] | (in[239] & in[172]); 
    assign layer_0[3620] = in[132] & ~in[129]; 
    assign layer_0[3621] = ~in[127]; 
    assign layer_0[3622] = in[158]; 
    assign layer_0[3623] = ~(in[207] ^ in[87]); 
    assign layer_0[3624] = ~(in[16] | in[4]); 
    assign layer_0[3625] = in[19] | in[125]; 
    assign layer_0[3626] = ~(in[115] | in[24]); 
    assign layer_0[3627] = ~in[112] | (in[112] & in[146]); 
    assign layer_0[3628] = ~in[119] | (in[194] & in[119]); 
    assign layer_0[3629] = ~in[100]; 
    assign layer_0[3630] = in[12]; 
    assign layer_0[3631] = ~in[100] | (in[100] & in[210]); 
    assign layer_0[3632] = ~(in[238] | in[209]); 
    assign layer_0[3633] = in[30] | in[155]; 
    assign layer_0[3634] = ~(in[138] ^ in[227]); 
    assign layer_0[3635] = in[47]; 
    assign layer_0[3636] = in[214] ^ in[202]; 
    assign layer_0[3637] = ~in[75]; 
    assign layer_0[3638] = in[58] & ~in[142]; 
    assign layer_0[3639] = in[52]; 
    assign layer_0[3640] = ~(in[44] & in[141]); 
    assign layer_0[3641] = in[170]; 
    assign layer_0[3642] = in[124]; 
    assign layer_0[3643] = ~(in[145] | in[42]); 
    assign layer_0[3644] = ~(in[191] ^ in[96]); 
    assign layer_0[3645] = ~in[14]; 
    assign layer_0[3646] = ~in[165] | (in[244] & in[165]); 
    assign layer_0[3647] = ~(in[128] & in[169]); 
    assign layer_0[3648] = in[136]; 
    assign layer_0[3649] = ~in[27] | (in[110] & in[27]); 
    assign layer_0[3650] = in[158] | in[149]; 
    assign layer_0[3651] = in[94] | in[49]; 
    assign layer_0[3652] = ~in[202]; 
    assign layer_0[3653] = ~in[132] | (in[132] & in[83]); 
    assign layer_0[3654] = ~in[15]; 
    assign layer_0[3655] = ~(in[130] ^ in[52]); 
    assign layer_0[3656] = ~in[25]; 
    assign layer_0[3657] = in[114] | in[84]; 
    assign layer_0[3658] = in[236]; 
    assign layer_0[3659] = in[155]; 
    assign layer_0[3660] = ~in[76]; 
    assign layer_0[3661] = in[43]; 
    assign layer_0[3662] = in[99]; 
    assign layer_0[3663] = in[217] & ~in[112]; 
    assign layer_0[3664] = ~in[96] | (in[96] & in[118]); 
    assign layer_0[3665] = ~(in[63] & in[145]); 
    assign layer_0[3666] = ~(in[219] | in[133]); 
    assign layer_0[3667] = in[218]; 
    assign layer_0[3668] = ~(in[103] & in[109]); 
    assign layer_0[3669] = in[134] & ~in[236]; 
    assign layer_0[3670] = ~in[209] | (in[209] & in[172]); 
    assign layer_0[3671] = ~in[156]; 
    assign layer_0[3672] = in[196] & in[140]; 
    assign layer_0[3673] = in[112] | in[210]; 
    assign layer_0[3674] = ~(in[175] | in[168]); 
    assign layer_0[3675] = ~in[175] | (in[175] & in[173]); 
    assign layer_0[3676] = ~in[59]; 
    assign layer_0[3677] = in[98] ^ in[186]; 
    assign layer_0[3678] = in[26]; 
    assign layer_0[3679] = in[47] ^ in[52]; 
    assign layer_0[3680] = ~in[253] | (in[253] & in[176]); 
    assign layer_0[3681] = in[178]; 
    assign layer_0[3682] = in[141] | in[175]; 
    assign layer_0[3683] = ~in[162] | (in[232] & in[162]); 
    assign layer_0[3684] = in[225] | in[187]; 
    assign layer_0[3685] = in[220] & ~in[95]; 
    assign layer_0[3686] = ~(in[35] & in[31]); 
    assign layer_0[3687] = in[189] | in[204]; 
    assign layer_0[3688] = ~(in[76] & in[78]); 
    assign layer_0[3689] = ~in[56]; 
    assign layer_0[3690] = in[82]; 
    assign layer_0[3691] = ~(in[254] | in[166]); 
    assign layer_0[3692] = ~in[143] | (in[224] & in[143]); 
    assign layer_0[3693] = ~in[14]; 
    assign layer_0[3694] = ~(in[213] ^ in[219]); 
    assign layer_0[3695] = ~in[122]; 
    assign layer_0[3696] = in[240] ^ in[220]; 
    assign layer_0[3697] = in[78] | in[109]; 
    assign layer_0[3698] = in[10] & in[0]; 
    assign layer_0[3699] = ~in[54]; 
    assign layer_0[3700] = ~(in[161] ^ in[133]); 
    assign layer_0[3701] = in[61]; 
    assign layer_0[3702] = ~in[121] | (in[159] & in[121]); 
    assign layer_0[3703] = ~in[108] | (in[52] & in[108]); 
    assign layer_0[3704] = ~in[154] | (in[131] & in[154]); 
    assign layer_0[3705] = in[213] ^ in[174]; 
    assign layer_0[3706] = ~in[57] | (in[57] & in[135]); 
    assign layer_0[3707] = in[16]; 
    assign layer_0[3708] = in[235] & in[225]; 
    assign layer_0[3709] = in[168] & ~in[229]; 
    assign layer_0[3710] = ~in[134]; 
    assign layer_0[3711] = in[227] & ~in[126]; 
    assign layer_0[3712] = ~in[63]; 
    assign layer_0[3713] = in[75] & ~in[123]; 
    assign layer_0[3714] = in[56]; 
    assign layer_0[3715] = in[187]; 
    assign layer_0[3716] = in[77] & ~in[100]; 
    assign layer_0[3717] = in[251] | in[164]; 
    assign layer_0[3718] = ~(in[85] & in[193]); 
    assign layer_0[3719] = in[192]; 
    assign layer_0[3720] = in[183]; 
    assign layer_0[3721] = in[243] & in[249]; 
    assign layer_0[3722] = in[57]; 
    assign layer_0[3723] = ~in[133] | (in[133] & in[93]); 
    assign layer_0[3724] = in[214]; 
    assign layer_0[3725] = in[70] & ~in[112]; 
    assign layer_0[3726] = in[86]; 
    assign layer_0[3727] = in[167] & ~in[174]; 
    assign layer_0[3728] = ~(in[7] & in[100]); 
    assign layer_0[3729] = in[132]; 
    assign layer_0[3730] = ~(in[167] | in[151]); 
    assign layer_0[3731] = ~in[147]; 
    assign layer_0[3732] = ~in[196]; 
    assign layer_0[3733] = ~(in[251] | in[171]); 
    assign layer_0[3734] = in[189] & ~in[106]; 
    assign layer_0[3735] = in[176] ^ in[143]; 
    assign layer_0[3736] = ~(in[145] & in[112]); 
    assign layer_0[3737] = ~in[195] | (in[226] & in[195]); 
    assign layer_0[3738] = ~in[217] | (in[217] & in[221]); 
    assign layer_0[3739] = ~in[159] | (in[159] & in[107]); 
    assign layer_0[3740] = ~in[235]; 
    assign layer_0[3741] = ~in[171] | (in[100] & in[171]); 
    assign layer_0[3742] = in[232] | in[138]; 
    assign layer_0[3743] = ~(in[7] ^ in[54]); 
    assign layer_0[3744] = in[142] | in[125]; 
    assign layer_0[3745] = in[32] | in[97]; 
    assign layer_0[3746] = ~in[9]; 
    assign layer_0[3747] = in[213] | in[217]; 
    assign layer_0[3748] = ~(in[130] | in[17]); 
    assign layer_0[3749] = in[29] & ~in[62]; 
    assign layer_0[3750] = ~(in[35] | in[12]); 
    assign layer_0[3751] = ~in[34]; 
    assign layer_0[3752] = in[158] | in[169]; 
    assign layer_0[3753] = ~in[204]; 
    assign layer_0[3754] = ~(in[241] & in[203]); 
    assign layer_0[3755] = ~in[129] | (in[4] & in[129]); 
    assign layer_0[3756] = in[31]; 
    assign layer_0[3757] = ~(in[164] ^ in[131]); 
    assign layer_0[3758] = ~(in[83] ^ in[179]); 
    assign layer_0[3759] = in[187] ^ in[166]; 
    assign layer_0[3760] = ~in[72] | (in[165] & in[72]); 
    assign layer_0[3761] = ~in[84] | (in[84] & in[62]); 
    assign layer_0[3762] = ~in[223]; 
    assign layer_0[3763] = ~(in[122] | in[0]); 
    assign layer_0[3764] = in[3] | in[41]; 
    assign layer_0[3765] = in[87] ^ in[212]; 
    assign layer_0[3766] = ~(in[44] & in[113]); 
    assign layer_0[3767] = in[83] ^ in[190]; 
    assign layer_0[3768] = in[146] ^ in[103]; 
    assign layer_0[3769] = in[45]; 
    assign layer_0[3770] = in[48]; 
    assign layer_0[3771] = in[123]; 
    assign layer_0[3772] = ~(in[163] ^ in[148]); 
    assign layer_0[3773] = ~in[0] | (in[7] & in[0]); 
    assign layer_0[3774] = in[83]; 
    assign layer_0[3775] = ~in[242] | (in[161] & in[242]); 
    assign layer_0[3776] = in[72] & ~in[35]; 
    assign layer_0[3777] = ~(in[224] ^ in[172]); 
    assign layer_0[3778] = in[201] & in[118]; 
    assign layer_0[3779] = in[203] ^ in[171]; 
    assign layer_0[3780] = ~in[192] | (in[192] & in[181]); 
    assign layer_0[3781] = in[12] & ~in[1]; 
    assign layer_0[3782] = ~in[182] | (in[182] & in[125]); 
    assign layer_0[3783] = in[200] & ~in[255]; 
    assign layer_0[3784] = ~(in[233] & in[145]); 
    assign layer_0[3785] = in[7] ^ in[92]; 
    assign layer_0[3786] = in[172]; 
    assign layer_0[3787] = ~(in[180] | in[225]); 
    assign layer_0[3788] = ~in[83]; 
    assign layer_0[3789] = in[13] & ~in[4]; 
    assign layer_0[3790] = in[103]; 
    assign layer_0[3791] = ~in[102]; 
    assign layer_0[3792] = in[181] ^ in[136]; 
    assign layer_0[3793] = in[141] & ~in[192]; 
    assign layer_0[3794] = ~in[107] | (in[107] & in[33]); 
    assign layer_0[3795] = in[189] | in[194]; 
    assign layer_0[3796] = in[125]; 
    assign layer_0[3797] = in[110] & in[92]; 
    assign layer_0[3798] = ~in[72]; 
    assign layer_0[3799] = ~(in[133] | in[252]); 
    assign layer_0[3800] = ~(in[71] & in[101]); 
    assign layer_0[3801] = ~in[109]; 
    assign layer_0[3802] = in[159] & ~in[240]; 
    assign layer_0[3803] = ~in[146] | (in[218] & in[146]); 
    assign layer_0[3804] = ~in[5] | (in[5] & in[9]); 
    assign layer_0[3805] = in[195] | in[239]; 
    assign layer_0[3806] = in[138] | in[17]; 
    assign layer_0[3807] = in[168]; 
    assign layer_0[3808] = in[242] & ~in[201]; 
    assign layer_0[3809] = ~in[136] | (in[136] & in[42]); 
    assign layer_0[3810] = ~(in[38] & in[94]); 
    assign layer_0[3811] = ~(in[162] & in[241]); 
    assign layer_0[3812] = in[13]; 
    assign layer_0[3813] = ~in[40]; 
    assign layer_0[3814] = in[116] & ~in[157]; 
    assign layer_0[3815] = ~(in[89] & in[117]); 
    assign layer_0[3816] = in[156] & ~in[249]; 
    assign layer_0[3817] = ~in[52] | (in[52] & in[4]); 
    assign layer_0[3818] = ~in[31] | (in[21] & in[31]); 
    assign layer_0[3819] = ~in[48]; 
    assign layer_0[3820] = ~in[133]; 
    assign layer_0[3821] = ~in[68] | (in[68] & in[0]); 
    assign layer_0[3822] = ~in[138]; 
    assign layer_0[3823] = in[168]; 
    assign layer_0[3824] = ~(in[161] | in[44]); 
    assign layer_0[3825] = ~(in[21] | in[51]); 
    assign layer_0[3826] = in[177] ^ in[214]; 
    assign layer_0[3827] = ~(in[171] | in[134]); 
    assign layer_0[3828] = in[218] ^ in[121]; 
    assign layer_0[3829] = ~(in[171] & in[59]); 
    assign layer_0[3830] = in[29] & in[69]; 
    assign layer_0[3831] = ~in[154] | (in[186] & in[154]); 
    assign layer_0[3832] = in[27]; 
    assign layer_0[3833] = in[156] & ~in[32]; 
    assign layer_0[3834] = in[212]; 
    assign layer_0[3835] = in[238] | in[168]; 
    assign layer_0[3836] = ~in[95]; 
    assign layer_0[3837] = in[106] ^ in[234]; 
    assign layer_0[3838] = ~in[166]; 
    assign layer_0[3839] = ~in[93]; 
    assign layer_0[3840] = in[89] & ~in[177]; 
    assign layer_0[3841] = in[34] & ~in[75]; 
    assign layer_0[3842] = in[102]; 
    assign layer_0[3843] = in[3] | in[17]; 
    assign layer_0[3844] = ~(in[41] | in[9]); 
    assign layer_0[3845] = in[154]; 
    assign layer_0[3846] = ~in[12] | (in[12] & in[46]); 
    assign layer_0[3847] = ~in[205]; 
    assign layer_0[3848] = ~(in[122] ^ in[155]); 
    assign layer_0[3849] = in[210] ^ in[165]; 
    assign layer_0[3850] = ~(in[199] | in[147]); 
    assign layer_0[3851] = in[226] & ~in[106]; 
    assign layer_0[3852] = ~in[121] | (in[226] & in[121]); 
    assign layer_0[3853] = ~in[150]; 
    assign layer_0[3854] = ~(in[209] ^ in[213]); 
    assign layer_0[3855] = in[160] & in[180]; 
    assign layer_0[3856] = ~in[99] | (in[99] & in[4]); 
    assign layer_0[3857] = ~(in[141] & in[149]); 
    assign layer_0[3858] = in[42]; 
    assign layer_0[3859] = ~(in[73] | in[1]); 
    assign layer_0[3860] = ~in[229] | (in[229] & in[221]); 
    assign layer_0[3861] = in[187]; 
    assign layer_0[3862] = ~(in[117] ^ in[129]); 
    assign layer_0[3863] = ~in[187] | (in[144] & in[187]); 
    assign layer_0[3864] = in[145]; 
    assign layer_0[3865] = in[84]; 
    assign layer_0[3866] = in[231] & ~in[174]; 
    assign layer_0[3867] = ~(in[200] ^ in[225]); 
    assign layer_0[3868] = in[139] & in[32]; 
    assign layer_0[3869] = in[92] | in[173]; 
    assign layer_0[3870] = in[82] & ~in[75]; 
    assign layer_0[3871] = in[128] ^ in[49]; 
    assign layer_0[3872] = ~(in[77] | in[189]); 
    assign layer_0[3873] = ~in[249] | (in[249] & in[218]); 
    assign layer_0[3874] = in[120] & ~in[218]; 
    assign layer_0[3875] = in[8]; 
    assign layer_0[3876] = in[52] & in[154]; 
    assign layer_0[3877] = ~in[147]; 
    assign layer_0[3878] = ~in[72] | (in[72] & in[11]); 
    assign layer_0[3879] = in[247] | in[200]; 
    assign layer_0[3880] = in[99]; 
    assign layer_0[3881] = ~in[30] | (in[30] & in[42]); 
    assign layer_0[3882] = ~(in[74] & in[165]); 
    assign layer_0[3883] = in[133] & ~in[170]; 
    assign layer_0[3884] = in[153] ^ in[188]; 
    assign layer_0[3885] = in[39]; 
    assign layer_0[3886] = in[252] & in[238]; 
    assign layer_0[3887] = in[62] & ~in[189]; 
    assign layer_0[3888] = ~(in[206] | in[191]); 
    assign layer_0[3889] = ~in[58] | (in[121] & in[58]); 
    assign layer_0[3890] = ~in[123] | (in[112] & in[123]); 
    assign layer_0[3891] = in[250] & ~in[235]; 
    assign layer_0[3892] = in[156] & ~in[216]; 
    assign layer_0[3893] = ~(in[207] ^ in[129]); 
    assign layer_0[3894] = ~in[194] | (in[146] & in[194]); 
    assign layer_0[3895] = ~(in[179] ^ in[149]); 
    assign layer_0[3896] = ~in[173]; 
    assign layer_0[3897] = in[253] & ~in[177]; 
    assign layer_0[3898] = in[187] & in[172]; 
    assign layer_0[3899] = ~in[55] | (in[55] & in[83]); 
    assign layer_0[3900] = ~(in[202] ^ in[180]); 
    assign layer_0[3901] = in[69] & ~in[120]; 
    assign layer_0[3902] = in[75] | in[51]; 
    assign layer_0[3903] = ~(in[94] ^ in[172]); 
    assign layer_0[3904] = ~in[7]; 
    assign layer_0[3905] = in[229] | in[242]; 
    assign layer_0[3906] = ~in[119]; 
    assign layer_0[3907] = ~in[180]; 
    assign layer_0[3908] = in[245] | in[202]; 
    assign layer_0[3909] = ~in[205] | (in[205] & in[201]); 
    assign layer_0[3910] = ~(in[229] ^ in[176]); 
    assign layer_0[3911] = ~in[133] | (in[133] & in[197]); 
    assign layer_0[3912] = in[220]; 
    assign layer_0[3913] = in[233] ^ in[183]; 
    assign layer_0[3914] = in[81] ^ in[89]; 
    assign layer_0[3915] = ~(in[83] & in[34]); 
    assign layer_0[3916] = ~(in[249] | in[201]); 
    assign layer_0[3917] = ~in[193]; 
    assign layer_0[3918] = ~in[44]; 
    assign layer_0[3919] = ~in[90] | (in[212] & in[90]); 
    assign layer_0[3920] = in[88] ^ in[153]; 
    assign layer_0[3921] = ~(in[201] & in[212]); 
    assign layer_0[3922] = in[241]; 
    assign layer_0[3923] = ~in[66] | (in[62] & in[66]); 
    assign layer_0[3924] = ~in[92] | (in[220] & in[92]); 
    assign layer_0[3925] = ~(in[129] ^ in[190]); 
    assign layer_0[3926] = in[90] | in[75]; 
    assign layer_0[3927] = in[59] & ~in[98]; 
    assign layer_0[3928] = in[184] & in[108]; 
    assign layer_0[3929] = in[242] & in[138]; 
    assign layer_0[3930] = in[67] & ~in[64]; 
    assign layer_0[3931] = in[110] ^ in[114]; 
    assign layer_0[3932] = in[26] | in[73]; 
    assign layer_0[3933] = ~in[143] | (in[36] & in[143]); 
    assign layer_0[3934] = ~in[118] | (in[118] & in[163]); 
    assign layer_0[3935] = ~in[182]; 
    assign layer_0[3936] = in[178] | in[104]; 
    assign layer_0[3937] = in[90] & in[173]; 
    assign layer_0[3938] = in[31] ^ in[20]; 
    assign layer_0[3939] = ~in[195] | (in[195] & in[219]); 
    assign layer_0[3940] = ~(in[194] | in[197]); 
    assign layer_0[3941] = in[139] ^ in[125]; 
    assign layer_0[3942] = ~(in[13] & in[46]); 
    assign layer_0[3943] = ~in[147]; 
    assign layer_0[3944] = ~in[163] | (in[109] & in[163]); 
    assign layer_0[3945] = ~in[228] | (in[170] & in[228]); 
    assign layer_0[3946] = in[121] | in[225]; 
    assign layer_0[3947] = in[43] | in[106]; 
    assign layer_0[3948] = in[137] & ~in[28]; 
    assign layer_0[3949] = ~(in[204] ^ in[145]); 
    assign layer_0[3950] = in[121] | in[197]; 
    assign layer_0[3951] = ~(in[124] | in[195]); 
    assign layer_0[3952] = in[145] | in[230]; 
    assign layer_0[3953] = in[211] & ~in[145]; 
    assign layer_0[3954] = ~(in[163] ^ in[137]); 
    assign layer_0[3955] = ~in[166] | (in[166] & in[156]); 
    assign layer_0[3956] = in[107] ^ in[82]; 
    assign layer_0[3957] = in[66] & ~in[111]; 
    assign layer_0[3958] = in[246] & ~in[247]; 
    assign layer_0[3959] = ~in[74] | (in[74] & in[2]); 
    assign layer_0[3960] = ~(in[241] | in[137]); 
    assign layer_0[3961] = in[213]; 
    assign layer_0[3962] = in[132] & ~in[226]; 
    assign layer_0[3963] = in[30] & in[158]; 
    assign layer_0[3964] = ~(in[87] ^ in[187]); 
    assign layer_0[3965] = in[61] ^ in[145]; 
    assign layer_0[3966] = in[254] | in[158]; 
    assign layer_0[3967] = in[91] ^ in[153]; 
    assign layer_0[3968] = ~in[3]; 
    assign layer_0[3969] = in[179]; 
    assign layer_0[3970] = ~(in[96] | in[182]); 
    assign layer_0[3971] = ~in[181] | (in[84] & in[181]); 
    assign layer_0[3972] = in[174] & in[240]; 
    assign layer_0[3973] = in[72] & ~in[24]; 
    assign layer_0[3974] = in[163] & ~in[141]; 
    assign layer_0[3975] = ~in[126] | (in[126] & in[237]); 
    assign layer_0[3976] = ~in[107]; 
    assign layer_0[3977] = ~in[93]; 
    assign layer_0[3978] = ~(in[61] ^ in[10]); 
    assign layer_0[3979] = in[163]; 
    assign layer_0[3980] = ~(in[238] & in[126]); 
    assign layer_0[3981] = ~in[224]; 
    assign layer_0[3982] = ~in[173]; 
    assign layer_0[3983] = ~(in[35] ^ in[37]); 
    assign layer_0[3984] = ~(in[139] ^ in[205]); 
    assign layer_0[3985] = ~in[211]; 
    assign layer_0[3986] = ~(in[193] ^ in[163]); 
    assign layer_0[3987] = ~in[174]; 
    assign layer_0[3988] = ~in[13] | (in[13] & in[95]); 
    assign layer_0[3989] = in[231]; 
    assign layer_0[3990] = ~in[150]; 
    assign layer_0[3991] = ~(in[196] ^ in[184]); 
    assign layer_0[3992] = in[41] | in[129]; 
    assign layer_0[3993] = ~in[189] | (in[189] & in[66]); 
    assign layer_0[3994] = in[129] & ~in[1]; 
    assign layer_0[3995] = in[157]; 
    assign layer_0[3996] = ~in[200]; 
    assign layer_0[3997] = in[95] | in[139]; 
    assign layer_0[3998] = in[59]; 
    assign layer_0[3999] = in[184] & in[175]; 
    // Layer 1 ============================================================
    assign layer_1[0] = layer_0[2944]; 
    assign layer_1[1] = ~(layer_0[3297] & layer_0[3176]); 
    assign layer_1[2] = layer_0[3837] & layer_0[3709]; 
    assign layer_1[3] = layer_0[2429] | layer_0[2506]; 
    assign layer_1[4] = layer_0[53] ^ layer_0[148]; 
    assign layer_1[5] = layer_0[793] & layer_0[792]; 
    assign layer_1[6] = ~layer_0[1331]; 
    assign layer_1[7] = ~layer_0[138] | (layer_0[138] & layer_0[208]); 
    assign layer_1[8] = ~(layer_0[3543] | layer_0[3468]); 
    assign layer_1[9] = layer_0[1345] ^ layer_0[1394]; 
    assign layer_1[10] = layer_0[1801]; 
    assign layer_1[11] = layer_0[2204] ^ layer_0[2298]; 
    assign layer_1[12] = layer_0[3081]; 
    assign layer_1[13] = ~layer_0[3326]; 
    assign layer_1[14] = ~(layer_0[3276] | layer_0[3262]); 
    assign layer_1[15] = ~layer_0[62] | (layer_0[62] & layer_0[17]); 
    assign layer_1[16] = ~layer_0[3787] | (layer_0[3788] & layer_0[3787]); 
    assign layer_1[17] = ~layer_0[779]; 
    assign layer_1[18] = layer_0[307]; 
    assign layer_1[19] = layer_0[2768] & layer_0[2751]; 
    assign layer_1[20] = ~layer_0[3407]; 
    assign layer_1[21] = layer_0[1478]; 
    assign layer_1[22] = ~(layer_0[3943] | layer_0[3874]); 
    assign layer_1[23] = ~layer_0[1360]; 
    assign layer_1[24] = ~layer_0[2662] | (layer_0[2662] & layer_0[2776]); 
    assign layer_1[25] = layer_0[3518] & ~layer_0[3527]; 
    assign layer_1[26] = layer_0[3248]; 
    assign layer_1[27] = layer_0[1168] ^ layer_0[1195]; 
    assign layer_1[28] = ~layer_0[3814]; 
    assign layer_1[29] = layer_0[3747] & ~layer_0[3621]; 
    assign layer_1[30] = layer_0[2394] & ~layer_0[2420]; 
    assign layer_1[31] = ~(layer_0[3726] | layer_0[3795]); 
    assign layer_1[32] = layer_0[3863] & layer_0[3978]; 
    assign layer_1[33] = ~layer_0[201]; 
    assign layer_1[34] = ~layer_0[335]; 
    assign layer_1[35] = ~layer_0[3856] | (layer_0[3849] & layer_0[3856]); 
    assign layer_1[36] = layer_0[592] & ~layer_0[505]; 
    assign layer_1[37] = ~layer_0[934] | (layer_0[1004] & layer_0[934]); 
    assign layer_1[38] = ~layer_0[584] | (layer_0[584] & layer_0[687]); 
    assign layer_1[39] = ~layer_0[1264] | (layer_0[1326] & layer_0[1264]); 
    assign layer_1[40] = ~layer_0[3867] | (layer_0[3867] & layer_0[3887]); 
    assign layer_1[41] = ~(layer_0[3966] ^ layer_0[3974]); 
    assign layer_1[42] = layer_0[1491] | layer_0[1427]; 
    assign layer_1[43] = ~(layer_0[3043] ^ layer_0[3095]); 
    assign layer_1[44] = layer_0[291] & ~layer_0[333]; 
    assign layer_1[45] = layer_0[3895]; 
    assign layer_1[46] = ~(layer_0[3083] & layer_0[3063]); 
    assign layer_1[47] = layer_0[804] ^ layer_0[716]; 
    assign layer_1[48] = ~layer_0[2949]; 
    assign layer_1[49] = layer_0[2009] & ~layer_0[2080]; 
    assign layer_1[50] = layer_0[1364]; 
    assign layer_1[51] = layer_0[1283]; 
    assign layer_1[52] = ~(layer_0[911] & layer_0[807]); 
    assign layer_1[53] = ~layer_0[2705] | (layer_0[2705] & layer_0[2617]); 
    assign layer_1[54] = ~layer_0[1428]; 
    assign layer_1[55] = layer_0[3948] & ~layer_0[3892]; 
    assign layer_1[56] = ~(layer_0[1440] ^ layer_0[1534]); 
    assign layer_1[57] = layer_0[3301] & layer_0[3398]; 
    assign layer_1[58] = ~(layer_0[1957] ^ layer_0[2022]); 
    assign layer_1[59] = layer_0[30]; 
    assign layer_1[60] = ~(layer_0[154] & layer_0[171]); 
    assign layer_1[61] = ~(layer_0[1451] ^ layer_0[1354]); 
    assign layer_1[62] = layer_0[2218]; 
    assign layer_1[63] = ~layer_0[700] | (layer_0[700] & layer_0[671]); 
    assign layer_1[64] = layer_0[3744] & layer_0[3700]; 
    assign layer_1[65] = layer_0[2313] & ~layer_0[2392]; 
    assign layer_1[66] = layer_0[3699]; 
    assign layer_1[67] = ~layer_0[1957] | (layer_0[1962] & layer_0[1957]); 
    assign layer_1[68] = layer_0[1411] & ~layer_0[1372]; 
    assign layer_1[69] = layer_0[1248] & ~layer_0[1172]; 
    assign layer_1[70] = ~layer_0[570]; 
    assign layer_1[71] = ~layer_0[2484] | (layer_0[2501] & layer_0[2484]); 
    assign layer_1[72] = ~(layer_0[2017] ^ layer_0[2062]); 
    assign layer_1[73] = layer_0[1928] & ~layer_0[1998]; 
    assign layer_1[74] = ~(layer_0[375] | layer_0[379]); 
    assign layer_1[75] = ~layer_0[1074] | (layer_0[1074] & layer_0[997]); 
    assign layer_1[76] = layer_0[1259] & ~layer_0[1155]; 
    assign layer_1[77] = ~(layer_0[3072] ^ layer_0[2976]); 
    assign layer_1[78] = ~layer_0[3674]; 
    assign layer_1[79] = layer_0[1151] & ~layer_0[1031]; 
    assign layer_1[80] = ~(layer_0[690] ^ layer_0[658]); 
    assign layer_1[81] = layer_0[1060] & ~layer_0[1033]; 
    assign layer_1[82] = layer_0[2565]; 
    assign layer_1[83] = layer_0[2672]; 
    assign layer_1[84] = ~layer_0[458]; 
    assign layer_1[85] = layer_0[496]; 
    assign layer_1[86] = ~layer_0[1519] | (layer_0[1519] & layer_0[1413]); 
    assign layer_1[87] = ~(layer_0[1140] | layer_0[1125]); 
    assign layer_1[88] = layer_0[1449]; 
    assign layer_1[89] = layer_0[2731] & ~layer_0[2653]; 
    assign layer_1[90] = ~layer_0[1833]; 
    assign layer_1[91] = layer_0[3647] & ~layer_0[3694]; 
    assign layer_1[92] = ~layer_0[911]; 
    assign layer_1[93] = ~layer_0[2357]; 
    assign layer_1[94] = layer_0[3839]; 
    assign layer_1[95] = layer_0[1241] ^ layer_0[1113]; 
    assign layer_1[96] = layer_0[2836] ^ layer_0[2714]; 
    assign layer_1[97] = ~layer_0[3964]; 
    assign layer_1[98] = ~layer_0[2582] | (layer_0[2582] & layer_0[2473]); 
    assign layer_1[99] = ~(layer_0[2537] & layer_0[2411]); 
    assign layer_1[100] = layer_0[3232]; 
    assign layer_1[101] = ~(layer_0[2104] ^ layer_0[2013]); 
    assign layer_1[102] = layer_0[1952] & ~layer_0[1994]; 
    assign layer_1[103] = layer_0[1919] & ~layer_0[1966]; 
    assign layer_1[104] = layer_0[2948] | layer_0[2851]; 
    assign layer_1[105] = ~(layer_0[3368] ^ layer_0[3477]); 
    assign layer_1[106] = layer_0[234] & layer_0[354]; 
    assign layer_1[107] = ~(layer_0[3385] | layer_0[3340]); 
    assign layer_1[108] = ~layer_0[3203] | (layer_0[3203] & layer_0[3138]); 
    assign layer_1[109] = layer_0[1968] ^ layer_0[1891]; 
    assign layer_1[110] = layer_0[3794] & layer_0[3837]; 
    assign layer_1[111] = layer_0[24]; 
    assign layer_1[112] = ~layer_0[1761]; 
    assign layer_1[113] = layer_0[2593]; 
    assign layer_1[114] = layer_0[1928] & layer_0[2051]; 
    assign layer_1[115] = layer_0[174]; 
    assign layer_1[116] = ~layer_0[632] | (layer_0[632] & layer_0[697]); 
    assign layer_1[117] = layer_0[1924]; 
    assign layer_1[118] = ~layer_0[3178]; 
    assign layer_1[119] = layer_0[3037]; 
    assign layer_1[120] = ~layer_0[2331]; 
    assign layer_1[121] = layer_0[1480]; 
    assign layer_1[122] = ~layer_0[1013] | (layer_0[1013] & layer_0[972]); 
    assign layer_1[123] = layer_0[3951] ^ layer_0[3914]; 
    assign layer_1[124] = ~(layer_0[3359] & layer_0[3406]); 
    assign layer_1[125] = ~(layer_0[1402] | layer_0[1420]); 
    assign layer_1[126] = layer_0[3275]; 
    assign layer_1[127] = ~(layer_0[1451] | layer_0[1513]); 
    assign layer_1[128] = ~layer_0[10]; 
    assign layer_1[129] = ~(layer_0[2277] & layer_0[2253]); 
    assign layer_1[130] = layer_0[3030] | layer_0[3092]; 
    assign layer_1[131] = ~(layer_0[3422] | layer_0[3356]); 
    assign layer_1[132] = layer_0[1686]; 
    assign layer_1[133] = layer_0[310]; 
    assign layer_1[134] = layer_0[3161]; 
    assign layer_1[135] = layer_0[1793] & ~layer_0[1702]; 
    assign layer_1[136] = layer_0[3524] & ~layer_0[3526]; 
    assign layer_1[137] = ~layer_0[193] | (layer_0[112] & layer_0[193]); 
    assign layer_1[138] = ~layer_0[2957]; 
    assign layer_1[139] = layer_0[3525] & ~layer_0[3613]; 
    assign layer_1[140] = ~layer_0[3355] | (layer_0[3355] & layer_0[3310]); 
    assign layer_1[141] = layer_0[3218] & layer_0[3207]; 
    assign layer_1[142] = ~layer_0[1985]; 
    assign layer_1[143] = ~layer_0[372] | (layer_0[484] & layer_0[372]); 
    assign layer_1[144] = ~layer_0[1097] | (layer_0[1097] & layer_0[1174]); 
    assign layer_1[145] = layer_0[259]; 
    assign layer_1[146] = ~(layer_0[1556] | layer_0[1621]); 
    assign layer_1[147] = ~(layer_0[1627] & layer_0[1634]); 
    assign layer_1[148] = ~(layer_0[3472] | layer_0[3559]); 
    assign layer_1[149] = layer_0[3241] ^ layer_0[3368]; 
    assign layer_1[150] = layer_0[1354] & ~layer_0[1233]; 
    assign layer_1[151] = ~layer_0[3510] | (layer_0[3465] & layer_0[3510]); 
    assign layer_1[152] = ~layer_0[3353] | (layer_0[3353] & layer_0[3323]); 
    assign layer_1[153] = layer_0[2473] ^ layer_0[2492]; 
    assign layer_1[154] = ~(layer_0[2361] | layer_0[2479]); 
    assign layer_1[155] = layer_0[3309]; 
    assign layer_1[156] = ~layer_0[1824] | (layer_0[1824] & layer_0[1826]); 
    assign layer_1[157] = ~layer_0[2132] | (layer_0[2154] & layer_0[2132]); 
    assign layer_1[158] = layer_0[2588]; 
    assign layer_1[159] = ~layer_0[257] | (layer_0[257] & layer_0[323]); 
    assign layer_1[160] = ~(layer_0[1820] & layer_0[1874]); 
    assign layer_1[161] = layer_0[2509]; 
    assign layer_1[162] = ~layer_0[1599] | (layer_0[1599] & layer_0[1555]); 
    assign layer_1[163] = ~(layer_0[3067] & layer_0[3105]); 
    assign layer_1[164] = layer_0[3471]; 
    assign layer_1[165] = ~layer_0[2231]; 
    assign layer_1[166] = ~(layer_0[46] ^ layer_0[95]); 
    assign layer_1[167] = layer_0[2491] & ~layer_0[2499]; 
    assign layer_1[168] = layer_0[1271] ^ layer_0[1335]; 
    assign layer_1[169] = ~(layer_0[3254] ^ layer_0[3263]); 
    assign layer_1[170] = layer_0[3383] | layer_0[3370]; 
    assign layer_1[171] = layer_0[2328] & ~layer_0[2356]; 
    assign layer_1[172] = layer_0[1919] | layer_0[1791]; 
    assign layer_1[173] = layer_0[3124]; 
    assign layer_1[174] = layer_0[2630]; 
    assign layer_1[175] = ~(layer_0[3270] | layer_0[3149]); 
    assign layer_1[176] = layer_0[2417] ^ layer_0[2462]; 
    assign layer_1[177] = layer_0[1396] & ~layer_0[1291]; 
    assign layer_1[178] = ~layer_0[859]; 
    assign layer_1[179] = layer_0[51]; 
    assign layer_1[180] = ~layer_0[1535] | (layer_0[1535] & layer_0[1510]); 
    assign layer_1[181] = ~layer_0[1065] | (layer_0[1065] & layer_0[1153]); 
    assign layer_1[182] = ~(layer_0[2962] | layer_0[2885]); 
    assign layer_1[183] = layer_0[3561]; 
    assign layer_1[184] = layer_0[3974] & layer_0[3847]; 
    assign layer_1[185] = ~(layer_0[2976] | layer_0[2984]); 
    assign layer_1[186] = ~layer_0[2152] | (layer_0[2152] & layer_0[2134]); 
    assign layer_1[187] = ~(layer_0[2616] & layer_0[2723]); 
    assign layer_1[188] = ~layer_0[1169]; 
    assign layer_1[189] = layer_0[1549] & ~layer_0[1676]; 
    assign layer_1[190] = layer_0[3145] & ~layer_0[3106]; 
    assign layer_1[191] = ~(layer_0[1586] ^ layer_0[1649]); 
    assign layer_1[192] = ~layer_0[3381]; 
    assign layer_1[193] = layer_0[3334]; 
    assign layer_1[194] = ~layer_0[2212] | (layer_0[2307] & layer_0[2212]); 
    assign layer_1[195] = layer_0[1633]; 
    assign layer_1[196] = layer_0[2685] ^ layer_0[2783]; 
    assign layer_1[197] = layer_0[3723] | layer_0[3622]; 
    assign layer_1[198] = ~layer_0[3998] | (layer_0[3998] & layer_0[3971]); 
    assign layer_1[199] = layer_0[292] | layer_0[306]; 
    assign layer_1[200] = layer_0[236] ^ layer_0[287]; 
    assign layer_1[201] = layer_0[3419]; 
    assign layer_1[202] = ~layer_0[3117]; 
    assign layer_1[203] = layer_0[469]; 
    assign layer_1[204] = ~layer_0[965]; 
    assign layer_1[205] = layer_0[1197] & ~layer_0[1319]; 
    assign layer_1[206] = ~layer_0[1576] | (layer_0[1631] & layer_0[1576]); 
    assign layer_1[207] = layer_0[3320]; 
    assign layer_1[208] = ~layer_0[2341]; 
    assign layer_1[209] = ~(layer_0[381] ^ layer_0[428]); 
    assign layer_1[210] = ~layer_0[495] | (layer_0[495] & layer_0[478]); 
    assign layer_1[211] = ~layer_0[3787] | (layer_0[3735] & layer_0[3787]); 
    assign layer_1[212] = ~(layer_0[1960] | layer_0[2042]); 
    assign layer_1[213] = ~layer_0[2531]; 
    assign layer_1[214] = ~(layer_0[3754] & layer_0[3671]); 
    assign layer_1[215] = layer_0[549] & ~layer_0[553]; 
    assign layer_1[216] = layer_0[915] & ~layer_0[983]; 
    assign layer_1[217] = ~(layer_0[673] & layer_0[555]); 
    assign layer_1[218] = layer_0[1622] & ~layer_0[1630]; 
    assign layer_1[219] = ~layer_0[3254]; 
    assign layer_1[220] = ~(layer_0[2493] ^ layer_0[2537]); 
    assign layer_1[221] = ~(layer_0[181] & layer_0[201]); 
    assign layer_1[222] = ~layer_0[1817] | (layer_0[1817] & layer_0[1772]); 
    assign layer_1[223] = layer_0[1392] & ~layer_0[1504]; 
    assign layer_1[224] = ~layer_0[2816] | (layer_0[2711] & layer_0[2816]); 
    assign layer_1[225] = ~layer_0[1946] | (layer_0[1840] & layer_0[1946]); 
    assign layer_1[226] = layer_0[1127] & ~layer_0[1011]; 
    assign layer_1[227] = layer_0[1039]; 
    assign layer_1[228] = layer_0[3458] & ~layer_0[3344]; 
    assign layer_1[229] = layer_0[3817] & ~layer_0[3842]; 
    assign layer_1[230] = ~layer_0[1367]; 
    assign layer_1[231] = ~layer_0[2493]; 
    assign layer_1[232] = ~(layer_0[2309] & layer_0[2223]); 
    assign layer_1[233] = layer_0[933] & layer_0[1058]; 
    assign layer_1[234] = layer_0[2323] & ~layer_0[2230]; 
    assign layer_1[235] = layer_0[2085] | layer_0[2027]; 
    assign layer_1[236] = layer_0[2431] & layer_0[2322]; 
    assign layer_1[237] = ~(layer_0[1855] & layer_0[1885]); 
    assign layer_1[238] = layer_0[64] & ~layer_0[132]; 
    assign layer_1[239] = ~layer_0[1597] | (layer_0[1597] & layer_0[1482]); 
    assign layer_1[240] = ~(layer_0[2726] & layer_0[2809]); 
    assign layer_1[241] = layer_0[3644] & ~layer_0[3634]; 
    assign layer_1[242] = ~layer_0[524]; 
    assign layer_1[243] = ~(layer_0[2766] | layer_0[2734]); 
    assign layer_1[244] = layer_0[3264]; 
    assign layer_1[245] = ~(layer_0[3780] | layer_0[3742]); 
    assign layer_1[246] = ~layer_0[3102] | (layer_0[3102] & layer_0[3016]); 
    assign layer_1[247] = ~layer_0[296]; 
    assign layer_1[248] = layer_0[507] & ~layer_0[565]; 
    assign layer_1[249] = layer_0[3587] & layer_0[3632]; 
    assign layer_1[250] = layer_0[667] & ~layer_0[760]; 
    assign layer_1[251] = layer_0[605]; 
    assign layer_1[252] = layer_0[1580] & ~layer_0[1463]; 
    assign layer_1[253] = layer_0[1082]; 
    assign layer_1[254] = layer_0[2539] & layer_0[2507]; 
    assign layer_1[255] = layer_0[2500] & layer_0[2605]; 
    assign layer_1[256] = ~(layer_0[366] ^ layer_0[386]); 
    assign layer_1[257] = ~layer_0[231] | (layer_0[231] & layer_0[190]); 
    assign layer_1[258] = layer_0[3678] & ~layer_0[3689]; 
    assign layer_1[259] = layer_0[1203]; 
    assign layer_1[260] = ~(layer_0[2067] & layer_0[2129]); 
    assign layer_1[261] = layer_0[3150]; 
    assign layer_1[262] = ~layer_0[3532]; 
    assign layer_1[263] = layer_0[3707] | layer_0[3610]; 
    assign layer_1[264] = layer_0[3008] ^ layer_0[2898]; 
    assign layer_1[265] = ~layer_0[819]; 
    assign layer_1[266] = layer_0[3219] & layer_0[3342]; 
    assign layer_1[267] = layer_0[1944] & ~layer_0[1979]; 
    assign layer_1[268] = layer_0[602]; 
    assign layer_1[269] = ~(layer_0[865] & layer_0[934]); 
    assign layer_1[270] = ~layer_0[2705]; 
    assign layer_1[271] = ~layer_0[1727]; 
    assign layer_1[272] = ~(layer_0[2071] ^ layer_0[2133]); 
    assign layer_1[273] = layer_0[2114] & ~layer_0[2219]; 
    assign layer_1[274] = ~(layer_0[843] & layer_0[729]); 
    assign layer_1[275] = ~layer_0[1703] | (layer_0[1675] & layer_0[1703]); 
    assign layer_1[276] = ~layer_0[3558]; 
    assign layer_1[277] = ~layer_0[1486]; 
    assign layer_1[278] = ~layer_0[541]; 
    assign layer_1[279] = ~layer_0[437]; 
    assign layer_1[280] = layer_0[1337] & ~layer_0[1328]; 
    assign layer_1[281] = ~(layer_0[3351] | layer_0[3449]); 
    assign layer_1[282] = ~layer_0[2571]; 
    assign layer_1[283] = ~layer_0[256] | (layer_0[256] & layer_0[358]); 
    assign layer_1[284] = layer_0[2734]; 
    assign layer_1[285] = layer_0[196]; 
    assign layer_1[286] = layer_0[2937] & ~layer_0[2822]; 
    assign layer_1[287] = ~layer_0[1827]; 
    assign layer_1[288] = ~(layer_0[3765] | layer_0[3777]); 
    assign layer_1[289] = ~layer_0[3286]; 
    assign layer_1[290] = ~(layer_0[2226] & layer_0[2202]); 
    assign layer_1[291] = layer_0[3848] | layer_0[3871]; 
    assign layer_1[292] = ~(layer_0[2267] ^ layer_0[2394]); 
    assign layer_1[293] = layer_0[1778]; 
    assign layer_1[294] = ~(layer_0[3574] & layer_0[3679]); 
    assign layer_1[295] = ~layer_0[3681] | (layer_0[3638] & layer_0[3681]); 
    assign layer_1[296] = ~layer_0[221]; 
    assign layer_1[297] = ~layer_0[1953] | (layer_0[2058] & layer_0[1953]); 
    assign layer_1[298] = layer_0[2102]; 
    assign layer_1[299] = layer_0[2193] ^ layer_0[2278]; 
    assign layer_1[300] = ~layer_0[1390] | (layer_0[1390] & layer_0[1388]); 
    assign layer_1[301] = ~(layer_0[1980] & layer_0[1961]); 
    assign layer_1[302] = ~(layer_0[3039] ^ layer_0[3098]); 
    assign layer_1[303] = ~(layer_0[506] & layer_0[574]); 
    assign layer_1[304] = ~layer_0[3694] | (layer_0[3611] & layer_0[3694]); 
    assign layer_1[305] = ~layer_0[3226]; 
    assign layer_1[306] = ~layer_0[1721]; 
    assign layer_1[307] = layer_0[3017] & ~layer_0[3094]; 
    assign layer_1[308] = layer_0[31] | layer_0[38]; 
    assign layer_1[309] = layer_0[2754] & layer_0[2778]; 
    assign layer_1[310] = ~layer_0[1048]; 
    assign layer_1[311] = ~layer_0[3895] | (layer_0[3895] & layer_0[3923]); 
    assign layer_1[312] = layer_0[2611] ^ layer_0[2653]; 
    assign layer_1[313] = ~(layer_0[27] & layer_0[39]); 
    assign layer_1[314] = ~layer_0[527] | (layer_0[615] & layer_0[527]); 
    assign layer_1[315] = layer_0[3833] & layer_0[3950]; 
    assign layer_1[316] = layer_0[1016] & ~layer_0[1118]; 
    assign layer_1[317] = ~layer_0[94] | (layer_0[94] & layer_0[33]); 
    assign layer_1[318] = layer_0[2328] & layer_0[2388]; 
    assign layer_1[319] = layer_0[3874] ^ layer_0[3809]; 
    assign layer_1[320] = ~layer_0[3147]; 
    assign layer_1[321] = layer_0[306] ^ layer_0[410]; 
    assign layer_1[322] = layer_0[3800]; 
    assign layer_1[323] = ~(layer_0[855] | layer_0[929]); 
    assign layer_1[324] = layer_0[3248] ^ layer_0[3137]; 
    assign layer_1[325] = ~(layer_0[1842] ^ layer_0[1843]); 
    assign layer_1[326] = layer_0[1967]; 
    assign layer_1[327] = ~(layer_0[191] | layer_0[188]); 
    assign layer_1[328] = layer_0[2658] | layer_0[2774]; 
    assign layer_1[329] = ~(layer_0[3243] | layer_0[3343]); 
    assign layer_1[330] = layer_0[172]; 
    assign layer_1[331] = ~layer_0[1183] | (layer_0[1310] & layer_0[1183]); 
    assign layer_1[332] = layer_0[704]; 
    assign layer_1[333] = ~layer_0[413]; 
    assign layer_1[334] = ~(layer_0[2980] | layer_0[2863]); 
    assign layer_1[335] = layer_0[2843] & ~layer_0[2739]; 
    assign layer_1[336] = layer_0[2260] & ~layer_0[2308]; 
    assign layer_1[337] = layer_0[1316] & layer_0[1427]; 
    assign layer_1[338] = layer_0[2225] & ~layer_0[2255]; 
    assign layer_1[339] = ~(layer_0[3394] & layer_0[3275]); 
    assign layer_1[340] = layer_0[1505]; 
    assign layer_1[341] = ~layer_0[3962]; 
    assign layer_1[342] = layer_0[612]; 
    assign layer_1[343] = ~layer_0[1033]; 
    assign layer_1[344] = layer_0[58]; 
    assign layer_1[345] = ~layer_0[643]; 
    assign layer_1[346] = layer_0[1330]; 
    assign layer_1[347] = layer_0[1181]; 
    assign layer_1[348] = layer_0[3467] & ~layer_0[3534]; 
    assign layer_1[349] = ~(layer_0[3734] ^ layer_0[3801]); 
    assign layer_1[350] = ~layer_0[730] | (layer_0[699] & layer_0[730]); 
    assign layer_1[351] = ~layer_0[2810] | (layer_0[2734] & layer_0[2810]); 
    assign layer_1[352] = layer_0[2499]; 
    assign layer_1[353] = layer_0[907]; 
    assign layer_1[354] = layer_0[407] & ~layer_0[302]; 
    assign layer_1[355] = ~(layer_0[2463] ^ layer_0[2409]); 
    assign layer_1[356] = ~layer_0[2125]; 
    assign layer_1[357] = layer_0[3394] | layer_0[3445]; 
    assign layer_1[358] = layer_0[2772] ^ layer_0[2725]; 
    assign layer_1[359] = ~layer_0[697]; 
    assign layer_1[360] = layer_0[1524] & layer_0[1484]; 
    assign layer_1[361] = ~layer_0[1423] | (layer_0[1334] & layer_0[1423]); 
    assign layer_1[362] = layer_0[2037]; 
    assign layer_1[363] = ~(layer_0[2120] ^ layer_0[2122]); 
    assign layer_1[364] = layer_0[3581] | layer_0[3502]; 
    assign layer_1[365] = layer_0[2407]; 
    assign layer_1[366] = ~layer_0[3631] | (layer_0[3539] & layer_0[3631]); 
    assign layer_1[367] = ~(layer_0[2483] | layer_0[2371]); 
    assign layer_1[368] = layer_0[577]; 
    assign layer_1[369] = layer_0[3132] ^ layer_0[3104]; 
    assign layer_1[370] = layer_0[2905]; 
    assign layer_1[371] = ~(layer_0[2059] ^ layer_0[1995]); 
    assign layer_1[372] = layer_0[2922] & ~layer_0[2863]; 
    assign layer_1[373] = layer_0[1622]; 
    assign layer_1[374] = layer_0[2237]; 
    assign layer_1[375] = layer_0[3262] & ~layer_0[3321]; 
    assign layer_1[376] = ~(layer_0[2216] | layer_0[2126]); 
    assign layer_1[377] = layer_0[536] | layer_0[439]; 
    assign layer_1[378] = ~(layer_0[593] | layer_0[506]); 
    assign layer_1[379] = layer_0[2460]; 
    assign layer_1[380] = ~layer_0[883] | (layer_0[932] & layer_0[883]); 
    assign layer_1[381] = ~layer_0[2413]; 
    assign layer_1[382] = layer_0[3849]; 
    assign layer_1[383] = layer_0[1328] | layer_0[1392]; 
    assign layer_1[384] = layer_0[2800]; 
    assign layer_1[385] = layer_0[2981] & ~layer_0[3001]; 
    assign layer_1[386] = layer_0[2201] & ~layer_0[2239]; 
    assign layer_1[387] = layer_0[3814] & ~layer_0[3695]; 
    assign layer_1[388] = ~layer_0[1669] | (layer_0[1767] & layer_0[1669]); 
    assign layer_1[389] = layer_0[3072]; 
    assign layer_1[390] = layer_0[3859] | layer_0[3957]; 
    assign layer_1[391] = layer_0[1427]; 
    assign layer_1[392] = ~layer_0[930]; 
    assign layer_1[393] = layer_0[1123]; 
    assign layer_1[394] = ~(layer_0[2368] & layer_0[2272]); 
    assign layer_1[395] = layer_0[1533] ^ layer_0[1522]; 
    assign layer_1[396] = layer_0[2753] ^ layer_0[2656]; 
    assign layer_1[397] = ~(layer_0[187] ^ layer_0[268]); 
    assign layer_1[398] = layer_0[434]; 
    assign layer_1[399] = ~layer_0[1569]; 
    assign layer_1[400] = layer_0[1072] & ~layer_0[1058]; 
    assign layer_1[401] = layer_0[2563] & ~layer_0[2685]; 
    assign layer_1[402] = ~layer_0[2916] | (layer_0[2806] & layer_0[2916]); 
    assign layer_1[403] = ~(layer_0[28] ^ layer_0[151]); 
    assign layer_1[404] = ~layer_0[1996]; 
    assign layer_1[405] = ~(layer_0[2810] ^ layer_0[2704]); 
    assign layer_1[406] = layer_0[875]; 
    assign layer_1[407] = layer_0[139] & ~layer_0[80]; 
    assign layer_1[408] = layer_0[3478] & ~layer_0[3517]; 
    assign layer_1[409] = ~layer_0[3529] | (layer_0[3529] & layer_0[3603]); 
    assign layer_1[410] = layer_0[3751] | layer_0[3836]; 
    assign layer_1[411] = ~layer_0[3722]; 
    assign layer_1[412] = ~layer_0[3614] | (layer_0[3528] & layer_0[3614]); 
    assign layer_1[413] = ~layer_0[960] | (layer_0[1007] & layer_0[960]); 
    assign layer_1[414] = layer_0[2197] ^ layer_0[2316]; 
    assign layer_1[415] = ~layer_0[2516]; 
    assign layer_1[416] = layer_0[3850]; 
    assign layer_1[417] = ~layer_0[1254]; 
    assign layer_1[418] = ~(layer_0[3997] | layer_0[3877]); 
    assign layer_1[419] = ~layer_0[172]; 
    assign layer_1[420] = layer_0[2432]; 
    assign layer_1[421] = ~(layer_0[1119] & layer_0[1137]); 
    assign layer_1[422] = ~(layer_0[791] | layer_0[887]); 
    assign layer_1[423] = ~(layer_0[3025] & layer_0[3152]); 
    assign layer_1[424] = layer_0[2935]; 
    assign layer_1[425] = layer_0[1382] & ~layer_0[1417]; 
    assign layer_1[426] = layer_0[1409] & layer_0[1357]; 
    assign layer_1[427] = ~(layer_0[450] & layer_0[404]); 
    assign layer_1[428] = ~(layer_0[729] & layer_0[746]); 
    assign layer_1[429] = ~(layer_0[3197] ^ layer_0[3152]); 
    assign layer_1[430] = ~layer_0[660] | (layer_0[660] & layer_0[754]); 
    assign layer_1[431] = layer_0[2856]; 
    assign layer_1[432] = ~(layer_0[1413] | layer_0[1451]); 
    assign layer_1[433] = ~layer_0[1720]; 
    assign layer_1[434] = ~layer_0[1256] | (layer_0[1342] & layer_0[1256]); 
    assign layer_1[435] = layer_0[3010]; 
    assign layer_1[436] = layer_0[2408]; 
    assign layer_1[437] = layer_0[733]; 
    assign layer_1[438] = ~layer_0[1155]; 
    assign layer_1[439] = layer_0[412]; 
    assign layer_1[440] = ~layer_0[1061] | (layer_0[1149] & layer_0[1061]); 
    assign layer_1[441] = layer_0[2093] & layer_0[2169]; 
    assign layer_1[442] = ~layer_0[3287]; 
    assign layer_1[443] = ~(layer_0[284] ^ layer_0[159]); 
    assign layer_1[444] = ~layer_0[3638]; 
    assign layer_1[445] = layer_0[1753] | layer_0[1829]; 
    assign layer_1[446] = layer_0[3823]; 
    assign layer_1[447] = ~layer_0[1105] | (layer_0[1076] & layer_0[1105]); 
    assign layer_1[448] = layer_0[1876] & ~layer_0[1960]; 
    assign layer_1[449] = layer_0[1191] ^ layer_0[1270]; 
    assign layer_1[450] = layer_0[3277]; 
    assign layer_1[451] = ~(layer_0[115] | layer_0[84]); 
    assign layer_1[452] = ~layer_0[501]; 
    assign layer_1[453] = ~(layer_0[2230] | layer_0[2145]); 
    assign layer_1[454] = ~layer_0[3280] | (layer_0[3280] & layer_0[3211]); 
    assign layer_1[455] = layer_0[3431]; 
    assign layer_1[456] = ~(layer_0[2131] & layer_0[2157]); 
    assign layer_1[457] = layer_0[2150] ^ layer_0[2029]; 
    assign layer_1[458] = layer_0[1465]; 
    assign layer_1[459] = ~(layer_0[2187] | layer_0[2280]); 
    assign layer_1[460] = ~layer_0[2082]; 
    assign layer_1[461] = ~(layer_0[972] ^ layer_0[984]); 
    assign layer_1[462] = ~layer_0[1167] | (layer_0[1167] & layer_0[1252]); 
    assign layer_1[463] = ~layer_0[202] | (layer_0[202] & layer_0[313]); 
    assign layer_1[464] = ~(layer_0[2805] ^ layer_0[2711]); 
    assign layer_1[465] = layer_0[3016]; 
    assign layer_1[466] = ~layer_0[474]; 
    assign layer_1[467] = ~layer_0[3303]; 
    assign layer_1[468] = ~(layer_0[3242] | layer_0[3349]); 
    assign layer_1[469] = ~(layer_0[1763] ^ layer_0[1771]); 
    assign layer_1[470] = layer_0[2288] & layer_0[2328]; 
    assign layer_1[471] = layer_0[92] | layer_0[12]; 
    assign layer_1[472] = ~layer_0[563] | (layer_0[487] & layer_0[563]); 
    assign layer_1[473] = ~layer_0[1840]; 
    assign layer_1[474] = layer_0[2062] & ~layer_0[2104]; 
    assign layer_1[475] = layer_0[3654]; 
    assign layer_1[476] = layer_0[716] ^ layer_0[795]; 
    assign layer_1[477] = layer_0[806] ^ layer_0[869]; 
    assign layer_1[478] = ~layer_0[2440]; 
    assign layer_1[479] = ~layer_0[3259] | (layer_0[3237] & layer_0[3259]); 
    assign layer_1[480] = layer_0[1293] & ~layer_0[1306]; 
    assign layer_1[481] = ~(layer_0[1452] | layer_0[1568]); 
    assign layer_1[482] = layer_0[3778] & ~layer_0[3765]; 
    assign layer_1[483] = layer_0[422]; 
    assign layer_1[484] = layer_0[3071]; 
    assign layer_1[485] = ~(layer_0[2652] ^ layer_0[2598]); 
    assign layer_1[486] = layer_0[3555] & layer_0[3581]; 
    assign layer_1[487] = layer_0[1614] & ~layer_0[1502]; 
    assign layer_1[488] = layer_0[2731] & ~layer_0[2763]; 
    assign layer_1[489] = layer_0[722] & ~layer_0[595]; 
    assign layer_1[490] = layer_0[3444] ^ layer_0[3418]; 
    assign layer_1[491] = ~(layer_0[3129] | layer_0[3071]); 
    assign layer_1[492] = ~layer_0[2119]; 
    assign layer_1[493] = ~(layer_0[3242] & layer_0[3258]); 
    assign layer_1[494] = ~layer_0[749]; 
    assign layer_1[495] = layer_0[2234] & ~layer_0[2313]; 
    assign layer_1[496] = ~(layer_0[2774] | layer_0[2816]); 
    assign layer_1[497] = layer_0[556] & layer_0[635]; 
    assign layer_1[498] = ~(layer_0[1035] | layer_0[913]); 
    assign layer_1[499] = ~layer_0[2160]; 
    assign layer_1[500] = ~layer_0[3495]; 
    assign layer_1[501] = ~(layer_0[922] & layer_0[940]); 
    assign layer_1[502] = layer_0[3560] & ~layer_0[3475]; 
    assign layer_1[503] = ~layer_0[3267] | (layer_0[3267] & layer_0[3191]); 
    assign layer_1[504] = ~layer_0[1362]; 
    assign layer_1[505] = ~(layer_0[2962] & layer_0[3036]); 
    assign layer_1[506] = ~(layer_0[974] ^ layer_0[855]); 
    assign layer_1[507] = layer_0[791]; 
    assign layer_1[508] = layer_0[1504] & ~layer_0[1596]; 
    assign layer_1[509] = layer_0[2475] ^ layer_0[2356]; 
    assign layer_1[510] = layer_0[2082]; 
    assign layer_1[511] = ~layer_0[2455]; 
    assign layer_1[512] = layer_0[3301] | layer_0[3303]; 
    assign layer_1[513] = layer_0[2684] & layer_0[2670]; 
    assign layer_1[514] = layer_0[235] ^ layer_0[342]; 
    assign layer_1[515] = layer_0[365]; 
    assign layer_1[516] = ~layer_0[190]; 
    assign layer_1[517] = layer_0[396] & layer_0[477]; 
    assign layer_1[518] = layer_0[2531]; 
    assign layer_1[519] = layer_0[702] & ~layer_0[689]; 
    assign layer_1[520] = ~layer_0[2795]; 
    assign layer_1[521] = ~(layer_0[3982] | layer_0[3994]); 
    assign layer_1[522] = ~layer_0[2971]; 
    assign layer_1[523] = ~(layer_0[2699] ^ layer_0[2607]); 
    assign layer_1[524] = ~layer_0[1384]; 
    assign layer_1[525] = layer_0[1382]; 
    assign layer_1[526] = layer_0[1639]; 
    assign layer_1[527] = ~layer_0[2859] | (layer_0[2859] & layer_0[2968]); 
    assign layer_1[528] = layer_0[57] ^ layer_0[51]; 
    assign layer_1[529] = ~layer_0[636]; 
    assign layer_1[530] = ~layer_0[3436]; 
    assign layer_1[531] = ~layer_0[3608]; 
    assign layer_1[532] = layer_0[38] | layer_0[45]; 
    assign layer_1[533] = ~layer_0[389]; 
    assign layer_1[534] = layer_0[1370] | layer_0[1327]; 
    assign layer_1[535] = ~(layer_0[105] | layer_0[73]); 
    assign layer_1[536] = ~(layer_0[951] & layer_0[943]); 
    assign layer_1[537] = ~layer_0[602] | (layer_0[602] & layer_0[671]); 
    assign layer_1[538] = ~(layer_0[3256] ^ layer_0[3167]); 
    assign layer_1[539] = ~layer_0[1702]; 
    assign layer_1[540] = ~layer_0[398]; 
    assign layer_1[541] = layer_0[3925] & ~layer_0[3926]; 
    assign layer_1[542] = layer_0[956]; 
    assign layer_1[543] = layer_0[2295] ^ layer_0[2269]; 
    assign layer_1[544] = ~layer_0[1959]; 
    assign layer_1[545] = layer_0[1754]; 
    assign layer_1[546] = ~(layer_0[689] | layer_0[805]); 
    assign layer_1[547] = ~layer_0[2145] | (layer_0[2047] & layer_0[2145]); 
    assign layer_1[548] = layer_0[2253] ^ layer_0[2229]; 
    assign layer_1[549] = layer_0[2371] ^ layer_0[2335]; 
    assign layer_1[550] = ~(layer_0[1390] ^ layer_0[1417]); 
    assign layer_1[551] = layer_0[2375]; 
    assign layer_1[552] = ~layer_0[3970]; 
    assign layer_1[553] = ~(layer_0[1918] | layer_0[1969]); 
    assign layer_1[554] = ~layer_0[2297] | (layer_0[2297] & layer_0[2310]); 
    assign layer_1[555] = layer_0[3825] & layer_0[3765]; 
    assign layer_1[556] = ~layer_0[3294]; 
    assign layer_1[557] = layer_0[1494]; 
    assign layer_1[558] = ~layer_0[2332] | (layer_0[2332] & layer_0[2314]); 
    assign layer_1[559] = layer_0[574] | layer_0[615]; 
    assign layer_1[560] = layer_0[3547] | layer_0[3448]; 
    assign layer_1[561] = layer_0[783]; 
    assign layer_1[562] = ~(layer_0[758] | layer_0[735]); 
    assign layer_1[563] = layer_0[1956] & ~layer_0[1970]; 
    assign layer_1[564] = layer_0[2142]; 
    assign layer_1[565] = layer_0[3393] & layer_0[3289]; 
    assign layer_1[566] = layer_0[621] ^ layer_0[723]; 
    assign layer_1[567] = layer_0[2584] | layer_0[2618]; 
    assign layer_1[568] = ~(layer_0[1229] ^ layer_0[1173]); 
    assign layer_1[569] = ~(layer_0[2348] & layer_0[2448]); 
    assign layer_1[570] = layer_0[2105]; 
    assign layer_1[571] = ~layer_0[3265] | (layer_0[3220] & layer_0[3265]); 
    assign layer_1[572] = ~(layer_0[491] | layer_0[426]); 
    assign layer_1[573] = ~layer_0[3568]; 
    assign layer_1[574] = ~layer_0[2487]; 
    assign layer_1[575] = ~(layer_0[2280] ^ layer_0[2186]); 
    assign layer_1[576] = ~(layer_0[2394] & layer_0[2507]); 
    assign layer_1[577] = layer_0[2288] ^ layer_0[2187]; 
    assign layer_1[578] = layer_0[1331] ^ layer_0[1405]; 
    assign layer_1[579] = layer_0[51] & layer_0[40]; 
    assign layer_1[580] = ~layer_0[3807]; 
    assign layer_1[581] = ~(layer_0[3431] | layer_0[3360]); 
    assign layer_1[582] = ~(layer_0[2083] ^ layer_0[2147]); 
    assign layer_1[583] = ~(layer_0[3037] & layer_0[3075]); 
    assign layer_1[584] = ~layer_0[3836]; 
    assign layer_1[585] = ~layer_0[2836]; 
    assign layer_1[586] = layer_0[885] & layer_0[827]; 
    assign layer_1[587] = ~(layer_0[614] ^ layer_0[726]); 
    assign layer_1[588] = layer_0[1201] | layer_0[1301]; 
    assign layer_1[589] = layer_0[3595] | layer_0[3646]; 
    assign layer_1[590] = ~layer_0[3928]; 
    assign layer_1[591] = layer_0[3368] & layer_0[3346]; 
    assign layer_1[592] = ~(layer_0[1223] ^ layer_0[1230]); 
    assign layer_1[593] = ~(layer_0[1315] ^ layer_0[1433]); 
    assign layer_1[594] = layer_0[1044] & layer_0[1011]; 
    assign layer_1[595] = ~(layer_0[3851] ^ layer_0[3923]); 
    assign layer_1[596] = ~layer_0[3873]; 
    assign layer_1[597] = layer_0[318] & layer_0[415]; 
    assign layer_1[598] = ~layer_0[3701]; 
    assign layer_1[599] = layer_0[1072]; 
    assign layer_1[600] = ~(layer_0[3989] | layer_0[3905]); 
    assign layer_1[601] = ~(layer_0[1847] ^ layer_0[1839]); 
    assign layer_1[602] = layer_0[2364]; 
    assign layer_1[603] = ~layer_0[166] | (layer_0[95] & layer_0[166]); 
    assign layer_1[604] = ~(layer_0[2821] ^ layer_0[2813]); 
    assign layer_1[605] = ~(layer_0[3309] | layer_0[3194]); 
    assign layer_1[606] = ~(layer_0[3644] & layer_0[3585]); 
    assign layer_1[607] = ~layer_0[1922]; 
    assign layer_1[608] = ~layer_0[93]; 
    assign layer_1[609] = layer_0[3802]; 
    assign layer_1[610] = layer_0[1192]; 
    assign layer_1[611] = layer_0[2805] & layer_0[2819]; 
    assign layer_1[612] = ~(layer_0[2758] | layer_0[2783]); 
    assign layer_1[613] = layer_0[1839]; 
    assign layer_1[614] = ~layer_0[1664]; 
    assign layer_1[615] = ~layer_0[2609]; 
    assign layer_1[616] = ~layer_0[3788]; 
    assign layer_1[617] = ~layer_0[1351] | (layer_0[1318] & layer_0[1351]); 
    assign layer_1[618] = layer_0[433]; 
    assign layer_1[619] = ~layer_0[3964]; 
    assign layer_1[620] = layer_0[3608]; 
    assign layer_1[621] = ~layer_0[1669]; 
    assign layer_1[622] = layer_0[1980] & ~layer_0[2053]; 
    assign layer_1[623] = ~layer_0[3874]; 
    assign layer_1[624] = layer_0[1589] | layer_0[1610]; 
    assign layer_1[625] = layer_0[1423] & ~layer_0[1434]; 
    assign layer_1[626] = ~layer_0[1320]; 
    assign layer_1[627] = ~(layer_0[3788] & layer_0[3763]); 
    assign layer_1[628] = ~(layer_0[671] & layer_0[552]); 
    assign layer_1[629] = layer_0[3233] & layer_0[3308]; 
    assign layer_1[630] = layer_0[427] ^ layer_0[367]; 
    assign layer_1[631] = ~(layer_0[3225] | layer_0[3118]); 
    assign layer_1[632] = layer_0[3461] & ~layer_0[3444]; 
    assign layer_1[633] = ~layer_0[2627] | (layer_0[2591] & layer_0[2627]); 
    assign layer_1[634] = layer_0[2655] & ~layer_0[2571]; 
    assign layer_1[635] = ~layer_0[2488] | (layer_0[2541] & layer_0[2488]); 
    assign layer_1[636] = layer_0[3599] & ~layer_0[3641]; 
    assign layer_1[637] = layer_0[3354] ^ layer_0[3257]; 
    assign layer_1[638] = ~layer_0[2935] | (layer_0[2935] & layer_0[2919]); 
    assign layer_1[639] = ~(layer_0[1851] ^ layer_0[1957]); 
    assign layer_1[640] = layer_0[3183] & ~layer_0[3239]; 
    assign layer_1[641] = ~layer_0[2436]; 
    assign layer_1[642] = ~layer_0[583]; 
    assign layer_1[643] = ~layer_0[3258]; 
    assign layer_1[644] = ~layer_0[1763]; 
    assign layer_1[645] = layer_0[298] ^ layer_0[209]; 
    assign layer_1[646] = ~layer_0[2649]; 
    assign layer_1[647] = ~layer_0[1794]; 
    assign layer_1[648] = layer_0[3143] & ~layer_0[3157]; 
    assign layer_1[649] = ~layer_0[886]; 
    assign layer_1[650] = ~layer_0[1297]; 
    assign layer_1[651] = layer_0[373] & ~layer_0[358]; 
    assign layer_1[652] = ~layer_0[2429]; 
    assign layer_1[653] = ~layer_0[1430]; 
    assign layer_1[654] = layer_0[836]; 
    assign layer_1[655] = ~layer_0[504]; 
    assign layer_1[656] = ~layer_0[3052]; 
    assign layer_1[657] = layer_0[1685] | layer_0[1727]; 
    assign layer_1[658] = ~(layer_0[3471] & layer_0[3478]); 
    assign layer_1[659] = ~(layer_0[124] ^ layer_0[131]); 
    assign layer_1[660] = ~(layer_0[3337] ^ layer_0[3291]); 
    assign layer_1[661] = layer_0[500]; 
    assign layer_1[662] = layer_0[1400]; 
    assign layer_1[663] = ~layer_0[3217]; 
    assign layer_1[664] = ~layer_0[1946] | (layer_0[1946] & layer_0[1855]); 
    assign layer_1[665] = ~layer_0[3442]; 
    assign layer_1[666] = ~layer_0[192]; 
    assign layer_1[667] = ~(layer_0[3680] ^ layer_0[3705]); 
    assign layer_1[668] = ~layer_0[3537] | (layer_0[3651] & layer_0[3537]); 
    assign layer_1[669] = ~(layer_0[2261] | layer_0[2371]); 
    assign layer_1[670] = layer_0[492] | layer_0[421]; 
    assign layer_1[671] = layer_0[1356] ^ layer_0[1481]; 
    assign layer_1[672] = layer_0[2879]; 
    assign layer_1[673] = layer_0[2883] | layer_0[2833]; 
    assign layer_1[674] = ~(layer_0[2221] & layer_0[2250]); 
    assign layer_1[675] = layer_0[1426] & layer_0[1435]; 
    assign layer_1[676] = layer_0[2231]; 
    assign layer_1[677] = ~layer_0[1344] | (layer_0[1257] & layer_0[1344]); 
    assign layer_1[678] = ~layer_0[3511] | (layer_0[3511] & layer_0[3488]); 
    assign layer_1[679] = ~(layer_0[1729] ^ layer_0[1642]); 
    assign layer_1[680] = layer_0[2365]; 
    assign layer_1[681] = layer_0[3200] & ~layer_0[3216]; 
    assign layer_1[682] = ~(layer_0[2024] ^ layer_0[2090]); 
    assign layer_1[683] = layer_0[679] & ~layer_0[735]; 
    assign layer_1[684] = layer_0[414] & ~layer_0[336]; 
    assign layer_1[685] = ~(layer_0[2809] & layer_0[2798]); 
    assign layer_1[686] = layer_0[1763]; 
    assign layer_1[687] = layer_0[12] ^ layer_0[106]; 
    assign layer_1[688] = ~(layer_0[3632] & layer_0[3528]); 
    assign layer_1[689] = layer_0[444] & ~layer_0[410]; 
    assign layer_1[690] = ~layer_0[3613]; 
    assign layer_1[691] = ~(layer_0[3242] ^ layer_0[3128]); 
    assign layer_1[692] = ~layer_0[172] | (layer_0[172] & layer_0[247]); 
    assign layer_1[693] = ~(layer_0[1720] & layer_0[1761]); 
    assign layer_1[694] = ~layer_0[2195]; 
    assign layer_1[695] = layer_0[9]; 
    assign layer_1[696] = ~(layer_0[2898] ^ layer_0[2940]); 
    assign layer_1[697] = layer_0[210] & ~layer_0[197]; 
    assign layer_1[698] = layer_0[1889] ^ layer_0[1783]; 
    assign layer_1[699] = layer_0[1736] ^ layer_0[1655]; 
    assign layer_1[700] = ~(layer_0[1450] ^ layer_0[1386]); 
    assign layer_1[701] = ~layer_0[1393]; 
    assign layer_1[702] = ~layer_0[586]; 
    assign layer_1[703] = layer_0[10]; 
    assign layer_1[704] = ~layer_0[3026]; 
    assign layer_1[705] = ~layer_0[1792]; 
    assign layer_1[706] = ~layer_0[3477]; 
    assign layer_1[707] = layer_0[564] & layer_0[610]; 
    assign layer_1[708] = layer_0[405] & ~layer_0[368]; 
    assign layer_1[709] = layer_0[2089] & ~layer_0[2037]; 
    assign layer_1[710] = ~layer_0[659]; 
    assign layer_1[711] = ~(layer_0[3366] | layer_0[3486]); 
    assign layer_1[712] = layer_0[22] & layer_0[143]; 
    assign layer_1[713] = layer_0[2215] & ~layer_0[2113]; 
    assign layer_1[714] = layer_0[2488] ^ layer_0[2445]; 
    assign layer_1[715] = layer_0[239]; 
    assign layer_1[716] = ~(layer_0[281] ^ layer_0[247]); 
    assign layer_1[717] = ~layer_0[461] | (layer_0[394] & layer_0[461]); 
    assign layer_1[718] = ~layer_0[740] | (layer_0[734] & layer_0[740]); 
    assign layer_1[719] = layer_0[1553] ^ layer_0[1550]; 
    assign layer_1[720] = layer_0[2484] & ~layer_0[2374]; 
    assign layer_1[721] = ~(layer_0[3123] & layer_0[3039]); 
    assign layer_1[722] = layer_0[3792] & layer_0[3776]; 
    assign layer_1[723] = layer_0[155]; 
    assign layer_1[724] = layer_0[2172]; 
    assign layer_1[725] = layer_0[3301] & layer_0[3215]; 
    assign layer_1[726] = ~layer_0[1148]; 
    assign layer_1[727] = ~(layer_0[2520] & layer_0[2488]); 
    assign layer_1[728] = layer_0[153] ^ layer_0[218]; 
    assign layer_1[729] = ~layer_0[527] | (layer_0[568] & layer_0[527]); 
    assign layer_1[730] = ~layer_0[360] | (layer_0[360] & layer_0[288]); 
    assign layer_1[731] = layer_0[2511] & ~layer_0[2614]; 
    assign layer_1[732] = layer_0[2451] & ~layer_0[2396]; 
    assign layer_1[733] = ~layer_0[2734]; 
    assign layer_1[734] = ~layer_0[3087]; 
    assign layer_1[735] = ~layer_0[547]; 
    assign layer_1[736] = ~(layer_0[3175] ^ layer_0[3146]); 
    assign layer_1[737] = ~layer_0[306]; 
    assign layer_1[738] = ~layer_0[3774]; 
    assign layer_1[739] = ~(layer_0[2074] ^ layer_0[2167]); 
    assign layer_1[740] = ~(layer_0[2084] ^ layer_0[1970]); 
    assign layer_1[741] = layer_0[2155] ^ layer_0[2044]; 
    assign layer_1[742] = layer_0[2156] ^ layer_0[2094]; 
    assign layer_1[743] = ~layer_0[1243]; 
    assign layer_1[744] = ~(layer_0[1489] & layer_0[1550]); 
    assign layer_1[745] = ~layer_0[657] | (layer_0[657] & layer_0[719]); 
    assign layer_1[746] = ~layer_0[327] | (layer_0[327] & layer_0[324]); 
    assign layer_1[747] = ~layer_0[2489]; 
    assign layer_1[748] = ~layer_0[962]; 
    assign layer_1[749] = ~layer_0[1600] | (layer_0[1600] & layer_0[1483]); 
    assign layer_1[750] = ~(layer_0[74] | layer_0[19]); 
    assign layer_1[751] = ~layer_0[358]; 
    assign layer_1[752] = layer_0[2109] ^ layer_0[2169]; 
    assign layer_1[753] = ~layer_0[1888] | (layer_0[1820] & layer_0[1888]); 
    assign layer_1[754] = layer_0[1618] | layer_0[1597]; 
    assign layer_1[755] = ~(layer_0[2493] ^ layer_0[2532]); 
    assign layer_1[756] = ~(layer_0[273] | layer_0[390]); 
    assign layer_1[757] = layer_0[118] ^ layer_0[101]; 
    assign layer_1[758] = ~(layer_0[2213] ^ layer_0[2202]); 
    assign layer_1[759] = ~layer_0[3877]; 
    assign layer_1[760] = ~(layer_0[439] | layer_0[485]); 
    assign layer_1[761] = layer_0[3056]; 
    assign layer_1[762] = ~layer_0[1828] | (layer_0[1828] & layer_0[1768]); 
    assign layer_1[763] = ~layer_0[1099] | (layer_0[1099] & layer_0[1068]); 
    assign layer_1[764] = layer_0[3429]; 
    assign layer_1[765] = ~layer_0[85]; 
    assign layer_1[766] = layer_0[880] & ~layer_0[833]; 
    assign layer_1[767] = ~(layer_0[2978] ^ layer_0[2888]); 
    assign layer_1[768] = layer_0[2378] | layer_0[2470]; 
    assign layer_1[769] = ~layer_0[1285] | (layer_0[1285] & layer_0[1277]); 
    assign layer_1[770] = layer_0[3036] | layer_0[3137]; 
    assign layer_1[771] = layer_0[2126]; 
    assign layer_1[772] = ~layer_0[1949]; 
    assign layer_1[773] = ~(layer_0[1482] & layer_0[1453]); 
    assign layer_1[774] = layer_0[3908] & layer_0[3945]; 
    assign layer_1[775] = layer_0[2319]; 
    assign layer_1[776] = ~layer_0[1314] | (layer_0[1314] & layer_0[1363]); 
    assign layer_1[777] = layer_0[1277] & ~layer_0[1281]; 
    assign layer_1[778] = layer_0[608] & layer_0[684]; 
    assign layer_1[779] = layer_0[1068]; 
    assign layer_1[780] = ~(layer_0[1703] | layer_0[1692]); 
    assign layer_1[781] = layer_0[1006]; 
    assign layer_1[782] = layer_0[3948]; 
    assign layer_1[783] = layer_0[106] & layer_0[98]; 
    assign layer_1[784] = ~layer_0[2882]; 
    assign layer_1[785] = ~layer_0[1612]; 
    assign layer_1[786] = layer_0[2628] | layer_0[2577]; 
    assign layer_1[787] = ~(layer_0[3750] ^ layer_0[3651]); 
    assign layer_1[788] = ~(layer_0[3824] & layer_0[3789]); 
    assign layer_1[789] = layer_0[1279]; 
    assign layer_1[790] = ~(layer_0[3549] | layer_0[3629]); 
    assign layer_1[791] = ~layer_0[3455] | (layer_0[3455] & layer_0[3567]); 
    assign layer_1[792] = layer_0[186]; 
    assign layer_1[793] = layer_0[1308] & ~layer_0[1277]; 
    assign layer_1[794] = layer_0[2477] ^ layer_0[2493]; 
    assign layer_1[795] = ~layer_0[1564] | (layer_0[1560] & layer_0[1564]); 
    assign layer_1[796] = ~(layer_0[2020] ^ layer_0[1948]); 
    assign layer_1[797] = ~layer_0[3991] | (layer_0[3996] & layer_0[3991]); 
    assign layer_1[798] = layer_0[3356] ^ layer_0[3483]; 
    assign layer_1[799] = ~(layer_0[3508] | layer_0[3618]); 
    assign layer_1[800] = layer_0[1185]; 
    assign layer_1[801] = layer_0[910] ^ layer_0[859]; 
    assign layer_1[802] = layer_0[1009] & layer_0[958]; 
    assign layer_1[803] = layer_0[182] ^ layer_0[227]; 
    assign layer_1[804] = layer_0[1218] & layer_0[1223]; 
    assign layer_1[805] = layer_0[801] & ~layer_0[910]; 
    assign layer_1[806] = layer_0[810] & ~layer_0[709]; 
    assign layer_1[807] = ~(layer_0[941] ^ layer_0[913]); 
    assign layer_1[808] = layer_0[873] | layer_0[826]; 
    assign layer_1[809] = ~layer_0[1493]; 
    assign layer_1[810] = layer_0[1766]; 
    assign layer_1[811] = ~layer_0[818] | (layer_0[818] & layer_0[726]); 
    assign layer_1[812] = ~(layer_0[2110] | layer_0[2043]); 
    assign layer_1[813] = layer_0[722] & layer_0[767]; 
    assign layer_1[814] = layer_0[511] & layer_0[443]; 
    assign layer_1[815] = layer_0[2528] & layer_0[2448]; 
    assign layer_1[816] = layer_0[2727] ^ layer_0[2623]; 
    assign layer_1[817] = ~(layer_0[2445] ^ layer_0[2396]); 
    assign layer_1[818] = layer_0[213] & ~layer_0[211]; 
    assign layer_1[819] = layer_0[2727] & layer_0[2818]; 
    assign layer_1[820] = ~(layer_0[790] & layer_0[763]); 
    assign layer_1[821] = layer_0[1301]; 
    assign layer_1[822] = layer_0[1783]; 
    assign layer_1[823] = layer_0[3973] & ~layer_0[3979]; 
    assign layer_1[824] = layer_0[673]; 
    assign layer_1[825] = layer_0[3444] | layer_0[3545]; 
    assign layer_1[826] = ~(layer_0[3680] & layer_0[3578]); 
    assign layer_1[827] = layer_0[2429]; 
    assign layer_1[828] = layer_0[1263] & ~layer_0[1266]; 
    assign layer_1[829] = layer_0[261] & ~layer_0[165]; 
    assign layer_1[830] = ~layer_0[260] | (layer_0[260] & layer_0[210]); 
    assign layer_1[831] = layer_0[1540] | layer_0[1626]; 
    assign layer_1[832] = layer_0[3201]; 
    assign layer_1[833] = ~(layer_0[1989] ^ layer_0[1982]); 
    assign layer_1[834] = ~layer_0[2847]; 
    assign layer_1[835] = layer_0[356] & ~layer_0[244]; 
    assign layer_1[836] = layer_0[2026] & ~layer_0[1966]; 
    assign layer_1[837] = layer_0[2250] & ~layer_0[2176]; 
    assign layer_1[838] = ~layer_0[860]; 
    assign layer_1[839] = layer_0[1265] & ~layer_0[1268]; 
    assign layer_1[840] = layer_0[3399]; 
    assign layer_1[841] = layer_0[632] & ~layer_0[594]; 
    assign layer_1[842] = ~(layer_0[1894] & layer_0[1847]); 
    assign layer_1[843] = ~(layer_0[2123] ^ layer_0[2129]); 
    assign layer_1[844] = layer_0[2319]; 
    assign layer_1[845] = ~(layer_0[2345] | layer_0[2274]); 
    assign layer_1[846] = ~layer_0[2176]; 
    assign layer_1[847] = ~(layer_0[3292] ^ layer_0[3217]); 
    assign layer_1[848] = ~layer_0[3412] | (layer_0[3412] & layer_0[3502]); 
    assign layer_1[849] = ~layer_0[1712]; 
    assign layer_1[850] = ~(layer_0[3821] & layer_0[3809]); 
    assign layer_1[851] = ~layer_0[2303]; 
    assign layer_1[852] = ~layer_0[3275] | (layer_0[3275] & layer_0[3220]); 
    assign layer_1[853] = layer_0[2675] & layer_0[2608]; 
    assign layer_1[854] = layer_0[892]; 
    assign layer_1[855] = layer_0[3102]; 
    assign layer_1[856] = ~layer_0[2582]; 
    assign layer_1[857] = ~layer_0[2851]; 
    assign layer_1[858] = ~(layer_0[135] & layer_0[161]); 
    assign layer_1[859] = layer_0[148] & ~layer_0[99]; 
    assign layer_1[860] = layer_0[733]; 
    assign layer_1[861] = ~(layer_0[3597] ^ layer_0[3706]); 
    assign layer_1[862] = layer_0[75] ^ layer_0[198]; 
    assign layer_1[863] = ~(layer_0[2883] & layer_0[2962]); 
    assign layer_1[864] = layer_0[2285] & ~layer_0[2390]; 
    assign layer_1[865] = ~layer_0[259]; 
    assign layer_1[866] = ~layer_0[2027]; 
    assign layer_1[867] = ~layer_0[2745] | (layer_0[2745] & layer_0[2846]); 
    assign layer_1[868] = ~layer_0[3467]; 
    assign layer_1[869] = ~(layer_0[3086] & layer_0[3014]); 
    assign layer_1[870] = layer_0[2587] & layer_0[2674]; 
    assign layer_1[871] = layer_0[1037] & ~layer_0[985]; 
    assign layer_1[872] = ~layer_0[1543]; 
    assign layer_1[873] = layer_0[446]; 
    assign layer_1[874] = ~(layer_0[1543] & layer_0[1485]); 
    assign layer_1[875] = layer_0[3888] & layer_0[3995]; 
    assign layer_1[876] = ~layer_0[3013] | (layer_0[3008] & layer_0[3013]); 
    assign layer_1[877] = ~(layer_0[478] ^ layer_0[506]); 
    assign layer_1[878] = layer_0[1560] | layer_0[1461]; 
    assign layer_1[879] = ~(layer_0[3051] | layer_0[3050]); 
    assign layer_1[880] = ~(layer_0[2497] | layer_0[2544]); 
    assign layer_1[881] = ~(layer_0[542] | layer_0[646]); 
    assign layer_1[882] = ~layer_0[3837] | (layer_0[3874] & layer_0[3837]); 
    assign layer_1[883] = ~layer_0[2572]; 
    assign layer_1[884] = layer_0[1409] & ~layer_0[1323]; 
    assign layer_1[885] = layer_0[209] & ~layer_0[154]; 
    assign layer_1[886] = layer_0[988] & ~layer_0[985]; 
    assign layer_1[887] = layer_0[157] & ~layer_0[217]; 
    assign layer_1[888] = layer_0[3509] & layer_0[3409]; 
    assign layer_1[889] = ~layer_0[1499]; 
    assign layer_1[890] = layer_0[1469] & ~layer_0[1510]; 
    assign layer_1[891] = ~(layer_0[3673] | layer_0[3575]); 
    assign layer_1[892] = ~(layer_0[1221] & layer_0[1290]); 
    assign layer_1[893] = ~(layer_0[1306] ^ layer_0[1282]); 
    assign layer_1[894] = ~(layer_0[2479] & layer_0[2475]); 
    assign layer_1[895] = layer_0[2322] & ~layer_0[2305]; 
    assign layer_1[896] = ~layer_0[2837]; 
    assign layer_1[897] = ~layer_0[2216]; 
    assign layer_1[898] = layer_0[2651] ^ layer_0[2557]; 
    assign layer_1[899] = layer_0[2849] ^ layer_0[2939]; 
    assign layer_1[900] = ~(layer_0[3843] ^ layer_0[3893]); 
    assign layer_1[901] = ~layer_0[947] | (layer_0[1043] & layer_0[947]); 
    assign layer_1[902] = ~layer_0[1788] | (layer_0[1890] & layer_0[1788]); 
    assign layer_1[903] = ~layer_0[948]; 
    assign layer_1[904] = layer_0[1278]; 
    assign layer_1[905] = ~layer_0[3577] | (layer_0[3518] & layer_0[3577]); 
    assign layer_1[906] = ~(layer_0[1857] | layer_0[1768]); 
    assign layer_1[907] = layer_0[1029] & ~layer_0[956]; 
    assign layer_1[908] = ~layer_0[3795] | (layer_0[3795] & layer_0[3806]); 
    assign layer_1[909] = ~(layer_0[1075] & layer_0[1103]); 
    assign layer_1[910] = layer_0[2150]; 
    assign layer_1[911] = ~layer_0[2153]; 
    assign layer_1[912] = ~layer_0[3941]; 
    assign layer_1[913] = layer_0[3194]; 
    assign layer_1[914] = layer_0[1815]; 
    assign layer_1[915] = ~layer_0[912] | (layer_0[912] & layer_0[869]); 
    assign layer_1[916] = ~layer_0[616] | (layer_0[652] & layer_0[616]); 
    assign layer_1[917] = ~(layer_0[2487] | layer_0[2453]); 
    assign layer_1[918] = ~layer_0[476]; 
    assign layer_1[919] = ~(layer_0[1696] ^ layer_0[1658]); 
    assign layer_1[920] = ~layer_0[3426] | (layer_0[3310] & layer_0[3426]); 
    assign layer_1[921] = layer_0[1544] ^ layer_0[1432]; 
    assign layer_1[922] = layer_0[1611]; 
    assign layer_1[923] = ~layer_0[667] | (layer_0[545] & layer_0[667]); 
    assign layer_1[924] = ~layer_0[2401]; 
    assign layer_1[925] = ~(layer_0[106] | layer_0[141]); 
    assign layer_1[926] = layer_0[162] & ~layer_0[175]; 
    assign layer_1[927] = ~layer_0[850]; 
    assign layer_1[928] = layer_0[1553] & ~layer_0[1594]; 
    assign layer_1[929] = ~layer_0[2480] | (layer_0[2480] & layer_0[2521]); 
    assign layer_1[930] = layer_0[1677]; 
    assign layer_1[931] = layer_0[943] & ~layer_0[964]; 
    assign layer_1[932] = layer_0[2404] & layer_0[2481]; 
    assign layer_1[933] = ~layer_0[2286]; 
    assign layer_1[934] = layer_0[2275] & layer_0[2206]; 
    assign layer_1[935] = ~layer_0[1914] | (layer_0[1941] & layer_0[1914]); 
    assign layer_1[936] = ~layer_0[2946]; 
    assign layer_1[937] = ~layer_0[3664] | (layer_0[3691] & layer_0[3664]); 
    assign layer_1[938] = ~(layer_0[173] ^ layer_0[52]); 
    assign layer_1[939] = ~layer_0[2108] | (layer_0[2108] & layer_0[2235]); 
    assign layer_1[940] = layer_0[2177]; 
    assign layer_1[941] = ~layer_0[215]; 
    assign layer_1[942] = layer_0[2527]; 
    assign layer_1[943] = ~(layer_0[24] | layer_0[118]); 
    assign layer_1[944] = ~layer_0[1055] | (layer_0[1055] & layer_0[1099]); 
    assign layer_1[945] = layer_0[2843] & ~layer_0[2924]; 
    assign layer_1[946] = layer_0[633] ^ layer_0[760]; 
    assign layer_1[947] = ~layer_0[974] | (layer_0[946] & layer_0[974]); 
    assign layer_1[948] = layer_0[3276] | layer_0[3178]; 
    assign layer_1[949] = layer_0[3074] & ~layer_0[3005]; 
    assign layer_1[950] = layer_0[753] & layer_0[752]; 
    assign layer_1[951] = layer_0[2864]; 
    assign layer_1[952] = ~layer_0[2969] | (layer_0[2969] & layer_0[2971]); 
    assign layer_1[953] = layer_0[1601] & ~layer_0[1632]; 
    assign layer_1[954] = layer_0[3158] | layer_0[3052]; 
    assign layer_1[955] = ~layer_0[1844] | (layer_0[1844] & layer_0[1736]); 
    assign layer_1[956] = ~layer_0[2808] | (layer_0[2808] & layer_0[2929]); 
    assign layer_1[957] = ~layer_0[2535] | (layer_0[2535] & layer_0[2623]); 
    assign layer_1[958] = ~layer_0[735]; 
    assign layer_1[959] = ~layer_0[2629] | (layer_0[2629] & layer_0[2523]); 
    assign layer_1[960] = layer_0[1485]; 
    assign layer_1[961] = layer_0[3570] & ~layer_0[3622]; 
    assign layer_1[962] = ~layer_0[3612]; 
    assign layer_1[963] = ~layer_0[369]; 
    assign layer_1[964] = layer_0[3656] & ~layer_0[3723]; 
    assign layer_1[965] = layer_0[2619] ^ layer_0[2666]; 
    assign layer_1[966] = layer_0[2021] & ~layer_0[2001]; 
    assign layer_1[967] = layer_0[971] ^ layer_0[857]; 
    assign layer_1[968] = ~(layer_0[1973] ^ layer_0[1998]); 
    assign layer_1[969] = ~(layer_0[1327] ^ layer_0[1204]); 
    assign layer_1[970] = layer_0[2648] | layer_0[2531]; 
    assign layer_1[971] = layer_0[2819]; 
    assign layer_1[972] = ~layer_0[861] | (layer_0[941] & layer_0[861]); 
    assign layer_1[973] = layer_0[1013] & ~layer_0[972]; 
    assign layer_1[974] = layer_0[328] | layer_0[264]; 
    assign layer_1[975] = layer_0[707]; 
    assign layer_1[976] = layer_0[564] ^ layer_0[536]; 
    assign layer_1[977] = layer_0[2423] ^ layer_0[2425]; 
    assign layer_1[978] = ~layer_0[883]; 
    assign layer_1[979] = ~(layer_0[1946] ^ layer_0[1923]); 
    assign layer_1[980] = layer_0[2775] ^ layer_0[2751]; 
    assign layer_1[981] = layer_0[2090]; 
    assign layer_1[982] = layer_0[2339] ^ layer_0[2340]; 
    assign layer_1[983] = ~layer_0[3327]; 
    assign layer_1[984] = ~layer_0[3576] | (layer_0[3576] & layer_0[3610]); 
    assign layer_1[985] = layer_0[3977]; 
    assign layer_1[986] = ~(layer_0[3066] & layer_0[3054]); 
    assign layer_1[987] = ~layer_0[807]; 
    assign layer_1[988] = layer_0[3870]; 
    assign layer_1[989] = ~(layer_0[2217] | layer_0[2248]); 
    assign layer_1[990] = ~(layer_0[307] & layer_0[187]); 
    assign layer_1[991] = ~layer_0[2946] | (layer_0[2946] & layer_0[2824]); 
    assign layer_1[992] = layer_0[2405]; 
    assign layer_1[993] = ~layer_0[848]; 
    assign layer_1[994] = ~(layer_0[3438] | layer_0[3477]); 
    assign layer_1[995] = layer_0[2293] & layer_0[2404]; 
    assign layer_1[996] = ~layer_0[3129]; 
    assign layer_1[997] = layer_0[636] ^ layer_0[688]; 
    assign layer_1[998] = layer_0[781]; 
    assign layer_1[999] = ~layer_0[3281]; 
    assign layer_1[1000] = ~(layer_0[741] ^ layer_0[680]); 
    assign layer_1[1001] = ~layer_0[1784] | (layer_0[1821] & layer_0[1784]); 
    assign layer_1[1002] = layer_0[1566] ^ layer_0[1546]; 
    assign layer_1[1003] = layer_0[1081]; 
    assign layer_1[1004] = layer_0[1555]; 
    assign layer_1[1005] = layer_0[1333] | layer_0[1274]; 
    assign layer_1[1006] = layer_0[720] ^ layer_0[685]; 
    assign layer_1[1007] = layer_0[757] ^ layer_0[785]; 
    assign layer_1[1008] = layer_0[2984]; 
    assign layer_1[1009] = ~(layer_0[1547] ^ layer_0[1667]); 
    assign layer_1[1010] = ~layer_0[3662]; 
    assign layer_1[1011] = ~(layer_0[2043] ^ layer_0[2045]); 
    assign layer_1[1012] = layer_0[2662]; 
    assign layer_1[1013] = ~(layer_0[3118] & layer_0[3069]); 
    assign layer_1[1014] = ~layer_0[1829] | (layer_0[1864] & layer_0[1829]); 
    assign layer_1[1015] = layer_0[3157]; 
    assign layer_1[1016] = ~layer_0[3889] | (layer_0[3889] & layer_0[3924]); 
    assign layer_1[1017] = ~(layer_0[3584] ^ layer_0[3517]); 
    assign layer_1[1018] = ~layer_0[3196] | (layer_0[3109] & layer_0[3196]); 
    assign layer_1[1019] = ~layer_0[229]; 
    assign layer_1[1020] = layer_0[2051]; 
    assign layer_1[1021] = layer_0[361] | layer_0[411]; 
    assign layer_1[1022] = ~layer_0[2407]; 
    assign layer_1[1023] = layer_0[2825] & ~layer_0[2764]; 
    assign layer_1[1024] = ~layer_0[704]; 
    assign layer_1[1025] = ~(layer_0[1746] ^ layer_0[1668]); 
    assign layer_1[1026] = ~layer_0[913]; 
    assign layer_1[1027] = ~(layer_0[3109] | layer_0[3062]); 
    assign layer_1[1028] = layer_0[2197] ^ layer_0[2149]; 
    assign layer_1[1029] = ~layer_0[2533]; 
    assign layer_1[1030] = layer_0[3208] & ~layer_0[3124]; 
    assign layer_1[1031] = layer_0[748] & layer_0[635]; 
    assign layer_1[1032] = layer_0[1008] | layer_0[1066]; 
    assign layer_1[1033] = ~layer_0[3991]; 
    assign layer_1[1034] = ~layer_0[554]; 
    assign layer_1[1035] = ~layer_0[795] | (layer_0[677] & layer_0[795]); 
    assign layer_1[1036] = layer_0[1587] ^ layer_0[1646]; 
    assign layer_1[1037] = layer_0[3259] & ~layer_0[3327]; 
    assign layer_1[1038] = ~layer_0[2194] | (layer_0[2194] & layer_0[2274]); 
    assign layer_1[1039] = ~(layer_0[3496] & layer_0[3572]); 
    assign layer_1[1040] = layer_0[1401] | layer_0[1397]; 
    assign layer_1[1041] = layer_0[1567] & ~layer_0[1517]; 
    assign layer_1[1042] = ~(layer_0[1574] ^ layer_0[1643]); 
    assign layer_1[1043] = ~layer_0[1028]; 
    assign layer_1[1044] = layer_0[1853] & ~layer_0[1975]; 
    assign layer_1[1045] = layer_0[2659] ^ layer_0[2558]; 
    assign layer_1[1046] = ~(layer_0[29] | layer_0[89]); 
    assign layer_1[1047] = layer_0[2269] & ~layer_0[2303]; 
    assign layer_1[1048] = layer_0[1646]; 
    assign layer_1[1049] = layer_0[3416] & layer_0[3467]; 
    assign layer_1[1050] = layer_0[3898] | layer_0[3786]; 
    assign layer_1[1051] = ~layer_0[1319] | (layer_0[1392] & layer_0[1319]); 
    assign layer_1[1052] = layer_0[419]; 
    assign layer_1[1053] = ~layer_0[2752] | (layer_0[2799] & layer_0[2752]); 
    assign layer_1[1054] = ~layer_0[1075] | (layer_0[1075] & layer_0[982]); 
    assign layer_1[1055] = ~layer_0[884]; 
    assign layer_1[1056] = layer_0[1225] & ~layer_0[1347]; 
    assign layer_1[1057] = ~layer_0[3772]; 
    assign layer_1[1058] = ~(layer_0[1796] | layer_0[1739]); 
    assign layer_1[1059] = layer_0[2044] ^ layer_0[2061]; 
    assign layer_1[1060] = ~layer_0[3945] | (layer_0[3944] & layer_0[3945]); 
    assign layer_1[1061] = ~(layer_0[1717] | layer_0[1739]); 
    assign layer_1[1062] = layer_0[2558]; 
    assign layer_1[1063] = layer_0[2098] | layer_0[2151]; 
    assign layer_1[1064] = ~(layer_0[776] & layer_0[881]); 
    assign layer_1[1065] = layer_0[423] | layer_0[342]; 
    assign layer_1[1066] = layer_0[2779] & layer_0[2862]; 
    assign layer_1[1067] = layer_0[2036]; 
    assign layer_1[1068] = layer_0[1552] & ~layer_0[1438]; 
    assign layer_1[1069] = ~(layer_0[1154] & layer_0[1129]); 
    assign layer_1[1070] = layer_0[2169]; 
    assign layer_1[1071] = layer_0[2056]; 
    assign layer_1[1072] = ~(layer_0[451] ^ layer_0[475]); 
    assign layer_1[1073] = ~layer_0[2492] | (layer_0[2492] & layer_0[2590]); 
    assign layer_1[1074] = ~layer_0[1977] | (layer_0[2000] & layer_0[1977]); 
    assign layer_1[1075] = ~layer_0[450] | (layer_0[396] & layer_0[450]); 
    assign layer_1[1076] = layer_0[3676] & ~layer_0[3745]; 
    assign layer_1[1077] = ~(layer_0[3518] | layer_0[3485]); 
    assign layer_1[1078] = layer_0[2047]; 
    assign layer_1[1079] = layer_0[3813] & layer_0[3872]; 
    assign layer_1[1080] = ~layer_0[2230]; 
    assign layer_1[1081] = ~(layer_0[3459] & layer_0[3562]); 
    assign layer_1[1082] = ~layer_0[2415] | (layer_0[2415] & layer_0[2342]); 
    assign layer_1[1083] = layer_0[1449] & ~layer_0[1462]; 
    assign layer_1[1084] = layer_0[1925] & ~layer_0[1860]; 
    assign layer_1[1085] = ~layer_0[332] | (layer_0[390] & layer_0[332]); 
    assign layer_1[1086] = layer_0[3314]; 
    assign layer_1[1087] = layer_0[1477]; 
    assign layer_1[1088] = ~layer_0[187]; 
    assign layer_1[1089] = ~(layer_0[472] ^ layer_0[392]); 
    assign layer_1[1090] = layer_0[3703]; 
    assign layer_1[1091] = ~layer_0[2445] | (layer_0[2539] & layer_0[2445]); 
    assign layer_1[1092] = layer_0[2879] ^ layer_0[2881]; 
    assign layer_1[1093] = ~layer_0[3188] | (layer_0[3188] & layer_0[3100]); 
    assign layer_1[1094] = layer_0[1508] & layer_0[1408]; 
    assign layer_1[1095] = ~layer_0[3615]; 
    assign layer_1[1096] = layer_0[1948] & layer_0[1909]; 
    assign layer_1[1097] = ~layer_0[212] | (layer_0[212] & layer_0[87]); 
    assign layer_1[1098] = layer_0[2691] ^ layer_0[2745]; 
    assign layer_1[1099] = layer_0[3584]; 
    assign layer_1[1100] = layer_0[716] ^ layer_0[817]; 
    assign layer_1[1101] = layer_0[3512]; 
    assign layer_1[1102] = layer_0[966] & ~layer_0[855]; 
    assign layer_1[1103] = layer_0[3689]; 
    assign layer_1[1104] = layer_0[3577]; 
    assign layer_1[1105] = layer_0[3825] & layer_0[3872]; 
    assign layer_1[1106] = ~(layer_0[2306] ^ layer_0[2215]); 
    assign layer_1[1107] = layer_0[1365] ^ layer_0[1468]; 
    assign layer_1[1108] = ~(layer_0[1428] ^ layer_0[1454]); 
    assign layer_1[1109] = layer_0[3519] & ~layer_0[3509]; 
    assign layer_1[1110] = ~layer_0[803] | (layer_0[675] & layer_0[803]); 
    assign layer_1[1111] = ~layer_0[3719]; 
    assign layer_1[1112] = ~(layer_0[1930] | layer_0[1877]); 
    assign layer_1[1113] = layer_0[1224]; 
    assign layer_1[1114] = layer_0[3361]; 
    assign layer_1[1115] = layer_0[1372] ^ layer_0[1375]; 
    assign layer_1[1116] = ~(layer_0[1353] ^ layer_0[1229]); 
    assign layer_1[1117] = layer_0[975] & layer_0[869]; 
    assign layer_1[1118] = layer_0[3491] & ~layer_0[3418]; 
    assign layer_1[1119] = ~(layer_0[2016] & layer_0[1951]); 
    assign layer_1[1120] = ~layer_0[2222]; 
    assign layer_1[1121] = layer_0[1108] & ~layer_0[1071]; 
    assign layer_1[1122] = layer_0[3296] & ~layer_0[3262]; 
    assign layer_1[1123] = layer_0[3211] | layer_0[3324]; 
    assign layer_1[1124] = layer_0[2724] & ~layer_0[2796]; 
    assign layer_1[1125] = ~(layer_0[3386] & layer_0[3427]); 
    assign layer_1[1126] = layer_0[1051] | layer_0[1002]; 
    assign layer_1[1127] = layer_0[2304] | layer_0[2319]; 
    assign layer_1[1128] = ~(layer_0[362] & layer_0[413]); 
    assign layer_1[1129] = layer_0[1406] & layer_0[1508]; 
    assign layer_1[1130] = layer_0[3878] | layer_0[3905]; 
    assign layer_1[1131] = layer_0[1025]; 
    assign layer_1[1132] = ~layer_0[1469] | (layer_0[1397] & layer_0[1469]); 
    assign layer_1[1133] = ~(layer_0[1103] ^ layer_0[992]); 
    assign layer_1[1134] = layer_0[3706]; 
    assign layer_1[1135] = layer_0[1093]; 
    assign layer_1[1136] = layer_0[468] ^ layer_0[380]; 
    assign layer_1[1137] = layer_0[3167] & ~layer_0[3128]; 
    assign layer_1[1138] = ~layer_0[243] | (layer_0[123] & layer_0[243]); 
    assign layer_1[1139] = ~(layer_0[3765] | layer_0[3820]); 
    assign layer_1[1140] = ~(layer_0[2434] ^ layer_0[2442]); 
    assign layer_1[1141] = ~layer_0[2830] | (layer_0[2702] & layer_0[2830]); 
    assign layer_1[1142] = layer_0[3764]; 
    assign layer_1[1143] = layer_0[1716]; 
    assign layer_1[1144] = layer_0[2769]; 
    assign layer_1[1145] = ~layer_0[2976]; 
    assign layer_1[1146] = ~layer_0[1082]; 
    assign layer_1[1147] = layer_0[1043]; 
    assign layer_1[1148] = ~layer_0[3953]; 
    assign layer_1[1149] = ~(layer_0[384] ^ layer_0[375]); 
    assign layer_1[1150] = ~(layer_0[3961] & layer_0[3955]); 
    assign layer_1[1151] = layer_0[2660] ^ layer_0[2691]; 
    assign layer_1[1152] = ~(layer_0[1503] & layer_0[1493]); 
    assign layer_1[1153] = ~layer_0[1528] | (layer_0[1528] & layer_0[1600]); 
    assign layer_1[1154] = ~layer_0[2738] | (layer_0[2778] & layer_0[2738]); 
    assign layer_1[1155] = layer_0[1124] ^ layer_0[1029]; 
    assign layer_1[1156] = layer_0[2247] & ~layer_0[2283]; 
    assign layer_1[1157] = ~layer_0[2031]; 
    assign layer_1[1158] = layer_0[498]; 
    assign layer_1[1159] = layer_0[3757]; 
    assign layer_1[1160] = ~layer_0[1199] | (layer_0[1262] & layer_0[1199]); 
    assign layer_1[1161] = ~(layer_0[2704] & layer_0[2730]); 
    assign layer_1[1162] = ~(layer_0[2775] & layer_0[2880]); 
    assign layer_1[1163] = layer_0[3037] & ~layer_0[2917]; 
    assign layer_1[1164] = ~layer_0[1165]; 
    assign layer_1[1165] = ~layer_0[346] | (layer_0[346] & layer_0[268]); 
    assign layer_1[1166] = ~(layer_0[374] ^ layer_0[437]); 
    assign layer_1[1167] = layer_0[1055] & ~layer_0[1173]; 
    assign layer_1[1168] = layer_0[3526]; 
    assign layer_1[1169] = layer_0[1942] & ~layer_0[1977]; 
    assign layer_1[1170] = ~layer_0[1530] | (layer_0[1530] & layer_0[1505]); 
    assign layer_1[1171] = ~layer_0[308]; 
    assign layer_1[1172] = layer_0[2667] & layer_0[2570]; 
    assign layer_1[1173] = ~layer_0[2916]; 
    assign layer_1[1174] = ~(layer_0[2539] | layer_0[2456]); 
    assign layer_1[1175] = layer_0[206]; 
    assign layer_1[1176] = ~(layer_0[2241] & layer_0[2259]); 
    assign layer_1[1177] = ~(layer_0[1744] | layer_0[1727]); 
    assign layer_1[1178] = ~layer_0[1981]; 
    assign layer_1[1179] = layer_0[2181]; 
    assign layer_1[1180] = ~layer_0[780] | (layer_0[801] & layer_0[780]); 
    assign layer_1[1181] = layer_0[526] | layer_0[463]; 
    assign layer_1[1182] = layer_0[2768]; 
    assign layer_1[1183] = ~(layer_0[3747] ^ layer_0[3852]); 
    assign layer_1[1184] = ~layer_0[1249] | (layer_0[1249] & layer_0[1204]); 
    assign layer_1[1185] = ~(layer_0[3758] | layer_0[3657]); 
    assign layer_1[1186] = layer_0[2927] & layer_0[2820]; 
    assign layer_1[1187] = layer_0[645]; 
    assign layer_1[1188] = ~layer_0[535]; 
    assign layer_1[1189] = ~(layer_0[1780] | layer_0[1792]); 
    assign layer_1[1190] = layer_0[1051]; 
    assign layer_1[1191] = ~layer_0[2932]; 
    assign layer_1[1192] = ~(layer_0[3199] ^ layer_0[3200]); 
    assign layer_1[1193] = layer_0[3456] & layer_0[3519]; 
    assign layer_1[1194] = layer_0[2719] & ~layer_0[2726]; 
    assign layer_1[1195] = layer_0[1113] & ~layer_0[1227]; 
    assign layer_1[1196] = ~layer_0[1349]; 
    assign layer_1[1197] = layer_0[20] & layer_0[85]; 
    assign layer_1[1198] = layer_0[3902] ^ layer_0[3908]; 
    assign layer_1[1199] = ~layer_0[432] | (layer_0[432] & layer_0[411]); 
    assign layer_1[1200] = layer_0[1132] & ~layer_0[1229]; 
    assign layer_1[1201] = ~layer_0[342]; 
    assign layer_1[1202] = ~layer_0[2792] | (layer_0[2838] & layer_0[2792]); 
    assign layer_1[1203] = layer_0[187] & ~layer_0[66]; 
    assign layer_1[1204] = ~(layer_0[2030] | layer_0[1989]); 
    assign layer_1[1205] = ~layer_0[1745]; 
    assign layer_1[1206] = ~layer_0[3732]; 
    assign layer_1[1207] = ~(layer_0[3268] ^ layer_0[3280]); 
    assign layer_1[1208] = layer_0[3418] | layer_0[3501]; 
    assign layer_1[1209] = ~layer_0[1254]; 
    assign layer_1[1210] = layer_0[2855]; 
    assign layer_1[1211] = ~(layer_0[764] ^ layer_0[716]); 
    assign layer_1[1212] = layer_0[2039] & ~layer_0[2137]; 
    assign layer_1[1213] = ~layer_0[108] | (layer_0[141] & layer_0[108]); 
    assign layer_1[1214] = layer_0[2380] ^ layer_0[2328]; 
    assign layer_1[1215] = layer_0[3658]; 
    assign layer_1[1216] = layer_0[1448]; 
    assign layer_1[1217] = ~(layer_0[3467] ^ layer_0[3493]); 
    assign layer_1[1218] = layer_0[1334] & ~layer_0[1327]; 
    assign layer_1[1219] = layer_0[1330]; 
    assign layer_1[1220] = layer_0[490] ^ layer_0[545]; 
    assign layer_1[1221] = layer_0[255] & layer_0[249]; 
    assign layer_1[1222] = layer_0[2600] | layer_0[2546]; 
    assign layer_1[1223] = ~layer_0[348] | (layer_0[348] & layer_0[411]); 
    assign layer_1[1224] = ~layer_0[2139] | (layer_0[2148] & layer_0[2139]); 
    assign layer_1[1225] = ~layer_0[735]; 
    assign layer_1[1226] = layer_0[2688] & layer_0[2671]; 
    assign layer_1[1227] = layer_0[2566]; 
    assign layer_1[1228] = ~layer_0[2030] | (layer_0[2030] & layer_0[2110]); 
    assign layer_1[1229] = layer_0[2223] | layer_0[2156]; 
    assign layer_1[1230] = ~layer_0[3659] | (layer_0[3696] & layer_0[3659]); 
    assign layer_1[1231] = layer_0[909] | layer_0[841]; 
    assign layer_1[1232] = ~(layer_0[2335] ^ layer_0[2329]); 
    assign layer_1[1233] = layer_0[1165] & ~layer_0[1080]; 
    assign layer_1[1234] = layer_0[2132] | layer_0[2147]; 
    assign layer_1[1235] = ~layer_0[1944]; 
    assign layer_1[1236] = ~layer_0[3506] | (layer_0[3482] & layer_0[3506]); 
    assign layer_1[1237] = ~layer_0[1353] | (layer_0[1353] & layer_0[1243]); 
    assign layer_1[1238] = ~(layer_0[636] & layer_0[728]); 
    assign layer_1[1239] = layer_0[3530] & layer_0[3650]; 
    assign layer_1[1240] = ~(layer_0[2274] | layer_0[2366]); 
    assign layer_1[1241] = layer_0[312]; 
    assign layer_1[1242] = ~layer_0[2249]; 
    assign layer_1[1243] = ~layer_0[376]; 
    assign layer_1[1244] = layer_0[1109] & ~layer_0[1038]; 
    assign layer_1[1245] = layer_0[1426]; 
    assign layer_1[1246] = layer_0[2216] & ~layer_0[2156]; 
    assign layer_1[1247] = ~(layer_0[1395] ^ layer_0[1401]); 
    assign layer_1[1248] = layer_0[1763] & ~layer_0[1769]; 
    assign layer_1[1249] = ~layer_0[3458]; 
    assign layer_1[1250] = ~layer_0[467]; 
    assign layer_1[1251] = ~layer_0[2520]; 
    assign layer_1[1252] = layer_0[733]; 
    assign layer_1[1253] = ~layer_0[2894]; 
    assign layer_1[1254] = layer_0[2017] ^ layer_0[1950]; 
    assign layer_1[1255] = layer_0[540] & layer_0[534]; 
    assign layer_1[1256] = ~layer_0[3865]; 
    assign layer_1[1257] = layer_0[2018]; 
    assign layer_1[1258] = ~layer_0[1620] | (layer_0[1620] & layer_0[1600]); 
    assign layer_1[1259] = ~layer_0[2456] | (layer_0[2362] & layer_0[2456]); 
    assign layer_1[1260] = layer_0[1548]; 
    assign layer_1[1261] = ~(layer_0[2550] ^ layer_0[2453]); 
    assign layer_1[1262] = ~(layer_0[15] ^ layer_0[85]); 
    assign layer_1[1263] = layer_0[601]; 
    assign layer_1[1264] = ~(layer_0[1178] ^ layer_0[1135]); 
    assign layer_1[1265] = layer_0[348] | layer_0[252]; 
    assign layer_1[1266] = ~(layer_0[1072] ^ layer_0[963]); 
    assign layer_1[1267] = ~(layer_0[2147] ^ layer_0[2158]); 
    assign layer_1[1268] = layer_0[76] | layer_0[161]; 
    assign layer_1[1269] = ~(layer_0[1067] ^ layer_0[1050]); 
    assign layer_1[1270] = ~(layer_0[3321] ^ layer_0[3323]); 
    assign layer_1[1271] = layer_0[3551] & ~layer_0[3561]; 
    assign layer_1[1272] = layer_0[2108] & ~layer_0[2125]; 
    assign layer_1[1273] = ~(layer_0[2582] & layer_0[2559]); 
    assign layer_1[1274] = ~layer_0[3530] | (layer_0[3448] & layer_0[3530]); 
    assign layer_1[1275] = ~layer_0[319]; 
    assign layer_1[1276] = layer_0[1635]; 
    assign layer_1[1277] = layer_0[3636]; 
    assign layer_1[1278] = ~(layer_0[1547] ^ layer_0[1471]); 
    assign layer_1[1279] = ~layer_0[2931] | (layer_0[2931] & layer_0[2944]); 
    assign layer_1[1280] = layer_0[1984] | layer_0[1923]; 
    assign layer_1[1281] = ~layer_0[2421] | (layer_0[2421] & layer_0[2517]); 
    assign layer_1[1282] = ~layer_0[1433]; 
    assign layer_1[1283] = layer_0[3074] | layer_0[3163]; 
    assign layer_1[1284] = layer_0[2072]; 
    assign layer_1[1285] = layer_0[427] & ~layer_0[426]; 
    assign layer_1[1286] = ~layer_0[3325]; 
    assign layer_1[1287] = ~(layer_0[510] | layer_0[468]); 
    assign layer_1[1288] = layer_0[682] & layer_0[624]; 
    assign layer_1[1289] = ~(layer_0[1757] & layer_0[1779]); 
    assign layer_1[1290] = layer_0[576] & layer_0[494]; 
    assign layer_1[1291] = ~layer_0[2690] | (layer_0[2690] & layer_0[2767]); 
    assign layer_1[1292] = layer_0[1252] & layer_0[1132]; 
    assign layer_1[1293] = layer_0[573] | layer_0[517]; 
    assign layer_1[1294] = layer_0[3173]; 
    assign layer_1[1295] = layer_0[2380] ^ layer_0[2314]; 
    assign layer_1[1296] = layer_0[3810] & ~layer_0[3906]; 
    assign layer_1[1297] = layer_0[2097] & ~layer_0[2198]; 
    assign layer_1[1298] = layer_0[308] ^ layer_0[339]; 
    assign layer_1[1299] = ~(layer_0[3526] & layer_0[3608]); 
    assign layer_1[1300] = ~(layer_0[4] & layer_0[24]); 
    assign layer_1[1301] = layer_0[571] & layer_0[459]; 
    assign layer_1[1302] = ~layer_0[384]; 
    assign layer_1[1303] = ~layer_0[966]; 
    assign layer_1[1304] = ~(layer_0[461] & layer_0[470]); 
    assign layer_1[1305] = ~layer_0[396]; 
    assign layer_1[1306] = layer_0[2502] ^ layer_0[2497]; 
    assign layer_1[1307] = ~(layer_0[719] & layer_0[700]); 
    assign layer_1[1308] = ~layer_0[3214]; 
    assign layer_1[1309] = layer_0[492]; 
    assign layer_1[1310] = layer_0[1821] & ~layer_0[1904]; 
    assign layer_1[1311] = ~layer_0[1177]; 
    assign layer_1[1312] = ~layer_0[2443] | (layer_0[2443] & layer_0[2469]); 
    assign layer_1[1313] = layer_0[9]; 
    assign layer_1[1314] = layer_0[3987]; 
    assign layer_1[1315] = ~layer_0[1287]; 
    assign layer_1[1316] = layer_0[631] & ~layer_0[627]; 
    assign layer_1[1317] = layer_0[3297] | layer_0[3319]; 
    assign layer_1[1318] = ~(layer_0[1043] & layer_0[1062]); 
    assign layer_1[1319] = layer_0[548]; 
    assign layer_1[1320] = ~layer_0[3242] | (layer_0[3242] & layer_0[3135]); 
    assign layer_1[1321] = layer_0[333] & layer_0[348]; 
    assign layer_1[1322] = ~(layer_0[2567] ^ layer_0[2466]); 
    assign layer_1[1323] = layer_0[1542]; 
    assign layer_1[1324] = layer_0[3151]; 
    assign layer_1[1325] = ~layer_0[1781]; 
    assign layer_1[1326] = ~(layer_0[1278] ^ layer_0[1334]); 
    assign layer_1[1327] = ~(layer_0[1172] | layer_0[1192]); 
    assign layer_1[1328] = layer_0[955]; 
    assign layer_1[1329] = layer_0[2715] | layer_0[2763]; 
    assign layer_1[1330] = ~(layer_0[2127] & layer_0[2186]); 
    assign layer_1[1331] = layer_0[942] | layer_0[823]; 
    assign layer_1[1332] = layer_0[2713] & layer_0[2645]; 
    assign layer_1[1333] = layer_0[2365] & ~layer_0[2436]; 
    assign layer_1[1334] = ~layer_0[2335] | (layer_0[2335] & layer_0[2367]); 
    assign layer_1[1335] = layer_0[372] & layer_0[485]; 
    assign layer_1[1336] = layer_0[906] | layer_0[858]; 
    assign layer_1[1337] = ~layer_0[1151]; 
    assign layer_1[1338] = ~(layer_0[2881] | layer_0[2826]); 
    assign layer_1[1339] = ~layer_0[760] | (layer_0[718] & layer_0[760]); 
    assign layer_1[1340] = ~layer_0[233] | (layer_0[233] & layer_0[153]); 
    assign layer_1[1341] = ~layer_0[206]; 
    assign layer_1[1342] = ~(layer_0[208] & layer_0[197]); 
    assign layer_1[1343] = ~layer_0[49] | (layer_0[49] & layer_0[65]); 
    assign layer_1[1344] = layer_0[2558]; 
    assign layer_1[1345] = layer_0[1341] & ~layer_0[1357]; 
    assign layer_1[1346] = layer_0[3311]; 
    assign layer_1[1347] = ~(layer_0[3666] ^ layer_0[3694]); 
    assign layer_1[1348] = ~layer_0[2987] | (layer_0[2987] & layer_0[3083]); 
    assign layer_1[1349] = layer_0[1569]; 
    assign layer_1[1350] = layer_0[1384] ^ layer_0[1493]; 
    assign layer_1[1351] = layer_0[365]; 
    assign layer_1[1352] = ~(layer_0[3674] ^ layer_0[3682]); 
    assign layer_1[1353] = ~layer_0[555] | (layer_0[555] & layer_0[672]); 
    assign layer_1[1354] = layer_0[1831] & layer_0[1887]; 
    assign layer_1[1355] = ~(layer_0[3006] ^ layer_0[2924]); 
    assign layer_1[1356] = layer_0[129] ^ layer_0[53]; 
    assign layer_1[1357] = ~layer_0[3578]; 
    assign layer_1[1358] = ~layer_0[53] | (layer_0[19] & layer_0[53]); 
    assign layer_1[1359] = ~(layer_0[2616] | layer_0[2500]); 
    assign layer_1[1360] = ~layer_0[286]; 
    assign layer_1[1361] = layer_0[1089]; 
    assign layer_1[1362] = ~layer_0[352]; 
    assign layer_1[1363] = layer_0[930] & ~layer_0[980]; 
    assign layer_1[1364] = layer_0[783]; 
    assign layer_1[1365] = layer_0[195] & ~layer_0[244]; 
    assign layer_1[1366] = layer_0[3512]; 
    assign layer_1[1367] = layer_0[1958] | layer_0[1892]; 
    assign layer_1[1368] = layer_0[3742] & layer_0[3864]; 
    assign layer_1[1369] = ~layer_0[3207] | (layer_0[3207] & layer_0[3142]); 
    assign layer_1[1370] = layer_0[129] & ~layer_0[155]; 
    assign layer_1[1371] = ~layer_0[111] | (layer_0[50] & layer_0[111]); 
    assign layer_1[1372] = layer_0[3644] & ~layer_0[3684]; 
    assign layer_1[1373] = layer_0[1468] & ~layer_0[1530]; 
    assign layer_1[1374] = ~layer_0[3293]; 
    assign layer_1[1375] = layer_0[1232]; 
    assign layer_1[1376] = ~(layer_0[1233] | layer_0[1302]); 
    assign layer_1[1377] = ~layer_0[823] | (layer_0[823] & layer_0[751]); 
    assign layer_1[1378] = ~layer_0[2777] | (layer_0[2777] & layer_0[2668]); 
    assign layer_1[1379] = ~(layer_0[412] & layer_0[401]); 
    assign layer_1[1380] = ~layer_0[111]; 
    assign layer_1[1381] = ~layer_0[3178] | (layer_0[3178] & layer_0[3221]); 
    assign layer_1[1382] = ~layer_0[945]; 
    assign layer_1[1383] = ~layer_0[3393]; 
    assign layer_1[1384] = layer_0[2054]; 
    assign layer_1[1385] = layer_0[3204] | layer_0[3228]; 
    assign layer_1[1386] = ~layer_0[459]; 
    assign layer_1[1387] = layer_0[112] & ~layer_0[23]; 
    assign layer_1[1388] = layer_0[2737]; 
    assign layer_1[1389] = ~(layer_0[3662] | layer_0[3690]); 
    assign layer_1[1390] = layer_0[2402]; 
    assign layer_1[1391] = layer_0[1420] | layer_0[1504]; 
    assign layer_1[1392] = ~layer_0[3459]; 
    assign layer_1[1393] = layer_0[2297]; 
    assign layer_1[1394] = layer_0[3884] & ~layer_0[3872]; 
    assign layer_1[1395] = ~layer_0[1220] | (layer_0[1220] & layer_0[1259]); 
    assign layer_1[1396] = layer_0[615] & ~layer_0[488]; 
    assign layer_1[1397] = layer_0[2727] & ~layer_0[2823]; 
    assign layer_1[1398] = ~(layer_0[3506] & layer_0[3563]); 
    assign layer_1[1399] = layer_0[40] & layer_0[135]; 
    assign layer_1[1400] = layer_0[711]; 
    assign layer_1[1401] = layer_0[3324]; 
    assign layer_1[1402] = layer_0[623]; 
    assign layer_1[1403] = ~layer_0[2639] | (layer_0[2732] & layer_0[2639]); 
    assign layer_1[1404] = layer_0[2850] & ~layer_0[2910]; 
    assign layer_1[1405] = ~layer_0[2845]; 
    assign layer_1[1406] = layer_0[3190] & layer_0[3081]; 
    assign layer_1[1407] = ~(layer_0[714] ^ layer_0[673]); 
    assign layer_1[1408] = ~layer_0[1900]; 
    assign layer_1[1409] = ~(layer_0[64] ^ layer_0[127]); 
    assign layer_1[1410] = layer_0[2385]; 
    assign layer_1[1411] = layer_0[1390] & ~layer_0[1381]; 
    assign layer_1[1412] = ~(layer_0[1663] | layer_0[1780]); 
    assign layer_1[1413] = ~layer_0[3987]; 
    assign layer_1[1414] = layer_0[1214] ^ layer_0[1216]; 
    assign layer_1[1415] = layer_0[1898] | layer_0[1940]; 
    assign layer_1[1416] = ~layer_0[1718]; 
    assign layer_1[1417] = ~layer_0[494] | (layer_0[494] & layer_0[594]); 
    assign layer_1[1418] = layer_0[1558]; 
    assign layer_1[1419] = ~layer_0[516]; 
    assign layer_1[1420] = ~layer_0[1826]; 
    assign layer_1[1421] = ~(layer_0[1934] | layer_0[1977]); 
    assign layer_1[1422] = layer_0[1608] ^ layer_0[1584]; 
    assign layer_1[1423] = ~(layer_0[1370] & layer_0[1405]); 
    assign layer_1[1424] = ~(layer_0[1736] & layer_0[1722]); 
    assign layer_1[1425] = ~layer_0[102]; 
    assign layer_1[1426] = layer_0[1639] ^ layer_0[1682]; 
    assign layer_1[1427] = layer_0[158] | layer_0[257]; 
    assign layer_1[1428] = layer_0[3934] ^ layer_0[3882]; 
    assign layer_1[1429] = layer_0[2555] & ~layer_0[2617]; 
    assign layer_1[1430] = ~layer_0[1677]; 
    assign layer_1[1431] = layer_0[3666] & ~layer_0[3765]; 
    assign layer_1[1432] = ~layer_0[1659]; 
    assign layer_1[1433] = layer_0[495]; 
    assign layer_1[1434] = layer_0[3810] & ~layer_0[3860]; 
    assign layer_1[1435] = ~layer_0[3438]; 
    assign layer_1[1436] = ~layer_0[79]; 
    assign layer_1[1437] = layer_0[2959]; 
    assign layer_1[1438] = layer_0[949] & ~layer_0[1063]; 
    assign layer_1[1439] = layer_0[854] | layer_0[915]; 
    assign layer_1[1440] = ~(layer_0[960] | layer_0[953]); 
    assign layer_1[1441] = layer_0[1946] ^ layer_0[2058]; 
    assign layer_1[1442] = layer_0[1912]; 
    assign layer_1[1443] = ~layer_0[1301]; 
    assign layer_1[1444] = layer_0[2282] & layer_0[2197]; 
    assign layer_1[1445] = ~layer_0[2764] | (layer_0[2764] & layer_0[2723]); 
    assign layer_1[1446] = ~layer_0[2430]; 
    assign layer_1[1447] = layer_0[2917] ^ layer_0[2967]; 
    assign layer_1[1448] = layer_0[34] & ~layer_0[60]; 
    assign layer_1[1449] = layer_0[1102] & layer_0[1003]; 
    assign layer_1[1450] = ~(layer_0[1159] | layer_0[1128]); 
    assign layer_1[1451] = layer_0[1687] | layer_0[1579]; 
    assign layer_1[1452] = layer_0[330] | layer_0[360]; 
    assign layer_1[1453] = layer_0[3838]; 
    assign layer_1[1454] = layer_0[2570] & ~layer_0[2505]; 
    assign layer_1[1455] = ~layer_0[1033] | (layer_0[1033] & layer_0[999]); 
    assign layer_1[1456] = layer_0[772] & ~layer_0[711]; 
    assign layer_1[1457] = ~(layer_0[1017] | layer_0[1049]); 
    assign layer_1[1458] = layer_0[148] | layer_0[73]; 
    assign layer_1[1459] = layer_0[572] & layer_0[574]; 
    assign layer_1[1460] = layer_0[123] & layer_0[88]; 
    assign layer_1[1461] = ~layer_0[2771] | (layer_0[2893] & layer_0[2771]); 
    assign layer_1[1462] = layer_0[1935]; 
    assign layer_1[1463] = layer_0[3116] & layer_0[3161]; 
    assign layer_1[1464] = layer_0[237]; 
    assign layer_1[1465] = layer_0[1033]; 
    assign layer_1[1466] = ~(layer_0[1207] | layer_0[1150]); 
    assign layer_1[1467] = layer_0[3267] & ~layer_0[3337]; 
    assign layer_1[1468] = ~layer_0[965]; 
    assign layer_1[1469] = layer_0[2687] ^ layer_0[2711]; 
    assign layer_1[1470] = ~(layer_0[1929] | layer_0[2021]); 
    assign layer_1[1471] = ~layer_0[3079]; 
    assign layer_1[1472] = ~(layer_0[2224] & layer_0[2121]); 
    assign layer_1[1473] = ~layer_0[3996]; 
    assign layer_1[1474] = layer_0[3406] ^ layer_0[3439]; 
    assign layer_1[1475] = layer_0[1872]; 
    assign layer_1[1476] = layer_0[399] & ~layer_0[466]; 
    assign layer_1[1477] = layer_0[902] ^ layer_0[968]; 
    assign layer_1[1478] = layer_0[3095]; 
    assign layer_1[1479] = ~layer_0[2406]; 
    assign layer_1[1480] = layer_0[1644] ^ layer_0[1534]; 
    assign layer_1[1481] = ~(layer_0[1461] | layer_0[1508]); 
    assign layer_1[1482] = ~layer_0[2416] | (layer_0[2329] & layer_0[2416]); 
    assign layer_1[1483] = layer_0[713] ^ layer_0[826]; 
    assign layer_1[1484] = ~layer_0[3573] | (layer_0[3643] & layer_0[3573]); 
    assign layer_1[1485] = ~layer_0[357] | (layer_0[357] & layer_0[320]); 
    assign layer_1[1486] = layer_0[3540] & layer_0[3569]; 
    assign layer_1[1487] = layer_0[73] | layer_0[42]; 
    assign layer_1[1488] = layer_0[3966] | layer_0[3893]; 
    assign layer_1[1489] = layer_0[2900] & layer_0[2918]; 
    assign layer_1[1490] = layer_0[609] & layer_0[577]; 
    assign layer_1[1491] = layer_0[272]; 
    assign layer_1[1492] = ~layer_0[1101]; 
    assign layer_1[1493] = layer_0[3015] ^ layer_0[3076]; 
    assign layer_1[1494] = layer_0[1050] | layer_0[970]; 
    assign layer_1[1495] = ~layer_0[781]; 
    assign layer_1[1496] = ~layer_0[2608] | (layer_0[2608] & layer_0[2724]); 
    assign layer_1[1497] = ~(layer_0[3705] ^ layer_0[3676]); 
    assign layer_1[1498] = layer_0[1121]; 
    assign layer_1[1499] = ~(layer_0[1542] & layer_0[1612]); 
    assign layer_1[1500] = ~layer_0[470] | (layer_0[596] & layer_0[470]); 
    assign layer_1[1501] = ~layer_0[2359] | (layer_0[2359] & layer_0[2405]); 
    assign layer_1[1502] = ~(layer_0[2532] & layer_0[2660]); 
    assign layer_1[1503] = layer_0[1936]; 
    assign layer_1[1504] = layer_0[89]; 
    assign layer_1[1505] = layer_0[1085] ^ layer_0[1100]; 
    assign layer_1[1506] = layer_0[104]; 
    assign layer_1[1507] = layer_0[2962]; 
    assign layer_1[1508] = ~(layer_0[1654] | layer_0[1750]); 
    assign layer_1[1509] = ~(layer_0[3694] ^ layer_0[3705]); 
    assign layer_1[1510] = layer_0[3143]; 
    assign layer_1[1511] = ~(layer_0[1028] | layer_0[1092]); 
    assign layer_1[1512] = ~(layer_0[3206] ^ layer_0[3145]); 
    assign layer_1[1513] = layer_0[2744] ^ layer_0[2723]; 
    assign layer_1[1514] = ~(layer_0[1836] ^ layer_0[1894]); 
    assign layer_1[1515] = ~layer_0[228] | (layer_0[228] & layer_0[190]); 
    assign layer_1[1516] = layer_0[3216] & layer_0[3149]; 
    assign layer_1[1517] = layer_0[1650] & ~layer_0[1619]; 
    assign layer_1[1518] = layer_0[3318]; 
    assign layer_1[1519] = ~layer_0[3672]; 
    assign layer_1[1520] = ~(layer_0[3143] & layer_0[3119]); 
    assign layer_1[1521] = layer_0[3355] ^ layer_0[3378]; 
    assign layer_1[1522] = ~(layer_0[639] | layer_0[699]); 
    assign layer_1[1523] = layer_0[3090]; 
    assign layer_1[1524] = ~layer_0[2264]; 
    assign layer_1[1525] = ~(layer_0[924] ^ layer_0[1008]); 
    assign layer_1[1526] = ~(layer_0[2475] | layer_0[2367]); 
    assign layer_1[1527] = layer_0[20] & layer_0[68]; 
    assign layer_1[1528] = ~layer_0[1466]; 
    assign layer_1[1529] = layer_0[2261] | layer_0[2266]; 
    assign layer_1[1530] = ~layer_0[3921] | (layer_0[3921] & layer_0[3858]); 
    assign layer_1[1531] = layer_0[2381] & layer_0[2374]; 
    assign layer_1[1532] = layer_0[625] & layer_0[612]; 
    assign layer_1[1533] = layer_0[2123] & ~layer_0[2081]; 
    assign layer_1[1534] = layer_0[3967] ^ layer_0[3845]; 
    assign layer_1[1535] = layer_0[774] ^ layer_0[831]; 
    assign layer_1[1536] = layer_0[321]; 
    assign layer_1[1537] = ~layer_0[3890]; 
    assign layer_1[1538] = ~layer_0[1817]; 
    assign layer_1[1539] = layer_0[68] ^ layer_0[119]; 
    assign layer_1[1540] = layer_0[3362] | layer_0[3415]; 
    assign layer_1[1541] = ~layer_0[3458]; 
    assign layer_1[1542] = ~(layer_0[23] | layer_0[131]); 
    assign layer_1[1543] = layer_0[1657] & ~layer_0[1667]; 
    assign layer_1[1544] = layer_0[3987]; 
    assign layer_1[1545] = layer_0[948]; 
    assign layer_1[1546] = layer_0[2792] & ~layer_0[2882]; 
    assign layer_1[1547] = layer_0[1137] & ~layer_0[1069]; 
    assign layer_1[1548] = layer_0[1091] & ~layer_0[1197]; 
    assign layer_1[1549] = layer_0[44] & ~layer_0[165]; 
    assign layer_1[1550] = layer_0[1280] & ~layer_0[1338]; 
    assign layer_1[1551] = layer_0[1025] ^ layer_0[983]; 
    assign layer_1[1552] = ~layer_0[2305]; 
    assign layer_1[1553] = layer_0[3668] | layer_0[3552]; 
    assign layer_1[1554] = layer_0[1148]; 
    assign layer_1[1555] = layer_0[3436] & ~layer_0[3354]; 
    assign layer_1[1556] = ~layer_0[1230]; 
    assign layer_1[1557] = ~layer_0[3304] | (layer_0[3223] & layer_0[3304]); 
    assign layer_1[1558] = layer_0[2200] & ~layer_0[2184]; 
    assign layer_1[1559] = ~(layer_0[2182] ^ layer_0[2212]); 
    assign layer_1[1560] = ~(layer_0[1786] | layer_0[1697]); 
    assign layer_1[1561] = ~layer_0[1648]; 
    assign layer_1[1562] = ~(layer_0[44] ^ layer_0[153]); 
    assign layer_1[1563] = ~layer_0[1451]; 
    assign layer_1[1564] = layer_0[3497]; 
    assign layer_1[1565] = layer_0[1252]; 
    assign layer_1[1566] = ~(layer_0[1830] & layer_0[1946]); 
    assign layer_1[1567] = layer_0[2905] | layer_0[2830]; 
    assign layer_1[1568] = layer_0[3865] ^ layer_0[3760]; 
    assign layer_1[1569] = layer_0[2479] & layer_0[2480]; 
    assign layer_1[1570] = layer_0[2458] ^ layer_0[2546]; 
    assign layer_1[1571] = layer_0[3727] ^ layer_0[3778]; 
    assign layer_1[1572] = layer_0[3092]; 
    assign layer_1[1573] = ~layer_0[343]; 
    assign layer_1[1574] = ~layer_0[3009]; 
    assign layer_1[1575] = ~(layer_0[3916] | layer_0[3906]); 
    assign layer_1[1576] = ~(layer_0[496] ^ layer_0[572]); 
    assign layer_1[1577] = ~layer_0[1003]; 
    assign layer_1[1578] = layer_0[2700]; 
    assign layer_1[1579] = ~(layer_0[1208] | layer_0[1116]); 
    assign layer_1[1580] = ~(layer_0[3737] ^ layer_0[3743]); 
    assign layer_1[1581] = ~layer_0[1324]; 
    assign layer_1[1582] = layer_0[2090] & ~layer_0[2040]; 
    assign layer_1[1583] = layer_0[2475] ^ layer_0[2389]; 
    assign layer_1[1584] = ~layer_0[1825]; 
    assign layer_1[1585] = layer_0[1628]; 
    assign layer_1[1586] = layer_0[2294] & layer_0[2348]; 
    assign layer_1[1587] = layer_0[870] | layer_0[936]; 
    assign layer_1[1588] = layer_0[2459] & ~layer_0[2438]; 
    assign layer_1[1589] = layer_0[192] & ~layer_0[263]; 
    assign layer_1[1590] = layer_0[565]; 
    assign layer_1[1591] = layer_0[2369] ^ layer_0[2310]; 
    assign layer_1[1592] = layer_0[3441]; 
    assign layer_1[1593] = layer_0[2814]; 
    assign layer_1[1594] = ~(layer_0[2386] ^ layer_0[2453]); 
    assign layer_1[1595] = ~(layer_0[3995] | layer_0[3869]); 
    assign layer_1[1596] = ~(layer_0[1417] & layer_0[1363]); 
    assign layer_1[1597] = layer_0[1005] & ~layer_0[1024]; 
    assign layer_1[1598] = ~(layer_0[311] | layer_0[384]); 
    assign layer_1[1599] = ~layer_0[1709] | (layer_0[1610] & layer_0[1709]); 
    assign layer_1[1600] = layer_0[594] | layer_0[628]; 
    assign layer_1[1601] = ~layer_0[1265] | (layer_0[1316] & layer_0[1265]); 
    assign layer_1[1602] = layer_0[811] & ~layer_0[785]; 
    assign layer_1[1603] = ~layer_0[3444]; 
    assign layer_1[1604] = ~layer_0[164]; 
    assign layer_1[1605] = ~layer_0[1881]; 
    assign layer_1[1606] = layer_0[3231] & layer_0[3314]; 
    assign layer_1[1607] = layer_0[1863]; 
    assign layer_1[1608] = ~(layer_0[2251] ^ layer_0[2212]); 
    assign layer_1[1609] = layer_0[1028]; 
    assign layer_1[1610] = ~(layer_0[3834] | layer_0[3813]); 
    assign layer_1[1611] = ~(layer_0[3892] ^ layer_0[3816]); 
    assign layer_1[1612] = ~layer_0[2597]; 
    assign layer_1[1613] = ~layer_0[465] | (layer_0[475] & layer_0[465]); 
    assign layer_1[1614] = ~(layer_0[893] & layer_0[807]); 
    assign layer_1[1615] = layer_0[2609] & ~layer_0[2547]; 
    assign layer_1[1616] = layer_0[2824] | layer_0[2779]; 
    assign layer_1[1617] = ~(layer_0[716] ^ layer_0[843]); 
    assign layer_1[1618] = ~layer_0[751]; 
    assign layer_1[1619] = layer_0[2181] & ~layer_0[2200]; 
    assign layer_1[1620] = layer_0[3045] & layer_0[3006]; 
    assign layer_1[1621] = ~layer_0[3188]; 
    assign layer_1[1622] = ~layer_0[2058]; 
    assign layer_1[1623] = ~layer_0[2834]; 
    assign layer_1[1624] = ~(layer_0[2839] | layer_0[2951]); 
    assign layer_1[1625] = ~(layer_0[2296] & layer_0[2269]); 
    assign layer_1[1626] = layer_0[2974] & ~layer_0[2908]; 
    assign layer_1[1627] = layer_0[3865] ^ layer_0[3992]; 
    assign layer_1[1628] = layer_0[454]; 
    assign layer_1[1629] = layer_0[830]; 
    assign layer_1[1630] = layer_0[2844] ^ layer_0[2858]; 
    assign layer_1[1631] = ~layer_0[3724]; 
    assign layer_1[1632] = ~(layer_0[3456] ^ layer_0[3530]); 
    assign layer_1[1633] = ~layer_0[3501] | (layer_0[3512] & layer_0[3501]); 
    assign layer_1[1634] = ~(layer_0[1182] | layer_0[1266]); 
    assign layer_1[1635] = layer_0[1333]; 
    assign layer_1[1636] = ~(layer_0[3908] ^ layer_0[3992]); 
    assign layer_1[1637] = layer_0[1140] & layer_0[1014]; 
    assign layer_1[1638] = ~(layer_0[2288] ^ layer_0[2376]); 
    assign layer_1[1639] = layer_0[1602]; 
    assign layer_1[1640] = layer_0[2639] & ~layer_0[2695]; 
    assign layer_1[1641] = ~layer_0[3899] | (layer_0[3918] & layer_0[3899]); 
    assign layer_1[1642] = ~layer_0[3015]; 
    assign layer_1[1643] = ~(layer_0[3077] | layer_0[3041]); 
    assign layer_1[1644] = ~layer_0[285]; 
    assign layer_1[1645] = ~(layer_0[3089] & layer_0[3188]); 
    assign layer_1[1646] = layer_0[3774] & layer_0[3693]; 
    assign layer_1[1647] = ~layer_0[394] | (layer_0[394] & layer_0[313]); 
    assign layer_1[1648] = layer_0[1042] ^ layer_0[1068]; 
    assign layer_1[1649] = ~layer_0[1652]; 
    assign layer_1[1650] = ~(layer_0[1092] & layer_0[1039]); 
    assign layer_1[1651] = ~(layer_0[1843] | layer_0[1785]); 
    assign layer_1[1652] = layer_0[728] ^ layer_0[761]; 
    assign layer_1[1653] = layer_0[689] ^ layer_0[676]; 
    assign layer_1[1654] = ~layer_0[1902]; 
    assign layer_1[1655] = ~layer_0[2784] | (layer_0[2784] & layer_0[2891]); 
    assign layer_1[1656] = ~(layer_0[169] ^ layer_0[122]); 
    assign layer_1[1657] = layer_0[701] | layer_0[761]; 
    assign layer_1[1658] = layer_0[3940] & ~layer_0[3861]; 
    assign layer_1[1659] = ~layer_0[1059]; 
    assign layer_1[1660] = ~layer_0[2649] | (layer_0[2718] & layer_0[2649]); 
    assign layer_1[1661] = ~(layer_0[3274] ^ layer_0[3402]); 
    assign layer_1[1662] = layer_0[975]; 
    assign layer_1[1663] = layer_0[2903] & layer_0[2817]; 
    assign layer_1[1664] = ~layer_0[3908]; 
    assign layer_1[1665] = layer_0[2065] & ~layer_0[2144]; 
    assign layer_1[1666] = layer_0[2306] & layer_0[2372]; 
    assign layer_1[1667] = layer_0[1697] & ~layer_0[1666]; 
    assign layer_1[1668] = layer_0[1028] ^ layer_0[1042]; 
    assign layer_1[1669] = ~layer_0[3349] | (layer_0[3349] & layer_0[3256]); 
    assign layer_1[1670] = ~(layer_0[2325] | layer_0[2267]); 
    assign layer_1[1671] = ~layer_0[482]; 
    assign layer_1[1672] = ~(layer_0[1403] | layer_0[1461]); 
    assign layer_1[1673] = layer_0[2174]; 
    assign layer_1[1674] = layer_0[556] & ~layer_0[648]; 
    assign layer_1[1675] = layer_0[1010] & ~layer_0[1082]; 
    assign layer_1[1676] = layer_0[319] ^ layer_0[293]; 
    assign layer_1[1677] = ~layer_0[637]; 
    assign layer_1[1678] = layer_0[3296] & ~layer_0[3168]; 
    assign layer_1[1679] = layer_0[2414] ^ layer_0[2394]; 
    assign layer_1[1680] = layer_0[1826]; 
    assign layer_1[1681] = ~layer_0[736] | (layer_0[721] & layer_0[736]); 
    assign layer_1[1682] = layer_0[2351]; 
    assign layer_1[1683] = ~(layer_0[2116] ^ layer_0[2148]); 
    assign layer_1[1684] = layer_0[3776] & layer_0[3807]; 
    assign layer_1[1685] = layer_0[272]; 
    assign layer_1[1686] = ~(layer_0[638] & layer_0[675]); 
    assign layer_1[1687] = ~(layer_0[3181] ^ layer_0[3167]); 
    assign layer_1[1688] = layer_0[3659]; 
    assign layer_1[1689] = ~(layer_0[178] & layer_0[193]); 
    assign layer_1[1690] = ~layer_0[2178] | (layer_0[2178] & layer_0[2187]); 
    assign layer_1[1691] = ~(layer_0[1164] & layer_0[1235]); 
    assign layer_1[1692] = ~(layer_0[2109] & layer_0[1996]); 
    assign layer_1[1693] = layer_0[2171]; 
    assign layer_1[1694] = layer_0[3521]; 
    assign layer_1[1695] = ~(layer_0[1037] & layer_0[1021]); 
    assign layer_1[1696] = ~(layer_0[3292] ^ layer_0[3321]); 
    assign layer_1[1697] = layer_0[3778] & ~layer_0[3833]; 
    assign layer_1[1698] = layer_0[211] | layer_0[257]; 
    assign layer_1[1699] = ~(layer_0[2688] & layer_0[2745]); 
    assign layer_1[1700] = layer_0[2516] & ~layer_0[2442]; 
    assign layer_1[1701] = layer_0[383]; 
    assign layer_1[1702] = ~(layer_0[345] | layer_0[234]); 
    assign layer_1[1703] = ~layer_0[708] | (layer_0[693] & layer_0[708]); 
    assign layer_1[1704] = ~layer_0[3540]; 
    assign layer_1[1705] = layer_0[3240] & ~layer_0[3173]; 
    assign layer_1[1706] = ~(layer_0[1963] ^ layer_0[1888]); 
    assign layer_1[1707] = layer_0[2876] & ~layer_0[2825]; 
    assign layer_1[1708] = ~(layer_0[3093] & layer_0[3161]); 
    assign layer_1[1709] = ~(layer_0[1558] ^ layer_0[1609]); 
    assign layer_1[1710] = layer_0[931] ^ layer_0[1037]; 
    assign layer_1[1711] = ~layer_0[1179]; 
    assign layer_1[1712] = layer_0[1103] & layer_0[1005]; 
    assign layer_1[1713] = ~layer_0[3393]; 
    assign layer_1[1714] = layer_0[1598] & layer_0[1617]; 
    assign layer_1[1715] = ~layer_0[208]; 
    assign layer_1[1716] = layer_0[1207] ^ layer_0[1097]; 
    assign layer_1[1717] = layer_0[2346] ^ layer_0[2379]; 
    assign layer_1[1718] = ~(layer_0[769] | layer_0[747]); 
    assign layer_1[1719] = layer_0[496] & ~layer_0[481]; 
    assign layer_1[1720] = ~layer_0[1439] | (layer_0[1422] & layer_0[1439]); 
    assign layer_1[1721] = layer_0[3702] ^ layer_0[3767]; 
    assign layer_1[1722] = ~(layer_0[3453] ^ layer_0[3363]); 
    assign layer_1[1723] = layer_0[1021] & ~layer_0[1010]; 
    assign layer_1[1724] = layer_0[1690]; 
    assign layer_1[1725] = ~(layer_0[1263] ^ layer_0[1349]); 
    assign layer_1[1726] = layer_0[1799] & ~layer_0[1812]; 
    assign layer_1[1727] = ~(layer_0[3269] ^ layer_0[3396]); 
    assign layer_1[1728] = layer_0[285]; 
    assign layer_1[1729] = ~(layer_0[1397] ^ layer_0[1369]); 
    assign layer_1[1730] = layer_0[3016]; 
    assign layer_1[1731] = ~layer_0[625] | (layer_0[593] & layer_0[625]); 
    assign layer_1[1732] = layer_0[1705]; 
    assign layer_1[1733] = ~(layer_0[1123] | layer_0[1199]); 
    assign layer_1[1734] = layer_0[1694] & ~layer_0[1631]; 
    assign layer_1[1735] = ~(layer_0[219] & layer_0[253]); 
    assign layer_1[1736] = ~layer_0[2640] | (layer_0[2640] & layer_0[2672]); 
    assign layer_1[1737] = ~(layer_0[3972] ^ layer_0[3906]); 
    assign layer_1[1738] = ~(layer_0[1216] ^ layer_0[1300]); 
    assign layer_1[1739] = ~(layer_0[873] | layer_0[961]); 
    assign layer_1[1740] = ~layer_0[1533] | (layer_0[1533] & layer_0[1480]); 
    assign layer_1[1741] = ~layer_0[2900] | (layer_0[2900] & layer_0[2964]); 
    assign layer_1[1742] = ~(layer_0[2440] ^ layer_0[2315]); 
    assign layer_1[1743] = ~(layer_0[3648] & layer_0[3753]); 
    assign layer_1[1744] = layer_0[2943] & ~layer_0[2907]; 
    assign layer_1[1745] = ~layer_0[1841] | (layer_0[1899] & layer_0[1841]); 
    assign layer_1[1746] = layer_0[1964] & layer_0[2031]; 
    assign layer_1[1747] = ~layer_0[2013]; 
    assign layer_1[1748] = layer_0[1455] & ~layer_0[1358]; 
    assign layer_1[1749] = ~layer_0[556]; 
    assign layer_1[1750] = ~layer_0[303] | (layer_0[303] & layer_0[297]); 
    assign layer_1[1751] = ~layer_0[1481]; 
    assign layer_1[1752] = ~layer_0[516]; 
    assign layer_1[1753] = layer_0[3177] ^ layer_0[3267]; 
    assign layer_1[1754] = ~layer_0[1804]; 
    assign layer_1[1755] = ~layer_0[2928] | (layer_0[2928] & layer_0[2923]); 
    assign layer_1[1756] = layer_0[900]; 
    assign layer_1[1757] = ~(layer_0[1069] & layer_0[1012]); 
    assign layer_1[1758] = layer_0[974] & ~layer_0[981]; 
    assign layer_1[1759] = ~(layer_0[504] ^ layer_0[399]); 
    assign layer_1[1760] = layer_0[275] & ~layer_0[254]; 
    assign layer_1[1761] = layer_0[1056] & ~layer_0[1024]; 
    assign layer_1[1762] = layer_0[3553]; 
    assign layer_1[1763] = ~layer_0[289] | (layer_0[289] & layer_0[398]); 
    assign layer_1[1764] = layer_0[2029] & layer_0[2038]; 
    assign layer_1[1765] = layer_0[1557] & ~layer_0[1446]; 
    assign layer_1[1766] = layer_0[3125] & layer_0[3179]; 
    assign layer_1[1767] = ~(layer_0[1335] ^ layer_0[1347]); 
    assign layer_1[1768] = layer_0[1540] & layer_0[1473]; 
    assign layer_1[1769] = ~layer_0[2715]; 
    assign layer_1[1770] = ~layer_0[3992]; 
    assign layer_1[1771] = ~(layer_0[2975] & layer_0[2956]); 
    assign layer_1[1772] = ~(layer_0[3487] & layer_0[3412]); 
    assign layer_1[1773] = ~layer_0[1984]; 
    assign layer_1[1774] = ~(layer_0[2530] & layer_0[2442]); 
    assign layer_1[1775] = layer_0[2023] & layer_0[2087]; 
    assign layer_1[1776] = ~layer_0[423]; 
    assign layer_1[1777] = layer_0[2425] | layer_0[2418]; 
    assign layer_1[1778] = ~layer_0[2464] | (layer_0[2464] & layer_0[2546]); 
    assign layer_1[1779] = ~(layer_0[29] | layer_0[127]); 
    assign layer_1[1780] = ~layer_0[2191]; 
    assign layer_1[1781] = ~(layer_0[3868] ^ layer_0[3844]); 
    assign layer_1[1782] = layer_0[1406] & layer_0[1453]; 
    assign layer_1[1783] = layer_0[1384]; 
    assign layer_1[1784] = ~layer_0[2623]; 
    assign layer_1[1785] = ~layer_0[3533]; 
    assign layer_1[1786] = layer_0[2715] ^ layer_0[2651]; 
    assign layer_1[1787] = ~layer_0[2868] | (layer_0[2990] & layer_0[2868]); 
    assign layer_1[1788] = layer_0[3952] | layer_0[3863]; 
    assign layer_1[1789] = layer_0[2199] & ~layer_0[2299]; 
    assign layer_1[1790] = layer_0[3108] ^ layer_0[3016]; 
    assign layer_1[1791] = layer_0[1749]; 
    assign layer_1[1792] = layer_0[648]; 
    assign layer_1[1793] = layer_0[1736]; 
    assign layer_1[1794] = layer_0[434]; 
    assign layer_1[1795] = layer_0[97] & ~layer_0[164]; 
    assign layer_1[1796] = ~(layer_0[122] | layer_0[159]); 
    assign layer_1[1797] = ~layer_0[3692]; 
    assign layer_1[1798] = ~(layer_0[3832] | layer_0[3782]); 
    assign layer_1[1799] = ~layer_0[3636] | (layer_0[3674] & layer_0[3636]); 
    assign layer_1[1800] = ~(layer_0[3878] & layer_0[3966]); 
    assign layer_1[1801] = layer_0[1624] & layer_0[1602]; 
    assign layer_1[1802] = ~layer_0[1691] | (layer_0[1748] & layer_0[1691]); 
    assign layer_1[1803] = layer_0[2512] ^ layer_0[2573]; 
    assign layer_1[1804] = layer_0[3713] & ~layer_0[3603]; 
    assign layer_1[1805] = ~layer_0[2262] | (layer_0[2270] & layer_0[2262]); 
    assign layer_1[1806] = ~layer_0[1586]; 
    assign layer_1[1807] = layer_0[2718] & ~layer_0[2629]; 
    assign layer_1[1808] = ~(layer_0[2620] ^ layer_0[2604]); 
    assign layer_1[1809] = layer_0[3696] | layer_0[3703]; 
    assign layer_1[1810] = ~(layer_0[315] & layer_0[372]); 
    assign layer_1[1811] = ~(layer_0[911] ^ layer_0[943]); 
    assign layer_1[1812] = layer_0[1347] ^ layer_0[1471]; 
    assign layer_1[1813] = layer_0[2575] & ~layer_0[2616]; 
    assign layer_1[1814] = ~(layer_0[48] ^ layer_0[147]); 
    assign layer_1[1815] = layer_0[1045] & layer_0[1040]; 
    assign layer_1[1816] = ~layer_0[2614]; 
    assign layer_1[1817] = ~(layer_0[1922] | layer_0[1989]); 
    assign layer_1[1818] = ~layer_0[3254] | (layer_0[3141] & layer_0[3254]); 
    assign layer_1[1819] = layer_0[1531] & ~layer_0[1504]; 
    assign layer_1[1820] = layer_0[691] & ~layer_0[696]; 
    assign layer_1[1821] = ~(layer_0[1230] ^ layer_0[1124]); 
    assign layer_1[1822] = layer_0[458]; 
    assign layer_1[1823] = ~layer_0[2436]; 
    assign layer_1[1824] = ~layer_0[1422]; 
    assign layer_1[1825] = ~(layer_0[1175] | layer_0[1181]); 
    assign layer_1[1826] = layer_0[320]; 
    assign layer_1[1827] = ~(layer_0[1610] ^ layer_0[1499]); 
    assign layer_1[1828] = ~(layer_0[3456] & layer_0[3391]); 
    assign layer_1[1829] = layer_0[2112] | layer_0[2074]; 
    assign layer_1[1830] = layer_0[3757] & ~layer_0[3694]; 
    assign layer_1[1831] = layer_0[940]; 
    assign layer_1[1832] = layer_0[2271] & ~layer_0[2246]; 
    assign layer_1[1833] = ~(layer_0[982] | layer_0[896]); 
    assign layer_1[1834] = ~layer_0[2148]; 
    assign layer_1[1835] = layer_0[3159] & ~layer_0[3248]; 
    assign layer_1[1836] = ~(layer_0[3548] ^ layer_0[3541]); 
    assign layer_1[1837] = ~(layer_0[1093] ^ layer_0[1034]); 
    assign layer_1[1838] = ~layer_0[3423]; 
    assign layer_1[1839] = ~(layer_0[1322] ^ layer_0[1360]); 
    assign layer_1[1840] = ~(layer_0[1279] & layer_0[1278]); 
    assign layer_1[1841] = layer_0[419] & ~layer_0[475]; 
    assign layer_1[1842] = ~layer_0[3945] | (layer_0[3945] & layer_0[3993]); 
    assign layer_1[1843] = ~(layer_0[842] & layer_0[946]); 
    assign layer_1[1844] = layer_0[923] & layer_0[921]; 
    assign layer_1[1845] = layer_0[1130] ^ layer_0[1120]; 
    assign layer_1[1846] = ~(layer_0[2670] | layer_0[2623]); 
    assign layer_1[1847] = layer_0[2675] ^ layer_0[2673]; 
    assign layer_1[1848] = ~layer_0[2706] | (layer_0[2815] & layer_0[2706]); 
    assign layer_1[1849] = ~(layer_0[1786] & layer_0[1868]); 
    assign layer_1[1850] = ~(layer_0[1757] & layer_0[1647]); 
    assign layer_1[1851] = ~(layer_0[1867] & layer_0[1925]); 
    assign layer_1[1852] = layer_0[2810]; 
    assign layer_1[1853] = ~(layer_0[1214] & layer_0[1284]); 
    assign layer_1[1854] = ~layer_0[1223] | (layer_0[1223] & layer_0[1113]); 
    assign layer_1[1855] = layer_0[3176]; 
    assign layer_1[1856] = ~layer_0[1869] | (layer_0[1869] & layer_0[1951]); 
    assign layer_1[1857] = ~layer_0[3952] | (layer_0[3992] & layer_0[3952]); 
    assign layer_1[1858] = ~layer_0[1311]; 
    assign layer_1[1859] = layer_0[1930] & ~layer_0[1971]; 
    assign layer_1[1860] = layer_0[2111] ^ layer_0[2130]; 
    assign layer_1[1861] = ~layer_0[1034] | (layer_0[1017] & layer_0[1034]); 
    assign layer_1[1862] = layer_0[2800]; 
    assign layer_1[1863] = layer_0[1473]; 
    assign layer_1[1864] = layer_0[1397] ^ layer_0[1396]; 
    assign layer_1[1865] = ~layer_0[2432]; 
    assign layer_1[1866] = layer_0[3186]; 
    assign layer_1[1867] = ~layer_0[3546]; 
    assign layer_1[1868] = layer_0[3036] ^ layer_0[3065]; 
    assign layer_1[1869] = ~(layer_0[2708] ^ layer_0[2634]); 
    assign layer_1[1870] = ~(layer_0[1097] ^ layer_0[1220]); 
    assign layer_1[1871] = ~(layer_0[289] ^ layer_0[412]); 
    assign layer_1[1872] = ~(layer_0[1786] & layer_0[1849]); 
    assign layer_1[1873] = layer_0[1679] & ~layer_0[1556]; 
    assign layer_1[1874] = layer_0[2952] & ~layer_0[3024]; 
    assign layer_1[1875] = ~layer_0[298] | (layer_0[298] & layer_0[281]); 
    assign layer_1[1876] = layer_0[799] | layer_0[698]; 
    assign layer_1[1877] = layer_0[1040] & ~layer_0[1063]; 
    assign layer_1[1878] = ~layer_0[1479] | (layer_0[1479] & layer_0[1572]); 
    assign layer_1[1879] = layer_0[2508] & ~layer_0[2445]; 
    assign layer_1[1880] = layer_0[2879]; 
    assign layer_1[1881] = layer_0[205] ^ layer_0[81]; 
    assign layer_1[1882] = ~(layer_0[1374] ^ layer_0[1277]); 
    assign layer_1[1883] = layer_0[2516] | layer_0[2424]; 
    assign layer_1[1884] = layer_0[2690] & ~layer_0[2764]; 
    assign layer_1[1885] = ~layer_0[3506] | (layer_0[3594] & layer_0[3506]); 
    assign layer_1[1886] = layer_0[1606] & ~layer_0[1658]; 
    assign layer_1[1887] = ~layer_0[3584] | (layer_0[3554] & layer_0[3584]); 
    assign layer_1[1888] = ~layer_0[3826]; 
    assign layer_1[1889] = layer_0[755] & ~layer_0[709]; 
    assign layer_1[1890] = layer_0[3128] & ~layer_0[3023]; 
    assign layer_1[1891] = layer_0[2567] ^ layer_0[2655]; 
    assign layer_1[1892] = ~(layer_0[3876] ^ layer_0[3855]); 
    assign layer_1[1893] = layer_0[2310] ^ layer_0[2380]; 
    assign layer_1[1894] = layer_0[537] ^ layer_0[488]; 
    assign layer_1[1895] = layer_0[56] & layer_0[158]; 
    assign layer_1[1896] = layer_0[1737] | layer_0[1839]; 
    assign layer_1[1897] = ~(layer_0[2176] ^ layer_0[2240]); 
    assign layer_1[1898] = layer_0[2945] | layer_0[2819]; 
    assign layer_1[1899] = ~(layer_0[921] ^ layer_0[1043]); 
    assign layer_1[1900] = ~layer_0[1591]; 
    assign layer_1[1901] = ~layer_0[2512]; 
    assign layer_1[1902] = layer_0[2203] & ~layer_0[2254]; 
    assign layer_1[1903] = ~layer_0[3730]; 
    assign layer_1[1904] = ~(layer_0[2114] ^ layer_0[2228]); 
    assign layer_1[1905] = layer_0[2127] & layer_0[2110]; 
    assign layer_1[1906] = ~layer_0[1988] | (layer_0[1886] & layer_0[1988]); 
    assign layer_1[1907] = layer_0[295] & layer_0[251]; 
    assign layer_1[1908] = ~layer_0[2102] | (layer_0[2102] & layer_0[2214]); 
    assign layer_1[1909] = ~(layer_0[1731] ^ layer_0[1694]); 
    assign layer_1[1910] = layer_0[2371] & layer_0[2320]; 
    assign layer_1[1911] = ~layer_0[1627]; 
    assign layer_1[1912] = ~(layer_0[1568] | layer_0[1491]); 
    assign layer_1[1913] = layer_0[3255] | layer_0[3324]; 
    assign layer_1[1914] = ~layer_0[2073] | (layer_0[2073] & layer_0[2198]); 
    assign layer_1[1915] = ~layer_0[2927]; 
    assign layer_1[1916] = ~(layer_0[2158] & layer_0[2104]); 
    assign layer_1[1917] = ~(layer_0[3471] & layer_0[3422]); 
    assign layer_1[1918] = ~layer_0[775] | (layer_0[872] & layer_0[775]); 
    assign layer_1[1919] = layer_0[2165] & ~layer_0[2091]; 
    assign layer_1[1920] = ~layer_0[1561]; 
    assign layer_1[1921] = layer_0[563] & layer_0[450]; 
    assign layer_1[1922] = ~layer_0[2047]; 
    assign layer_1[1923] = ~(layer_0[3771] ^ layer_0[3662]); 
    assign layer_1[1924] = layer_0[1203] & layer_0[1320]; 
    assign layer_1[1925] = ~layer_0[1784]; 
    assign layer_1[1926] = ~(layer_0[3724] ^ layer_0[3783]); 
    assign layer_1[1927] = ~layer_0[222]; 
    assign layer_1[1928] = ~layer_0[2452]; 
    assign layer_1[1929] = layer_0[2619] & layer_0[2691]; 
    assign layer_1[1930] = ~layer_0[795] | (layer_0[704] & layer_0[795]); 
    assign layer_1[1931] = layer_0[2422]; 
    assign layer_1[1932] = ~layer_0[1545] | (layer_0[1501] & layer_0[1545]); 
    assign layer_1[1933] = ~(layer_0[3697] ^ layer_0[3666]); 
    assign layer_1[1934] = layer_0[364]; 
    assign layer_1[1935] = ~(layer_0[2798] | layer_0[2693]); 
    assign layer_1[1936] = ~layer_0[1856] | (layer_0[1856] & layer_0[1746]); 
    assign layer_1[1937] = layer_0[72] & ~layer_0[193]; 
    assign layer_1[1938] = layer_0[3053]; 
    assign layer_1[1939] = layer_0[49] & ~layer_0[137]; 
    assign layer_1[1940] = ~(layer_0[3422] & layer_0[3379]); 
    assign layer_1[1941] = layer_0[2493] & ~layer_0[2571]; 
    assign layer_1[1942] = layer_0[3345] & layer_0[3447]; 
    assign layer_1[1943] = ~(layer_0[3724] ^ layer_0[3664]); 
    assign layer_1[1944] = ~layer_0[1271] | (layer_0[1271] & layer_0[1278]); 
    assign layer_1[1945] = ~(layer_0[3088] ^ layer_0[3005]); 
    assign layer_1[1946] = ~layer_0[752]; 
    assign layer_1[1947] = layer_0[3805] & layer_0[3722]; 
    assign layer_1[1948] = layer_0[2680] & ~layer_0[2716]; 
    assign layer_1[1949] = layer_0[3157] ^ layer_0[3121]; 
    assign layer_1[1950] = ~(layer_0[2291] ^ layer_0[2194]); 
    assign layer_1[1951] = ~layer_0[650]; 
    assign layer_1[1952] = ~(layer_0[1606] ^ layer_0[1616]); 
    assign layer_1[1953] = layer_0[2770] ^ layer_0[2721]; 
    assign layer_1[1954] = ~layer_0[2064]; 
    assign layer_1[1955] = layer_0[1650]; 
    assign layer_1[1956] = layer_0[240] & layer_0[246]; 
    assign layer_1[1957] = layer_0[1272]; 
    assign layer_1[1958] = layer_0[143]; 
    assign layer_1[1959] = ~(layer_0[3948] ^ layer_0[3973]); 
    assign layer_1[1960] = ~layer_0[238]; 
    assign layer_1[1961] = ~layer_0[1027] | (layer_0[1147] & layer_0[1027]); 
    assign layer_1[1962] = ~layer_0[1867]; 
    assign layer_1[1963] = ~(layer_0[934] ^ layer_0[888]); 
    assign layer_1[1964] = ~(layer_0[1525] & layer_0[1409]); 
    assign layer_1[1965] = layer_0[3864]; 
    assign layer_1[1966] = layer_0[2754]; 
    assign layer_1[1967] = ~(layer_0[1800] & layer_0[1809]); 
    assign layer_1[1968] = ~layer_0[308] | (layer_0[222] & layer_0[308]); 
    assign layer_1[1969] = ~(layer_0[1321] ^ layer_0[1423]); 
    assign layer_1[1970] = ~(layer_0[890] | layer_0[999]); 
    assign layer_1[1971] = layer_0[2109] & ~layer_0[2199]; 
    assign layer_1[1972] = layer_0[597] & layer_0[690]; 
    assign layer_1[1973] = layer_0[339] & ~layer_0[267]; 
    assign layer_1[1974] = ~layer_0[688]; 
    assign layer_1[1975] = layer_0[1740] & ~layer_0[1733]; 
    assign layer_1[1976] = layer_0[1394]; 
    assign layer_1[1977] = ~(layer_0[3792] & layer_0[3688]); 
    assign layer_1[1978] = ~layer_0[3653]; 
    assign layer_1[1979] = ~(layer_0[3806] ^ layer_0[3741]); 
    assign layer_1[1980] = layer_0[1558] ^ layer_0[1562]; 
    assign layer_1[1981] = layer_0[1945] ^ layer_0[1824]; 
    assign layer_1[1982] = layer_0[3888]; 
    assign layer_1[1983] = layer_0[3633] ^ layer_0[3538]; 
    assign layer_1[1984] = layer_0[1592] | layer_0[1476]; 
    assign layer_1[1985] = layer_0[2814] & ~layer_0[2842]; 
    assign layer_1[1986] = layer_0[3903] & ~layer_0[3963]; 
    assign layer_1[1987] = ~(layer_0[3629] ^ layer_0[3723]); 
    assign layer_1[1988] = layer_0[1771] | layer_0[1860]; 
    assign layer_1[1989] = layer_0[820] & layer_0[800]; 
    assign layer_1[1990] = layer_0[758]; 
    assign layer_1[1991] = ~(layer_0[64] | layer_0[7]); 
    assign layer_1[1992] = layer_0[2412] | layer_0[2358]; 
    assign layer_1[1993] = layer_0[1653]; 
    assign layer_1[1994] = ~(layer_0[3921] | layer_0[3906]); 
    assign layer_1[1995] = layer_0[1446] ^ layer_0[1560]; 
    assign layer_1[1996] = ~layer_0[2647]; 
    assign layer_1[1997] = ~layer_0[505]; 
    assign layer_1[1998] = layer_0[3669]; 
    assign layer_1[1999] = layer_0[356]; 
    assign layer_1[2000] = layer_0[2560] & ~layer_0[2452]; 
    assign layer_1[2001] = layer_0[3603] & ~layer_0[3636]; 
    assign layer_1[2002] = ~layer_0[3601]; 
    assign layer_1[2003] = layer_0[3337] ^ layer_0[3210]; 
    assign layer_1[2004] = ~layer_0[2054]; 
    assign layer_1[2005] = layer_0[125]; 
    assign layer_1[2006] = ~(layer_0[185] & layer_0[303]); 
    assign layer_1[2007] = ~(layer_0[3527] ^ layer_0[3450]); 
    assign layer_1[2008] = layer_0[1456] & ~layer_0[1583]; 
    assign layer_1[2009] = ~layer_0[2651] | (layer_0[2651] & layer_0[2633]); 
    assign layer_1[2010] = layer_0[3962] | layer_0[3992]; 
    assign layer_1[2011] = layer_0[569]; 
    assign layer_1[2012] = layer_0[512] ^ layer_0[579]; 
    assign layer_1[2013] = ~layer_0[3137] | (layer_0[3129] & layer_0[3137]); 
    assign layer_1[2014] = layer_0[1969] & ~layer_0[2021]; 
    assign layer_1[2015] = ~layer_0[2705]; 
    assign layer_1[2016] = layer_0[672]; 
    assign layer_1[2017] = ~layer_0[2046]; 
    assign layer_1[2018] = layer_0[2545] & layer_0[2523]; 
    assign layer_1[2019] = layer_0[2324] & ~layer_0[2348]; 
    assign layer_1[2020] = layer_0[1343] & layer_0[1260]; 
    assign layer_1[2021] = ~layer_0[1171] | (layer_0[1116] & layer_0[1171]); 
    assign layer_1[2022] = layer_0[2692] & layer_0[2727]; 
    assign layer_1[2023] = layer_0[3019] ^ layer_0[3036]; 
    assign layer_1[2024] = layer_0[2919] & ~layer_0[3041]; 
    assign layer_1[2025] = layer_0[853] ^ layer_0[862]; 
    assign layer_1[2026] = ~layer_0[3172] | (layer_0[3246] & layer_0[3172]); 
    assign layer_1[2027] = ~(layer_0[174] ^ layer_0[79]); 
    assign layer_1[2028] = ~layer_0[1506] | (layer_0[1470] & layer_0[1506]); 
    assign layer_1[2029] = ~(layer_0[1613] | layer_0[1490]); 
    assign layer_1[2030] = layer_0[2857]; 
    assign layer_1[2031] = layer_0[2323] | layer_0[2325]; 
    assign layer_1[2032] = layer_0[3738]; 
    assign layer_1[2033] = layer_0[2569] & ~layer_0[2648]; 
    assign layer_1[2034] = ~(layer_0[848] ^ layer_0[793]); 
    assign layer_1[2035] = layer_0[1514] & layer_0[1581]; 
    assign layer_1[2036] = layer_0[3661] ^ layer_0[3762]; 
    assign layer_1[2037] = layer_0[2983] | layer_0[3097]; 
    assign layer_1[2038] = ~layer_0[3370] | (layer_0[3370] & layer_0[3301]); 
    assign layer_1[2039] = layer_0[3732] | layer_0[3769]; 
    assign layer_1[2040] = ~layer_0[187]; 
    assign layer_1[2041] = layer_0[3000]; 
    assign layer_1[2042] = layer_0[1509] ^ layer_0[1489]; 
    assign layer_1[2043] = ~layer_0[3196]; 
    assign layer_1[2044] = ~(layer_0[1124] & layer_0[1060]); 
    assign layer_1[2045] = ~(layer_0[774] & layer_0[803]); 
    assign layer_1[2046] = ~(layer_0[117] & layer_0[166]); 
    assign layer_1[2047] = ~(layer_0[1416] ^ layer_0[1508]); 
    assign layer_1[2048] = layer_0[1545] & ~layer_0[1496]; 
    assign layer_1[2049] = ~layer_0[3421]; 
    assign layer_1[2050] = layer_0[1956] | layer_0[1883]; 
    assign layer_1[2051] = ~layer_0[114]; 
    assign layer_1[2052] = ~layer_0[3970] | (layer_0[3953] & layer_0[3970]); 
    assign layer_1[2053] = ~layer_0[1053] | (layer_0[1053] & layer_0[1112]); 
    assign layer_1[2054] = layer_0[3639] | layer_0[3572]; 
    assign layer_1[2055] = layer_0[3337] & ~layer_0[3307]; 
    assign layer_1[2056] = ~layer_0[1511]; 
    assign layer_1[2057] = layer_0[3894] & ~layer_0[3798]; 
    assign layer_1[2058] = ~(layer_0[3987] ^ layer_0[3913]); 
    assign layer_1[2059] = ~layer_0[397]; 
    assign layer_1[2060] = ~(layer_0[3199] & layer_0[3294]); 
    assign layer_1[2061] = layer_0[3100]; 
    assign layer_1[2062] = layer_0[3521]; 
    assign layer_1[2063] = layer_0[236]; 
    assign layer_1[2064] = ~layer_0[241]; 
    assign layer_1[2065] = layer_0[2351]; 
    assign layer_1[2066] = layer_0[258]; 
    assign layer_1[2067] = layer_0[1949] & ~layer_0[1964]; 
    assign layer_1[2068] = layer_0[3646]; 
    assign layer_1[2069] = layer_0[1580] & layer_0[1548]; 
    assign layer_1[2070] = ~(layer_0[183] ^ layer_0[114]); 
    assign layer_1[2071] = layer_0[681] ^ layer_0[614]; 
    assign layer_1[2072] = ~layer_0[848]; 
    assign layer_1[2073] = ~(layer_0[1273] | layer_0[1376]); 
    assign layer_1[2074] = layer_0[2843] & ~layer_0[2824]; 
    assign layer_1[2075] = layer_0[1300] | layer_0[1377]; 
    assign layer_1[2076] = layer_0[1844] & ~layer_0[1788]; 
    assign layer_1[2077] = layer_0[2357]; 
    assign layer_1[2078] = ~(layer_0[1980] ^ layer_0[1942]); 
    assign layer_1[2079] = layer_0[1774] | layer_0[1830]; 
    assign layer_1[2080] = ~layer_0[2890]; 
    assign layer_1[2081] = ~(layer_0[446] & layer_0[364]); 
    assign layer_1[2082] = layer_0[2807]; 
    assign layer_1[2083] = layer_0[2640] ^ layer_0[2557]; 
    assign layer_1[2084] = ~(layer_0[1747] ^ layer_0[1818]); 
    assign layer_1[2085] = layer_0[3977] & ~layer_0[3997]; 
    assign layer_1[2086] = layer_0[1510] & layer_0[1505]; 
    assign layer_1[2087] = layer_0[3912] & ~layer_0[3943]; 
    assign layer_1[2088] = ~layer_0[3890]; 
    assign layer_1[2089] = layer_0[399]; 
    assign layer_1[2090] = layer_0[446] | layer_0[359]; 
    assign layer_1[2091] = ~layer_0[1183]; 
    assign layer_1[2092] = layer_0[3375]; 
    assign layer_1[2093] = ~(layer_0[107] & layer_0[163]); 
    assign layer_1[2094] = ~layer_0[119]; 
    assign layer_1[2095] = ~(layer_0[178] | layer_0[105]); 
    assign layer_1[2096] = layer_0[1989] & ~layer_0[1912]; 
    assign layer_1[2097] = layer_0[3467] & ~layer_0[3474]; 
    assign layer_1[2098] = layer_0[1905] ^ layer_0[1895]; 
    assign layer_1[2099] = layer_0[1820] ^ layer_0[1862]; 
    assign layer_1[2100] = layer_0[3101] ^ layer_0[3128]; 
    assign layer_1[2101] = layer_0[690]; 
    assign layer_1[2102] = layer_0[1034]; 
    assign layer_1[2103] = ~layer_0[503]; 
    assign layer_1[2104] = ~(layer_0[1717] ^ layer_0[1631]); 
    assign layer_1[2105] = layer_0[409] ^ layer_0[358]; 
    assign layer_1[2106] = layer_0[922] & ~layer_0[920]; 
    assign layer_1[2107] = ~(layer_0[499] & layer_0[538]); 
    assign layer_1[2108] = layer_0[1802]; 
    assign layer_1[2109] = ~layer_0[1612] | (layer_0[1528] & layer_0[1612]); 
    assign layer_1[2110] = ~layer_0[3286] | (layer_0[3286] & layer_0[3176]); 
    assign layer_1[2111] = layer_0[3307] ^ layer_0[3217]; 
    assign layer_1[2112] = ~(layer_0[1781] ^ layer_0[1807]); 
    assign layer_1[2113] = ~(layer_0[371] | layer_0[249]); 
    assign layer_1[2114] = layer_0[3587] & layer_0[3649]; 
    assign layer_1[2115] = ~layer_0[3068]; 
    assign layer_1[2116] = layer_0[2705]; 
    assign layer_1[2117] = layer_0[774] & ~layer_0[790]; 
    assign layer_1[2118] = layer_0[2644] ^ layer_0[2530]; 
    assign layer_1[2119] = layer_0[1513]; 
    assign layer_1[2120] = layer_0[1410] | layer_0[1338]; 
    assign layer_1[2121] = ~layer_0[2497] | (layer_0[2517] & layer_0[2497]); 
    assign layer_1[2122] = ~layer_0[1969] | (layer_0[1969] & layer_0[2020]); 
    assign layer_1[2123] = ~(layer_0[2028] & layer_0[1906]); 
    assign layer_1[2124] = layer_0[158]; 
    assign layer_1[2125] = layer_0[718]; 
    assign layer_1[2126] = ~(layer_0[775] ^ layer_0[772]); 
    assign layer_1[2127] = layer_0[1671]; 
    assign layer_1[2128] = ~(layer_0[932] | layer_0[806]); 
    assign layer_1[2129] = ~layer_0[3178]; 
    assign layer_1[2130] = ~(layer_0[737] ^ layer_0[864]); 
    assign layer_1[2131] = ~layer_0[2243]; 
    assign layer_1[2132] = layer_0[3604] | layer_0[3592]; 
    assign layer_1[2133] = ~layer_0[3621]; 
    assign layer_1[2134] = layer_0[510] & ~layer_0[487]; 
    assign layer_1[2135] = ~layer_0[775]; 
    assign layer_1[2136] = ~layer_0[3523]; 
    assign layer_1[2137] = ~(layer_0[2654] & layer_0[2572]); 
    assign layer_1[2138] = layer_0[1539] & layer_0[1612]; 
    assign layer_1[2139] = layer_0[1357] | layer_0[1445]; 
    assign layer_1[2140] = ~layer_0[2416] | (layer_0[2328] & layer_0[2416]); 
    assign layer_1[2141] = layer_0[370] | layer_0[279]; 
    assign layer_1[2142] = ~layer_0[2245]; 
    assign layer_1[2143] = ~layer_0[1666]; 
    assign layer_1[2144] = layer_0[2883]; 
    assign layer_1[2145] = ~(layer_0[3749] ^ layer_0[3765]); 
    assign layer_1[2146] = layer_0[1375] | layer_0[1390]; 
    assign layer_1[2147] = layer_0[3618] & ~layer_0[3564]; 
    assign layer_1[2148] = layer_0[2694] | layer_0[2646]; 
    assign layer_1[2149] = ~(layer_0[3981] & layer_0[3948]); 
    assign layer_1[2150] = layer_0[3398]; 
    assign layer_1[2151] = layer_0[355] ^ layer_0[426]; 
    assign layer_1[2152] = layer_0[494] & ~layer_0[386]; 
    assign layer_1[2153] = layer_0[2813] ^ layer_0[2850]; 
    assign layer_1[2154] = ~layer_0[2205]; 
    assign layer_1[2155] = ~(layer_0[2146] ^ layer_0[2252]); 
    assign layer_1[2156] = ~(layer_0[682] | layer_0[643]); 
    assign layer_1[2157] = layer_0[3336] ^ layer_0[3348]; 
    assign layer_1[2158] = ~(layer_0[1450] | layer_0[1361]); 
    assign layer_1[2159] = layer_0[2726] ^ layer_0[2851]; 
    assign layer_1[2160] = ~layer_0[1599]; 
    assign layer_1[2161] = ~layer_0[659] | (layer_0[659] & layer_0[567]); 
    assign layer_1[2162] = ~(layer_0[2352] & layer_0[2437]); 
    assign layer_1[2163] = layer_0[1684] & ~layer_0[1724]; 
    assign layer_1[2164] = ~layer_0[3407]; 
    assign layer_1[2165] = ~layer_0[2510]; 
    assign layer_1[2166] = layer_0[385] & ~layer_0[475]; 
    assign layer_1[2167] = ~(layer_0[1552] & layer_0[1620]); 
    assign layer_1[2168] = layer_0[638]; 
    assign layer_1[2169] = layer_0[1942] & ~layer_0[1932]; 
    assign layer_1[2170] = ~(layer_0[863] ^ layer_0[864]); 
    assign layer_1[2171] = layer_0[1354]; 
    assign layer_1[2172] = layer_0[1848] | layer_0[1961]; 
    assign layer_1[2173] = layer_0[3343] ^ layer_0[3368]; 
    assign layer_1[2174] = ~(layer_0[2445] ^ layer_0[2451]); 
    assign layer_1[2175] = layer_0[2132] & layer_0[2123]; 
    assign layer_1[2176] = layer_0[2012] ^ layer_0[2070]; 
    assign layer_1[2177] = ~(layer_0[3406] & layer_0[3361]); 
    assign layer_1[2178] = ~layer_0[3490] | (layer_0[3391] & layer_0[3490]); 
    assign layer_1[2179] = layer_0[843] & layer_0[965]; 
    assign layer_1[2180] = layer_0[3925] ^ layer_0[3889]; 
    assign layer_1[2181] = layer_0[3807] & layer_0[3866]; 
    assign layer_1[2182] = ~layer_0[701]; 
    assign layer_1[2183] = ~layer_0[1198]; 
    assign layer_1[2184] = layer_0[2982] & layer_0[2989]; 
    assign layer_1[2185] = layer_0[954] & ~layer_0[903]; 
    assign layer_1[2186] = ~(layer_0[1282] | layer_0[1402]); 
    assign layer_1[2187] = ~(layer_0[2302] | layer_0[2287]); 
    assign layer_1[2188] = layer_0[575] | layer_0[539]; 
    assign layer_1[2189] = layer_0[2705] & ~layer_0[2649]; 
    assign layer_1[2190] = ~layer_0[601] | (layer_0[726] & layer_0[601]); 
    assign layer_1[2191] = ~(layer_0[2101] ^ layer_0[2014]); 
    assign layer_1[2192] = layer_0[950]; 
    assign layer_1[2193] = layer_0[1470] & ~layer_0[1374]; 
    assign layer_1[2194] = ~layer_0[2081]; 
    assign layer_1[2195] = layer_0[3953] | layer_0[3967]; 
    assign layer_1[2196] = layer_0[756] | layer_0[801]; 
    assign layer_1[2197] = ~layer_0[3070] | (layer_0[3070] & layer_0[3114]); 
    assign layer_1[2198] = layer_0[3866]; 
    assign layer_1[2199] = ~(layer_0[3004] | layer_0[2923]); 
    assign layer_1[2200] = layer_0[2711]; 
    assign layer_1[2201] = ~layer_0[768]; 
    assign layer_1[2202] = ~layer_0[320] | (layer_0[320] & layer_0[377]); 
    assign layer_1[2203] = layer_0[410] & ~layer_0[359]; 
    assign layer_1[2204] = layer_0[14] & ~layer_0[48]; 
    assign layer_1[2205] = layer_0[3506] & ~layer_0[3416]; 
    assign layer_1[2206] = ~layer_0[3858] | (layer_0[3858] & layer_0[3828]); 
    assign layer_1[2207] = ~layer_0[716]; 
    assign layer_1[2208] = layer_0[865] & layer_0[764]; 
    assign layer_1[2209] = layer_0[2160]; 
    assign layer_1[2210] = ~layer_0[2349]; 
    assign layer_1[2211] = ~layer_0[2101] | (layer_0[2101] & layer_0[2040]); 
    assign layer_1[2212] = layer_0[112] | layer_0[146]; 
    assign layer_1[2213] = ~(layer_0[2862] ^ layer_0[2879]); 
    assign layer_1[2214] = layer_0[1891]; 
    assign layer_1[2215] = ~layer_0[1274]; 
    assign layer_1[2216] = layer_0[86]; 
    assign layer_1[2217] = ~layer_0[2199]; 
    assign layer_1[2218] = layer_0[3983] | layer_0[3994]; 
    assign layer_1[2219] = layer_0[1940] & ~layer_0[1929]; 
    assign layer_1[2220] = ~layer_0[35]; 
    assign layer_1[2221] = layer_0[173] & ~layer_0[281]; 
    assign layer_1[2222] = layer_0[3689] | layer_0[3634]; 
    assign layer_1[2223] = layer_0[1773]; 
    assign layer_1[2224] = ~(layer_0[975] ^ layer_0[1017]); 
    assign layer_1[2225] = ~layer_0[27] | (layer_0[20] & layer_0[27]); 
    assign layer_1[2226] = layer_0[3544]; 
    assign layer_1[2227] = layer_0[1579] ^ layer_0[1628]; 
    assign layer_1[2228] = ~(layer_0[3472] | layer_0[3585]); 
    assign layer_1[2229] = layer_0[134] & ~layer_0[20]; 
    assign layer_1[2230] = layer_0[33] & ~layer_0[82]; 
    assign layer_1[2231] = ~layer_0[2498] | (layer_0[2498] & layer_0[2414]); 
    assign layer_1[2232] = layer_0[3491] & layer_0[3405]; 
    assign layer_1[2233] = ~layer_0[2742]; 
    assign layer_1[2234] = layer_0[683] & layer_0[640]; 
    assign layer_1[2235] = ~(layer_0[38] | layer_0[91]); 
    assign layer_1[2236] = layer_0[1948]; 
    assign layer_1[2237] = ~(layer_0[3856] & layer_0[3764]); 
    assign layer_1[2238] = ~(layer_0[1693] & layer_0[1773]); 
    assign layer_1[2239] = ~layer_0[3611]; 
    assign layer_1[2240] = layer_0[1791]; 
    assign layer_1[2241] = ~(layer_0[96] ^ layer_0[16]); 
    assign layer_1[2242] = layer_0[2297] & layer_0[2306]; 
    assign layer_1[2243] = ~(layer_0[1276] | layer_0[1199]); 
    assign layer_1[2244] = ~(layer_0[1259] ^ layer_0[1208]); 
    assign layer_1[2245] = ~(layer_0[1855] | layer_0[1870]); 
    assign layer_1[2246] = layer_0[1184] | layer_0[1160]; 
    assign layer_1[2247] = layer_0[1895] & ~layer_0[1798]; 
    assign layer_1[2248] = layer_0[554] & ~layer_0[663]; 
    assign layer_1[2249] = ~layer_0[1286] | (layer_0[1286] & layer_0[1223]); 
    assign layer_1[2250] = layer_0[2793]; 
    assign layer_1[2251] = ~layer_0[2131] | (layer_0[2168] & layer_0[2131]); 
    assign layer_1[2252] = ~layer_0[799] | (layer_0[688] & layer_0[799]); 
    assign layer_1[2253] = layer_0[2553] ^ layer_0[2509]; 
    assign layer_1[2254] = layer_0[2726]; 
    assign layer_1[2255] = ~layer_0[1898]; 
    assign layer_1[2256] = layer_0[3176] & ~layer_0[3230]; 
    assign layer_1[2257] = layer_0[3180] ^ layer_0[3195]; 
    assign layer_1[2258] = ~layer_0[3423]; 
    assign layer_1[2259] = layer_0[3113] & ~layer_0[3081]; 
    assign layer_1[2260] = layer_0[2259] & layer_0[2370]; 
    assign layer_1[2261] = layer_0[3130] & ~layer_0[3170]; 
    assign layer_1[2262] = layer_0[3105] & ~layer_0[3222]; 
    assign layer_1[2263] = ~layer_0[1217] | (layer_0[1249] & layer_0[1217]); 
    assign layer_1[2264] = layer_0[3387] & layer_0[3433]; 
    assign layer_1[2265] = layer_0[3044]; 
    assign layer_1[2266] = ~(layer_0[1064] & layer_0[1128]); 
    assign layer_1[2267] = layer_0[560] & layer_0[453]; 
    assign layer_1[2268] = ~layer_0[1979]; 
    assign layer_1[2269] = layer_0[2432] & ~layer_0[2385]; 
    assign layer_1[2270] = ~(layer_0[3190] & layer_0[3218]); 
    assign layer_1[2271] = ~layer_0[830]; 
    assign layer_1[2272] = layer_0[1047] | layer_0[1062]; 
    assign layer_1[2273] = layer_0[3361] ^ layer_0[3401]; 
    assign layer_1[2274] = ~layer_0[833]; 
    assign layer_1[2275] = layer_0[3242] & ~layer_0[3223]; 
    assign layer_1[2276] = layer_0[2783]; 
    assign layer_1[2277] = layer_0[3431] | layer_0[3502]; 
    assign layer_1[2278] = layer_0[516] & layer_0[403]; 
    assign layer_1[2279] = layer_0[1594] & layer_0[1591]; 
    assign layer_1[2280] = layer_0[3959] & ~layer_0[3850]; 
    assign layer_1[2281] = ~(layer_0[293] & layer_0[315]); 
    assign layer_1[2282] = layer_0[634] ^ layer_0[584]; 
    assign layer_1[2283] = ~layer_0[519] | (layer_0[519] & layer_0[423]); 
    assign layer_1[2284] = layer_0[3066] & layer_0[3094]; 
    assign layer_1[2285] = ~layer_0[3110]; 
    assign layer_1[2286] = layer_0[984] | layer_0[1086]; 
    assign layer_1[2287] = ~layer_0[2833] | (layer_0[2833] & layer_0[2708]); 
    assign layer_1[2288] = ~(layer_0[1099] ^ layer_0[1133]); 
    assign layer_1[2289] = layer_0[969] | layer_0[922]; 
    assign layer_1[2290] = ~layer_0[2761] | (layer_0[2863] & layer_0[2761]); 
    assign layer_1[2291] = ~layer_0[3475] | (layer_0[3469] & layer_0[3475]); 
    assign layer_1[2292] = layer_0[2075]; 
    assign layer_1[2293] = layer_0[1147] & layer_0[1269]; 
    assign layer_1[2294] = ~layer_0[1993] | (layer_0[1957] & layer_0[1993]); 
    assign layer_1[2295] = layer_0[3327]; 
    assign layer_1[2296] = layer_0[113] ^ layer_0[109]; 
    assign layer_1[2297] = ~(layer_0[1054] | layer_0[1019]); 
    assign layer_1[2298] = layer_0[2067] ^ layer_0[1958]; 
    assign layer_1[2299] = layer_0[1604] ^ layer_0[1580]; 
    assign layer_1[2300] = layer_0[1563] & ~layer_0[1528]; 
    assign layer_1[2301] = layer_0[3601]; 
    assign layer_1[2302] = layer_0[1366] & ~layer_0[1388]; 
    assign layer_1[2303] = layer_0[2448] ^ layer_0[2329]; 
    assign layer_1[2304] = ~layer_0[464]; 
    assign layer_1[2305] = ~(layer_0[2100] ^ layer_0[2041]); 
    assign layer_1[2306] = layer_0[1453]; 
    assign layer_1[2307] = ~(layer_0[503] ^ layer_0[552]); 
    assign layer_1[2308] = ~layer_0[1731]; 
    assign layer_1[2309] = ~layer_0[2751]; 
    assign layer_1[2310] = ~(layer_0[1959] & layer_0[2049]); 
    assign layer_1[2311] = layer_0[278]; 
    assign layer_1[2312] = layer_0[1623]; 
    assign layer_1[2313] = ~layer_0[477] | (layer_0[477] & layer_0[575]); 
    assign layer_1[2314] = ~(layer_0[1182] ^ layer_0[1197]); 
    assign layer_1[2315] = ~(layer_0[3657] ^ layer_0[3568]); 
    assign layer_1[2316] = ~layer_0[2756] | (layer_0[2756] & layer_0[2783]); 
    assign layer_1[2317] = layer_0[3907] | layer_0[3989]; 
    assign layer_1[2318] = layer_0[2038]; 
    assign layer_1[2319] = layer_0[1573] & ~layer_0[1696]; 
    assign layer_1[2320] = layer_0[2483] | layer_0[2424]; 
    assign layer_1[2321] = ~layer_0[1092]; 
    assign layer_1[2322] = layer_0[1315] & ~layer_0[1232]; 
    assign layer_1[2323] = layer_0[3507] ^ layer_0[3626]; 
    assign layer_1[2324] = ~(layer_0[444] ^ layer_0[319]); 
    assign layer_1[2325] = layer_0[585] ^ layer_0[695]; 
    assign layer_1[2326] = ~layer_0[2896] | (layer_0[2896] & layer_0[2793]); 
    assign layer_1[2327] = layer_0[2203] & layer_0[2205]; 
    assign layer_1[2328] = layer_0[2916] ^ layer_0[2865]; 
    assign layer_1[2329] = layer_0[2072] ^ layer_0[2061]; 
    assign layer_1[2330] = ~layer_0[3477] | (layer_0[3540] & layer_0[3477]); 
    assign layer_1[2331] = layer_0[517] | layer_0[427]; 
    assign layer_1[2332] = ~layer_0[1087]; 
    assign layer_1[2333] = ~(layer_0[1835] & layer_0[1740]); 
    assign layer_1[2334] = layer_0[132] & layer_0[58]; 
    assign layer_1[2335] = layer_0[3541]; 
    assign layer_1[2336] = layer_0[383] & ~layer_0[384]; 
    assign layer_1[2337] = layer_0[205] & layer_0[115]; 
    assign layer_1[2338] = ~layer_0[3363]; 
    assign layer_1[2339] = ~layer_0[1140]; 
    assign layer_1[2340] = layer_0[712] & ~layer_0[806]; 
    assign layer_1[2341] = layer_0[501] & ~layer_0[549]; 
    assign layer_1[2342] = ~layer_0[2088] | (layer_0[2027] & layer_0[2088]); 
    assign layer_1[2343] = layer_0[2570] & layer_0[2575]; 
    assign layer_1[2344] = ~(layer_0[2379] | layer_0[2361]); 
    assign layer_1[2345] = ~(layer_0[3102] | layer_0[3115]); 
    assign layer_1[2346] = layer_0[1068] ^ layer_0[951]; 
    assign layer_1[2347] = layer_0[1946] & ~layer_0[1971]; 
    assign layer_1[2348] = layer_0[628]; 
    assign layer_1[2349] = layer_0[3039] & ~layer_0[3153]; 
    assign layer_1[2350] = layer_0[2188] ^ layer_0[2121]; 
    assign layer_1[2351] = layer_0[184] & ~layer_0[145]; 
    assign layer_1[2352] = layer_0[113]; 
    assign layer_1[2353] = ~layer_0[1821] | (layer_0[1760] & layer_0[1821]); 
    assign layer_1[2354] = ~layer_0[3067]; 
    assign layer_1[2355] = layer_0[2385]; 
    assign layer_1[2356] = ~(layer_0[759] | layer_0[727]); 
    assign layer_1[2357] = layer_0[1185]; 
    assign layer_1[2358] = layer_0[1155] | layer_0[1282]; 
    assign layer_1[2359] = ~(layer_0[3674] & layer_0[3612]); 
    assign layer_1[2360] = ~(layer_0[622] & layer_0[520]); 
    assign layer_1[2361] = layer_0[2809] | layer_0[2722]; 
    assign layer_1[2362] = ~(layer_0[1420] ^ layer_0[1411]); 
    assign layer_1[2363] = ~(layer_0[237] & layer_0[281]); 
    assign layer_1[2364] = layer_0[3048] ^ layer_0[2949]; 
    assign layer_1[2365] = ~layer_0[1555]; 
    assign layer_1[2366] = ~layer_0[1410]; 
    assign layer_1[2367] = ~(layer_0[1279] ^ layer_0[1351]); 
    assign layer_1[2368] = layer_0[353] & ~layer_0[412]; 
    assign layer_1[2369] = layer_0[3974] & layer_0[3932]; 
    assign layer_1[2370] = layer_0[1376] | layer_0[1326]; 
    assign layer_1[2371] = ~(layer_0[926] ^ layer_0[918]); 
    assign layer_1[2372] = layer_0[1723]; 
    assign layer_1[2373] = layer_0[143]; 
    assign layer_1[2374] = layer_0[527] | layer_0[520]; 
    assign layer_1[2375] = layer_0[3658] ^ layer_0[3573]; 
    assign layer_1[2376] = layer_0[328] ^ layer_0[363]; 
    assign layer_1[2377] = layer_0[2319] & layer_0[2212]; 
    assign layer_1[2378] = layer_0[813] & layer_0[728]; 
    assign layer_1[2379] = ~layer_0[636]; 
    assign layer_1[2380] = layer_0[3994] & ~layer_0[3951]; 
    assign layer_1[2381] = ~layer_0[714] | (layer_0[714] & layer_0[826]); 
    assign layer_1[2382] = ~(layer_0[3632] & layer_0[3542]); 
    assign layer_1[2383] = layer_0[22] & ~layer_0[9]; 
    assign layer_1[2384] = layer_0[3448]; 
    assign layer_1[2385] = layer_0[625] & layer_0[544]; 
    assign layer_1[2386] = ~layer_0[210]; 
    assign layer_1[2387] = layer_0[2165] ^ layer_0[2285]; 
    assign layer_1[2388] = ~layer_0[2170]; 
    assign layer_1[2389] = layer_0[689] | layer_0[726]; 
    assign layer_1[2390] = ~layer_0[3737] | (layer_0[3705] & layer_0[3737]); 
    assign layer_1[2391] = ~layer_0[607] | (layer_0[504] & layer_0[607]); 
    assign layer_1[2392] = ~(layer_0[3226] | layer_0[3267]); 
    assign layer_1[2393] = ~layer_0[294] | (layer_0[294] & layer_0[311]); 
    assign layer_1[2394] = layer_0[1226] & layer_0[1230]; 
    assign layer_1[2395] = ~(layer_0[1335] & layer_0[1450]); 
    assign layer_1[2396] = ~layer_0[1100]; 
    assign layer_1[2397] = ~layer_0[2914] | (layer_0[3039] & layer_0[2914]); 
    assign layer_1[2398] = layer_0[1483] & ~layer_0[1572]; 
    assign layer_1[2399] = layer_0[1950] & ~layer_0[1994]; 
    assign layer_1[2400] = layer_0[3468]; 
    assign layer_1[2401] = ~(layer_0[3816] | layer_0[3749]); 
    assign layer_1[2402] = ~layer_0[3111] | (layer_0[3111] & layer_0[3094]); 
    assign layer_1[2403] = layer_0[2243] & layer_0[2357]; 
    assign layer_1[2404] = ~(layer_0[3145] | layer_0[3154]); 
    assign layer_1[2405] = ~layer_0[3044]; 
    assign layer_1[2406] = layer_0[2649] & layer_0[2575]; 
    assign layer_1[2407] = ~layer_0[3298] | (layer_0[3298] & layer_0[3411]); 
    assign layer_1[2408] = layer_0[1852] | layer_0[1750]; 
    assign layer_1[2409] = ~(layer_0[2712] | layer_0[2789]); 
    assign layer_1[2410] = ~layer_0[2928]; 
    assign layer_1[2411] = layer_0[3339]; 
    assign layer_1[2412] = layer_0[2489] ^ layer_0[2597]; 
    assign layer_1[2413] = layer_0[546] ^ layer_0[522]; 
    assign layer_1[2414] = layer_0[3605] ^ layer_0[3637]; 
    assign layer_1[2415] = layer_0[1937]; 
    assign layer_1[2416] = layer_0[3959] & ~layer_0[3974]; 
    assign layer_1[2417] = ~(layer_0[3144] ^ layer_0[3096]); 
    assign layer_1[2418] = layer_0[3568] & ~layer_0[3581]; 
    assign layer_1[2419] = ~layer_0[3447] | (layer_0[3447] & layer_0[3519]); 
    assign layer_1[2420] = ~(layer_0[2497] ^ layer_0[2621]); 
    assign layer_1[2421] = ~(layer_0[2575] ^ layer_0[2687]); 
    assign layer_1[2422] = ~(layer_0[3426] & layer_0[3371]); 
    assign layer_1[2423] = layer_0[3259]; 
    assign layer_1[2424] = ~layer_0[3971]; 
    assign layer_1[2425] = layer_0[3681]; 
    assign layer_1[2426] = layer_0[1258] ^ layer_0[1372]; 
    assign layer_1[2427] = ~layer_0[697] | (layer_0[814] & layer_0[697]); 
    assign layer_1[2428] = layer_0[1232] ^ layer_0[1334]; 
    assign layer_1[2429] = ~(layer_0[523] | layer_0[491]); 
    assign layer_1[2430] = ~(layer_0[971] ^ layer_0[1015]); 
    assign layer_1[2431] = ~layer_0[305]; 
    assign layer_1[2432] = ~layer_0[3353] | (layer_0[3353] & layer_0[3283]); 
    assign layer_1[2433] = ~(layer_0[653] ^ layer_0[596]); 
    assign layer_1[2434] = layer_0[2695]; 
    assign layer_1[2435] = ~(layer_0[3350] | layer_0[3329]); 
    assign layer_1[2436] = layer_0[952]; 
    assign layer_1[2437] = ~layer_0[3706] | (layer_0[3706] & layer_0[3791]); 
    assign layer_1[2438] = layer_0[2978] & ~layer_0[2963]; 
    assign layer_1[2439] = ~layer_0[1606] | (layer_0[1506] & layer_0[1606]); 
    assign layer_1[2440] = layer_0[2243] | layer_0[2234]; 
    assign layer_1[2441] = ~layer_0[8] | (layer_0[51] & layer_0[8]); 
    assign layer_1[2442] = layer_0[3199] & ~layer_0[3231]; 
    assign layer_1[2443] = ~(layer_0[2223] | layer_0[2266]); 
    assign layer_1[2444] = ~(layer_0[1405] & layer_0[1434]); 
    assign layer_1[2445] = layer_0[746] & layer_0[642]; 
    assign layer_1[2446] = layer_0[3630]; 
    assign layer_1[2447] = layer_0[2741] & layer_0[2860]; 
    assign layer_1[2448] = ~layer_0[474]; 
    assign layer_1[2449] = layer_0[541] ^ layer_0[520]; 
    assign layer_1[2450] = ~(layer_0[872] | layer_0[956]); 
    assign layer_1[2451] = layer_0[1697]; 
    assign layer_1[2452] = ~(layer_0[93] & layer_0[102]); 
    assign layer_1[2453] = layer_0[1171]; 
    assign layer_1[2454] = layer_0[451] & ~layer_0[367]; 
    assign layer_1[2455] = layer_0[2155] & ~layer_0[2207]; 
    assign layer_1[2456] = layer_0[745]; 
    assign layer_1[2457] = layer_0[2675] & ~layer_0[2673]; 
    assign layer_1[2458] = layer_0[215] ^ layer_0[95]; 
    assign layer_1[2459] = layer_0[181] ^ layer_0[204]; 
    assign layer_1[2460] = ~(layer_0[661] ^ layer_0[738]); 
    assign layer_1[2461] = ~layer_0[1679]; 
    assign layer_1[2462] = layer_0[2203] & ~layer_0[2217]; 
    assign layer_1[2463] = ~(layer_0[539] | layer_0[432]); 
    assign layer_1[2464] = layer_0[3293] & ~layer_0[3308]; 
    assign layer_1[2465] = layer_0[2234] ^ layer_0[2271]; 
    assign layer_1[2466] = ~(layer_0[2262] & layer_0[2216]); 
    assign layer_1[2467] = layer_0[3261] & ~layer_0[3380]; 
    assign layer_1[2468] = layer_0[3000]; 
    assign layer_1[2469] = layer_0[2906] & layer_0[3012]; 
    assign layer_1[2470] = layer_0[1839] & ~layer_0[1871]; 
    assign layer_1[2471] = ~layer_0[577]; 
    assign layer_1[2472] = ~layer_0[745] | (layer_0[745] & layer_0[688]); 
    assign layer_1[2473] = ~layer_0[3250]; 
    assign layer_1[2474] = ~layer_0[612] | (layer_0[612] & layer_0[636]); 
    assign layer_1[2475] = ~layer_0[875] | (layer_0[765] & layer_0[875]); 
    assign layer_1[2476] = layer_0[806] & ~layer_0[832]; 
    assign layer_1[2477] = ~layer_0[1073]; 
    assign layer_1[2478] = ~layer_0[1634]; 
    assign layer_1[2479] = layer_0[3714]; 
    assign layer_1[2480] = layer_0[310] ^ layer_0[285]; 
    assign layer_1[2481] = ~(layer_0[2957] | layer_0[2873]); 
    assign layer_1[2482] = ~(layer_0[3079] ^ layer_0[3096]); 
    assign layer_1[2483] = ~(layer_0[3665] ^ layer_0[3782]); 
    assign layer_1[2484] = ~(layer_0[2991] ^ layer_0[2896]); 
    assign layer_1[2485] = layer_0[3442] | layer_0[3451]; 
    assign layer_1[2486] = ~layer_0[1277]; 
    assign layer_1[2487] = ~layer_0[236]; 
    assign layer_1[2488] = layer_0[3200] ^ layer_0[3117]; 
    assign layer_1[2489] = layer_0[3933] & ~layer_0[3898]; 
    assign layer_1[2490] = ~(layer_0[2427] & layer_0[2513]); 
    assign layer_1[2491] = ~layer_0[3118] | (layer_0[3174] & layer_0[3118]); 
    assign layer_1[2492] = ~layer_0[3987]; 
    assign layer_1[2493] = ~layer_0[3757] | (layer_0[3802] & layer_0[3757]); 
    assign layer_1[2494] = ~layer_0[3914] | (layer_0[3914] & layer_0[3954]); 
    assign layer_1[2495] = layer_0[3526] ^ layer_0[3558]; 
    assign layer_1[2496] = layer_0[146]; 
    assign layer_1[2497] = ~layer_0[1015]; 
    assign layer_1[2498] = ~(layer_0[2914] | layer_0[3034]); 
    assign layer_1[2499] = ~layer_0[2743]; 
    assign layer_1[2500] = ~layer_0[905]; 
    assign layer_1[2501] = ~(layer_0[2984] & layer_0[2869]); 
    assign layer_1[2502] = layer_0[905] | layer_0[858]; 
    assign layer_1[2503] = layer_0[1348]; 
    assign layer_1[2504] = layer_0[89] & ~layer_0[71]; 
    assign layer_1[2505] = ~layer_0[3146] | (layer_0[3102] & layer_0[3146]); 
    assign layer_1[2506] = layer_0[555] ^ layer_0[622]; 
    assign layer_1[2507] = layer_0[964] | layer_0[1075]; 
    assign layer_1[2508] = layer_0[2462] ^ layer_0[2534]; 
    assign layer_1[2509] = ~layer_0[685]; 
    assign layer_1[2510] = ~layer_0[324]; 
    assign layer_1[2511] = layer_0[1417] ^ layer_0[1347]; 
    assign layer_1[2512] = ~(layer_0[1639] ^ layer_0[1638]); 
    assign layer_1[2513] = ~layer_0[408] | (layer_0[408] & layer_0[324]); 
    assign layer_1[2514] = layer_0[234]; 
    assign layer_1[2515] = ~layer_0[526]; 
    assign layer_1[2516] = layer_0[3137] & ~layer_0[3210]; 
    assign layer_1[2517] = ~layer_0[3913] | (layer_0[3913] & layer_0[3901]); 
    assign layer_1[2518] = ~(layer_0[2763] | layer_0[2664]); 
    assign layer_1[2519] = ~(layer_0[2405] | layer_0[2398]); 
    assign layer_1[2520] = ~(layer_0[621] & layer_0[579]); 
    assign layer_1[2521] = layer_0[501]; 
    assign layer_1[2522] = ~layer_0[2523] | (layer_0[2523] & layer_0[2539]); 
    assign layer_1[2523] = layer_0[1025] & ~layer_0[1149]; 
    assign layer_1[2524] = ~layer_0[3955] | (layer_0[3885] & layer_0[3955]); 
    assign layer_1[2525] = ~(layer_0[3823] ^ layer_0[3697]); 
    assign layer_1[2526] = layer_0[1634]; 
    assign layer_1[2527] = layer_0[975] ^ layer_0[852]; 
    assign layer_1[2528] = ~layer_0[2592] | (layer_0[2592] & layer_0[2646]); 
    assign layer_1[2529] = layer_0[1452]; 
    assign layer_1[2530] = layer_0[3107] | layer_0[3233]; 
    assign layer_1[2531] = ~(layer_0[3765] ^ layer_0[3722]); 
    assign layer_1[2532] = layer_0[2980]; 
    assign layer_1[2533] = layer_0[2598]; 
    assign layer_1[2534] = layer_0[2111] & ~layer_0[2216]; 
    assign layer_1[2535] = layer_0[2733] ^ layer_0[2849]; 
    assign layer_1[2536] = ~layer_0[3361]; 
    assign layer_1[2537] = ~(layer_0[545] | layer_0[422]); 
    assign layer_1[2538] = layer_0[1958] ^ layer_0[1908]; 
    assign layer_1[2539] = layer_0[311] & layer_0[186]; 
    assign layer_1[2540] = ~(layer_0[794] | layer_0[916]); 
    assign layer_1[2541] = layer_0[3384] & ~layer_0[3275]; 
    assign layer_1[2542] = ~(layer_0[2615] | layer_0[2572]); 
    assign layer_1[2543] = ~layer_0[3228] | (layer_0[3228] & layer_0[3330]); 
    assign layer_1[2544] = layer_0[2214]; 
    assign layer_1[2545] = ~(layer_0[137] ^ layer_0[95]); 
    assign layer_1[2546] = ~(layer_0[1223] ^ layer_0[1345]); 
    assign layer_1[2547] = layer_0[1838] & ~layer_0[1773]; 
    assign layer_1[2548] = ~(layer_0[1986] & layer_0[1900]); 
    assign layer_1[2549] = ~(layer_0[1581] & layer_0[1475]); 
    assign layer_1[2550] = ~layer_0[1828]; 
    assign layer_1[2551] = ~(layer_0[1423] & layer_0[1451]); 
    assign layer_1[2552] = layer_0[3836] & ~layer_0[3927]; 
    assign layer_1[2553] = layer_0[3604] & ~layer_0[3642]; 
    assign layer_1[2554] = layer_0[1835] & ~layer_0[1726]; 
    assign layer_1[2555] = layer_0[2426] & ~layer_0[2503]; 
    assign layer_1[2556] = layer_0[1004]; 
    assign layer_1[2557] = layer_0[120] & layer_0[194]; 
    assign layer_1[2558] = ~(layer_0[30] & layer_0[100]); 
    assign layer_1[2559] = layer_0[200] & ~layer_0[206]; 
    assign layer_1[2560] = ~(layer_0[1516] | layer_0[1462]); 
    assign layer_1[2561] = ~(layer_0[3853] ^ layer_0[3885]); 
    assign layer_1[2562] = ~layer_0[131] | (layer_0[131] & layer_0[58]); 
    assign layer_1[2563] = ~(layer_0[2059] | layer_0[1947]); 
    assign layer_1[2564] = ~(layer_0[2613] | layer_0[2686]); 
    assign layer_1[2565] = layer_0[1452] | layer_0[1325]; 
    assign layer_1[2566] = ~(layer_0[590] ^ layer_0[643]); 
    assign layer_1[2567] = ~layer_0[3055]; 
    assign layer_1[2568] = layer_0[899] ^ layer_0[778]; 
    assign layer_1[2569] = layer_0[3835] & ~layer_0[3807]; 
    assign layer_1[2570] = layer_0[1993]; 
    assign layer_1[2571] = ~(layer_0[489] | layer_0[552]); 
    assign layer_1[2572] = ~layer_0[1400] | (layer_0[1400] & layer_0[1300]); 
    assign layer_1[2573] = ~layer_0[1502]; 
    assign layer_1[2574] = layer_0[3129] & layer_0[3078]; 
    assign layer_1[2575] = layer_0[2350] & ~layer_0[2421]; 
    assign layer_1[2576] = layer_0[1899]; 
    assign layer_1[2577] = ~(layer_0[2495] | layer_0[2371]); 
    assign layer_1[2578] = layer_0[2523] & ~layer_0[2618]; 
    assign layer_1[2579] = ~layer_0[901] | (layer_0[855] & layer_0[901]); 
    assign layer_1[2580] = ~layer_0[2759]; 
    assign layer_1[2581] = layer_0[2376] & ~layer_0[2291]; 
    assign layer_1[2582] = ~(layer_0[1006] | layer_0[982]); 
    assign layer_1[2583] = ~(layer_0[2987] & layer_0[3105]); 
    assign layer_1[2584] = ~(layer_0[1558] & layer_0[1548]); 
    assign layer_1[2585] = ~(layer_0[1684] | layer_0[1637]); 
    assign layer_1[2586] = layer_0[2159] | layer_0[2239]; 
    assign layer_1[2587] = ~layer_0[1337] | (layer_0[1298] & layer_0[1337]); 
    assign layer_1[2588] = layer_0[2803] & layer_0[2708]; 
    assign layer_1[2589] = ~(layer_0[3477] | layer_0[3545]); 
    assign layer_1[2590] = layer_0[3050] & ~layer_0[3166]; 
    assign layer_1[2591] = ~layer_0[1427]; 
    assign layer_1[2592] = layer_0[1767] & ~layer_0[1791]; 
    assign layer_1[2593] = ~layer_0[708]; 
    assign layer_1[2594] = ~layer_0[2971]; 
    assign layer_1[2595] = ~(layer_0[2232] & layer_0[2121]); 
    assign layer_1[2596] = ~layer_0[558]; 
    assign layer_1[2597] = ~layer_0[2276] | (layer_0[2358] & layer_0[2276]); 
    assign layer_1[2598] = layer_0[669] & layer_0[573]; 
    assign layer_1[2599] = ~layer_0[887]; 
    assign layer_1[2600] = ~(layer_0[3771] ^ layer_0[3744]); 
    assign layer_1[2601] = layer_0[3475]; 
    assign layer_1[2602] = layer_0[764] & ~layer_0[790]; 
    assign layer_1[2603] = layer_0[1967] & ~layer_0[2086]; 
    assign layer_1[2604] = ~(layer_0[1294] ^ layer_0[1272]); 
    assign layer_1[2605] = ~(layer_0[1953] & layer_0[2065]); 
    assign layer_1[2606] = ~layer_0[655]; 
    assign layer_1[2607] = layer_0[661] & ~layer_0[571]; 
    assign layer_1[2608] = ~(layer_0[1354] ^ layer_0[1314]); 
    assign layer_1[2609] = layer_0[1867] & ~layer_0[1744]; 
    assign layer_1[2610] = ~layer_0[1541]; 
    assign layer_1[2611] = ~layer_0[753]; 
    assign layer_1[2612] = layer_0[741] & layer_0[780]; 
    assign layer_1[2613] = layer_0[2682] | layer_0[2808]; 
    assign layer_1[2614] = layer_0[626] & layer_0[643]; 
    assign layer_1[2615] = layer_0[3935]; 
    assign layer_1[2616] = ~layer_0[3702]; 
    assign layer_1[2617] = layer_0[1883]; 
    assign layer_1[2618] = layer_0[1550]; 
    assign layer_1[2619] = layer_0[2988]; 
    assign layer_1[2620] = ~(layer_0[2274] | layer_0[2378]); 
    assign layer_1[2621] = layer_0[2752] ^ layer_0[2856]; 
    assign layer_1[2622] = layer_0[1028] | layer_0[969]; 
    assign layer_1[2623] = layer_0[2586]; 
    assign layer_1[2624] = layer_0[3451] & layer_0[3491]; 
    assign layer_1[2625] = layer_0[938] & ~layer_0[956]; 
    assign layer_1[2626] = layer_0[1483]; 
    assign layer_1[2627] = layer_0[3622] | layer_0[3570]; 
    assign layer_1[2628] = ~(layer_0[1942] | layer_0[1957]); 
    assign layer_1[2629] = ~layer_0[2435]; 
    assign layer_1[2630] = ~layer_0[401] | (layer_0[336] & layer_0[401]); 
    assign layer_1[2631] = layer_0[3502] & ~layer_0[3484]; 
    assign layer_1[2632] = layer_0[3186]; 
    assign layer_1[2633] = ~(layer_0[3201] & layer_0[3326]); 
    assign layer_1[2634] = ~layer_0[3455]; 
    assign layer_1[2635] = layer_0[3066] ^ layer_0[3171]; 
    assign layer_1[2636] = ~(layer_0[2064] | layer_0[2159]); 
    assign layer_1[2637] = layer_0[2158]; 
    assign layer_1[2638] = ~layer_0[2082]; 
    assign layer_1[2639] = ~layer_0[608]; 
    assign layer_1[2640] = ~layer_0[3019]; 
    assign layer_1[2641] = layer_0[2798] & layer_0[2788]; 
    assign layer_1[2642] = ~layer_0[1225]; 
    assign layer_1[2643] = layer_0[386] & ~layer_0[366]; 
    assign layer_1[2644] = layer_0[883] & ~layer_0[902]; 
    assign layer_1[2645] = layer_0[1855]; 
    assign layer_1[2646] = ~(layer_0[2703] | layer_0[2821]); 
    assign layer_1[2647] = ~(layer_0[1386] ^ layer_0[1331]); 
    assign layer_1[2648] = layer_0[3256]; 
    assign layer_1[2649] = ~layer_0[485]; 
    assign layer_1[2650] = ~(layer_0[2732] ^ layer_0[2727]); 
    assign layer_1[2651] = ~layer_0[2737] | (layer_0[2737] & layer_0[2635]); 
    assign layer_1[2652] = layer_0[651] & layer_0[777]; 
    assign layer_1[2653] = ~(layer_0[2004] & layer_0[1954]); 
    assign layer_1[2654] = ~layer_0[2866]; 
    assign layer_1[2655] = layer_0[2811] & layer_0[2694]; 
    assign layer_1[2656] = ~layer_0[1950] | (layer_0[1892] & layer_0[1950]); 
    assign layer_1[2657] = ~layer_0[1664]; 
    assign layer_1[2658] = layer_0[281] ^ layer_0[397]; 
    assign layer_1[2659] = layer_0[198]; 
    assign layer_1[2660] = layer_0[2538]; 
    assign layer_1[2661] = layer_0[2252] ^ layer_0[2274]; 
    assign layer_1[2662] = layer_0[2395] & layer_0[2480]; 
    assign layer_1[2663] = layer_0[1852]; 
    assign layer_1[2664] = layer_0[3592]; 
    assign layer_1[2665] = ~layer_0[2418]; 
    assign layer_1[2666] = layer_0[3783] & ~layer_0[3738]; 
    assign layer_1[2667] = ~(layer_0[3486] ^ layer_0[3531]); 
    assign layer_1[2668] = ~layer_0[1641] | (layer_0[1641] & layer_0[1706]); 
    assign layer_1[2669] = ~layer_0[328]; 
    assign layer_1[2670] = layer_0[276] & layer_0[363]; 
    assign layer_1[2671] = ~layer_0[3882]; 
    assign layer_1[2672] = ~(layer_0[1783] ^ layer_0[1730]); 
    assign layer_1[2673] = ~layer_0[2727] | (layer_0[2734] & layer_0[2727]); 
    assign layer_1[2674] = ~layer_0[2387]; 
    assign layer_1[2675] = ~layer_0[332]; 
    assign layer_1[2676] = ~layer_0[412]; 
    assign layer_1[2677] = layer_0[123] & ~layer_0[222]; 
    assign layer_1[2678] = ~layer_0[393]; 
    assign layer_1[2679] = layer_0[3263]; 
    assign layer_1[2680] = layer_0[3547]; 
    assign layer_1[2681] = ~layer_0[1827] | (layer_0[1719] & layer_0[1827]); 
    assign layer_1[2682] = ~(layer_0[445] ^ layer_0[390]); 
    assign layer_1[2683] = layer_0[672] & ~layer_0[703]; 
    assign layer_1[2684] = ~(layer_0[792] ^ layer_0[722]); 
    assign layer_1[2685] = ~layer_0[3455] | (layer_0[3535] & layer_0[3455]); 
    assign layer_1[2686] = layer_0[2858]; 
    assign layer_1[2687] = layer_0[219]; 
    assign layer_1[2688] = layer_0[373] & ~layer_0[457]; 
    assign layer_1[2689] = ~layer_0[1467] | (layer_0[1465] & layer_0[1467]); 
    assign layer_1[2690] = layer_0[1866] ^ layer_0[1773]; 
    assign layer_1[2691] = layer_0[2049]; 
    assign layer_1[2692] = ~(layer_0[616] | layer_0[546]); 
    assign layer_1[2693] = layer_0[3705]; 
    assign layer_1[2694] = ~layer_0[983] | (layer_0[1023] & layer_0[983]); 
    assign layer_1[2695] = ~layer_0[3101]; 
    assign layer_1[2696] = layer_0[2670] & ~layer_0[2755]; 
    assign layer_1[2697] = layer_0[3221] & layer_0[3126]; 
    assign layer_1[2698] = ~layer_0[547]; 
    assign layer_1[2699] = layer_0[942] ^ layer_0[1028]; 
    assign layer_1[2700] = layer_0[2887]; 
    assign layer_1[2701] = layer_0[1795]; 
    assign layer_1[2702] = ~(layer_0[49] & layer_0[95]); 
    assign layer_1[2703] = layer_0[2462] & layer_0[2350]; 
    assign layer_1[2704] = layer_0[955]; 
    assign layer_1[2705] = ~layer_0[2697]; 
    assign layer_1[2706] = ~(layer_0[355] | layer_0[408]); 
    assign layer_1[2707] = ~layer_0[374] | (layer_0[374] & layer_0[291]); 
    assign layer_1[2708] = layer_0[146]; 
    assign layer_1[2709] = layer_0[1223]; 
    assign layer_1[2710] = ~layer_0[1666]; 
    assign layer_1[2711] = layer_0[1866] & ~layer_0[1803]; 
    assign layer_1[2712] = ~layer_0[798] | (layer_0[721] & layer_0[798]); 
    assign layer_1[2713] = ~layer_0[3024] | (layer_0[3024] & layer_0[2965]); 
    assign layer_1[2714] = ~(layer_0[2477] ^ layer_0[2524]); 
    assign layer_1[2715] = ~(layer_0[3729] | layer_0[3685]); 
    assign layer_1[2716] = ~layer_0[1900]; 
    assign layer_1[2717] = ~layer_0[1794]; 
    assign layer_1[2718] = layer_0[694] & ~layer_0[723]; 
    assign layer_1[2719] = ~layer_0[2697]; 
    assign layer_1[2720] = layer_0[1744]; 
    assign layer_1[2721] = layer_0[2122] & ~layer_0[2027]; 
    assign layer_1[2722] = layer_0[1771] | layer_0[1813]; 
    assign layer_1[2723] = ~(layer_0[1146] ^ layer_0[1160]); 
    assign layer_1[2724] = layer_0[1402] | layer_0[1421]; 
    assign layer_1[2725] = ~layer_0[2044] | (layer_0[2022] & layer_0[2044]); 
    assign layer_1[2726] = layer_0[395] & layer_0[294]; 
    assign layer_1[2727] = layer_0[170]; 
    assign layer_1[2728] = ~(layer_0[381] | layer_0[439]); 
    assign layer_1[2729] = ~layer_0[1735] | (layer_0[1735] & layer_0[1656]); 
    assign layer_1[2730] = ~layer_0[690]; 
    assign layer_1[2731] = layer_0[2614]; 
    assign layer_1[2732] = layer_0[3068]; 
    assign layer_1[2733] = ~(layer_0[2220] ^ layer_0[2204]); 
    assign layer_1[2734] = ~(layer_0[3189] & layer_0[3185]); 
    assign layer_1[2735] = ~layer_0[3086] | (layer_0[3181] & layer_0[3086]); 
    assign layer_1[2736] = ~(layer_0[2761] ^ layer_0[2873]); 
    assign layer_1[2737] = layer_0[1265] & ~layer_0[1292]; 
    assign layer_1[2738] = ~(layer_0[2133] | layer_0[2205]); 
    assign layer_1[2739] = ~layer_0[1503]; 
    assign layer_1[2740] = layer_0[2724]; 
    assign layer_1[2741] = ~(layer_0[1030] | layer_0[957]); 
    assign layer_1[2742] = layer_0[572] & ~layer_0[604]; 
    assign layer_1[2743] = layer_0[227]; 
    assign layer_1[2744] = ~layer_0[1521] | (layer_0[1521] & layer_0[1541]); 
    assign layer_1[2745] = layer_0[3660] & ~layer_0[3705]; 
    assign layer_1[2746] = layer_0[325] ^ layer_0[345]; 
    assign layer_1[2747] = layer_0[3548]; 
    assign layer_1[2748] = layer_0[2430] ^ layer_0[2306]; 
    assign layer_1[2749] = layer_0[1518]; 
    assign layer_1[2750] = ~layer_0[2994]; 
    assign layer_1[2751] = ~layer_0[2376]; 
    assign layer_1[2752] = ~(layer_0[3790] & layer_0[3785]); 
    assign layer_1[2753] = layer_0[2671] & ~layer_0[2678]; 
    assign layer_1[2754] = layer_0[1960]; 
    assign layer_1[2755] = ~(layer_0[2600] | layer_0[2700]); 
    assign layer_1[2756] = ~layer_0[2258] | (layer_0[2258] & layer_0[2247]); 
    assign layer_1[2757] = layer_0[2342] & ~layer_0[2402]; 
    assign layer_1[2758] = layer_0[3812] | layer_0[3831]; 
    assign layer_1[2759] = ~(layer_0[2626] & layer_0[2727]); 
    assign layer_1[2760] = layer_0[3544] & layer_0[3562]; 
    assign layer_1[2761] = layer_0[2362] & layer_0[2258]; 
    assign layer_1[2762] = layer_0[2160] & ~layer_0[2256]; 
    assign layer_1[2763] = layer_0[1683]; 
    assign layer_1[2764] = ~(layer_0[3075] | layer_0[3172]); 
    assign layer_1[2765] = layer_0[845] | layer_0[879]; 
    assign layer_1[2766] = ~layer_0[1501]; 
    assign layer_1[2767] = ~(layer_0[1773] | layer_0[1744]); 
    assign layer_1[2768] = ~(layer_0[83] & layer_0[165]); 
    assign layer_1[2769] = layer_0[1014]; 
    assign layer_1[2770] = layer_0[3900] & ~layer_0[3865]; 
    assign layer_1[2771] = layer_0[2121] | layer_0[2086]; 
    assign layer_1[2772] = ~layer_0[2125] | (layer_0[2125] & layer_0[2199]); 
    assign layer_1[2773] = layer_0[1373] & layer_0[1434]; 
    assign layer_1[2774] = ~layer_0[574]; 
    assign layer_1[2775] = layer_0[1931] | layer_0[2002]; 
    assign layer_1[2776] = ~layer_0[1857]; 
    assign layer_1[2777] = ~layer_0[817]; 
    assign layer_1[2778] = layer_0[2438] | layer_0[2378]; 
    assign layer_1[2779] = ~layer_0[555]; 
    assign layer_1[2780] = layer_0[224] & ~layer_0[206]; 
    assign layer_1[2781] = layer_0[1185]; 
    assign layer_1[2782] = layer_0[1620] & ~layer_0[1508]; 
    assign layer_1[2783] = ~layer_0[182]; 
    assign layer_1[2784] = ~layer_0[1782] | (layer_0[1782] & layer_0[1708]); 
    assign layer_1[2785] = ~(layer_0[3100] | layer_0[3204]); 
    assign layer_1[2786] = layer_0[1236] & ~layer_0[1244]; 
    assign layer_1[2787] = layer_0[2532]; 
    assign layer_1[2788] = ~layer_0[3036]; 
    assign layer_1[2789] = layer_0[3134] ^ layer_0[3093]; 
    assign layer_1[2790] = layer_0[1235] & layer_0[1337]; 
    assign layer_1[2791] = ~(layer_0[1155] | layer_0[1072]); 
    assign layer_1[2792] = ~layer_0[165]; 
    assign layer_1[2793] = layer_0[2770] ^ layer_0[2756]; 
    assign layer_1[2794] = ~(layer_0[896] | layer_0[806]); 
    assign layer_1[2795] = ~layer_0[1260] | (layer_0[1331] & layer_0[1260]); 
    assign layer_1[2796] = ~(layer_0[1320] & layer_0[1433]); 
    assign layer_1[2797] = ~(layer_0[1914] & layer_0[1915]); 
    assign layer_1[2798] = layer_0[223]; 
    assign layer_1[2799] = ~layer_0[325]; 
    assign layer_1[2800] = layer_0[3363]; 
    assign layer_1[2801] = layer_0[3438] ^ layer_0[3442]; 
    assign layer_1[2802] = layer_0[39] & ~layer_0[38]; 
    assign layer_1[2803] = layer_0[1218] ^ layer_0[1196]; 
    assign layer_1[2804] = ~layer_0[1208] | (layer_0[1208] & layer_0[1317]); 
    assign layer_1[2805] = ~(layer_0[34] ^ layer_0[84]); 
    assign layer_1[2806] = ~(layer_0[3416] & layer_0[3297]); 
    assign layer_1[2807] = layer_0[2840] & layer_0[2738]; 
    assign layer_1[2808] = layer_0[2679] | layer_0[2647]; 
    assign layer_1[2809] = layer_0[3513] & ~layer_0[3442]; 
    assign layer_1[2810] = ~(layer_0[1101] | layer_0[1045]); 
    assign layer_1[2811] = layer_0[3836] & ~layer_0[3795]; 
    assign layer_1[2812] = layer_0[1541]; 
    assign layer_1[2813] = layer_0[3981] ^ layer_0[3886]; 
    assign layer_1[2814] = layer_0[3836] & ~layer_0[3866]; 
    assign layer_1[2815] = ~(layer_0[1789] ^ layer_0[1909]); 
    assign layer_1[2816] = layer_0[2827] & layer_0[2907]; 
    assign layer_1[2817] = ~layer_0[3602] | (layer_0[3690] & layer_0[3602]); 
    assign layer_1[2818] = layer_0[2763] & ~layer_0[2791]; 
    assign layer_1[2819] = layer_0[674] & ~layer_0[711]; 
    assign layer_1[2820] = layer_0[2768] ^ layer_0[2671]; 
    assign layer_1[2821] = layer_0[2316]; 
    assign layer_1[2822] = ~layer_0[3678]; 
    assign layer_1[2823] = layer_0[3390] & ~layer_0[3483]; 
    assign layer_1[2824] = ~layer_0[209] | (layer_0[209] & layer_0[208]); 
    assign layer_1[2825] = layer_0[3954] | layer_0[3960]; 
    assign layer_1[2826] = layer_0[3173]; 
    assign layer_1[2827] = ~layer_0[3211] | (layer_0[3211] & layer_0[3240]); 
    assign layer_1[2828] = ~layer_0[50] | (layer_0[50] & layer_0[112]); 
    assign layer_1[2829] = layer_0[1534]; 
    assign layer_1[2830] = layer_0[2914] & ~layer_0[2863]; 
    assign layer_1[2831] = ~(layer_0[325] & layer_0[272]); 
    assign layer_1[2832] = layer_0[269] | layer_0[351]; 
    assign layer_1[2833] = ~layer_0[3462]; 
    assign layer_1[2834] = layer_0[3755] ^ layer_0[3644]; 
    assign layer_1[2835] = layer_0[3930] ^ layer_0[3967]; 
    assign layer_1[2836] = layer_0[2459]; 
    assign layer_1[2837] = ~layer_0[3668]; 
    assign layer_1[2838] = layer_0[3403] | layer_0[3420]; 
    assign layer_1[2839] = layer_0[1894]; 
    assign layer_1[2840] = layer_0[2751] & ~layer_0[2636]; 
    assign layer_1[2841] = layer_0[1844] & layer_0[1909]; 
    assign layer_1[2842] = ~layer_0[3924]; 
    assign layer_1[2843] = layer_0[2180] ^ layer_0[2273]; 
    assign layer_1[2844] = ~layer_0[1699]; 
    assign layer_1[2845] = ~layer_0[1330]; 
    assign layer_1[2846] = layer_0[2681] & ~layer_0[2622]; 
    assign layer_1[2847] = layer_0[1671] ^ layer_0[1777]; 
    assign layer_1[2848] = layer_0[565] ^ layer_0[582]; 
    assign layer_1[2849] = ~layer_0[3645]; 
    assign layer_1[2850] = ~layer_0[3919]; 
    assign layer_1[2851] = layer_0[3545]; 
    assign layer_1[2852] = ~(layer_0[2535] & layer_0[2424]); 
    assign layer_1[2853] = layer_0[267] | layer_0[191]; 
    assign layer_1[2854] = layer_0[834]; 
    assign layer_1[2855] = layer_0[2608]; 
    assign layer_1[2856] = layer_0[2536]; 
    assign layer_1[2857] = layer_0[3667] & layer_0[3646]; 
    assign layer_1[2858] = ~(layer_0[2898] | layer_0[2889]); 
    assign layer_1[2859] = ~layer_0[1604]; 
    assign layer_1[2860] = layer_0[671]; 
    assign layer_1[2861] = layer_0[1981] ^ layer_0[2066]; 
    assign layer_1[2862] = layer_0[1410]; 
    assign layer_1[2863] = layer_0[1634]; 
    assign layer_1[2864] = layer_0[954]; 
    assign layer_1[2865] = layer_0[349] | layer_0[355]; 
    assign layer_1[2866] = layer_0[1827] ^ layer_0[1802]; 
    assign layer_1[2867] = ~(layer_0[2975] ^ layer_0[3000]); 
    assign layer_1[2868] = ~(layer_0[2779] ^ layer_0[2657]); 
    assign layer_1[2869] = layer_0[2588]; 
    assign layer_1[2870] = layer_0[2630] & layer_0[2620]; 
    assign layer_1[2871] = ~(layer_0[3781] ^ layer_0[3875]); 
    assign layer_1[2872] = layer_0[972] & ~layer_0[1015]; 
    assign layer_1[2873] = layer_0[3755] | layer_0[3822]; 
    assign layer_1[2874] = layer_0[1901]; 
    assign layer_1[2875] = ~layer_0[731] | (layer_0[804] & layer_0[731]); 
    assign layer_1[2876] = layer_0[3750] & layer_0[3772]; 
    assign layer_1[2877] = ~layer_0[403] | (layer_0[418] & layer_0[403]); 
    assign layer_1[2878] = ~layer_0[2362]; 
    assign layer_1[2879] = ~(layer_0[1329] ^ layer_0[1334]); 
    assign layer_1[2880] = ~layer_0[1514]; 
    assign layer_1[2881] = ~layer_0[1039]; 
    assign layer_1[2882] = ~layer_0[2866]; 
    assign layer_1[2883] = layer_0[3211] ^ layer_0[3141]; 
    assign layer_1[2884] = layer_0[2034] ^ layer_0[1956]; 
    assign layer_1[2885] = ~(layer_0[95] | layer_0[91]); 
    assign layer_1[2886] = layer_0[3364]; 
    assign layer_1[2887] = ~layer_0[1546]; 
    assign layer_1[2888] = layer_0[1134] | layer_0[1189]; 
    assign layer_1[2889] = ~(layer_0[2027] & layer_0[2123]); 
    assign layer_1[2890] = layer_0[1822] ^ layer_0[1779]; 
    assign layer_1[2891] = layer_0[1694] & ~layer_0[1584]; 
    assign layer_1[2892] = layer_0[3515]; 
    assign layer_1[2893] = ~layer_0[501] | (layer_0[434] & layer_0[501]); 
    assign layer_1[2894] = ~(layer_0[555] & layer_0[574]); 
    assign layer_1[2895] = ~layer_0[42]; 
    assign layer_1[2896] = layer_0[2826] & layer_0[2810]; 
    assign layer_1[2897] = layer_0[630] ^ layer_0[608]; 
    assign layer_1[2898] = layer_0[3312] & layer_0[3304]; 
    assign layer_1[2899] = layer_0[3343] & layer_0[3379]; 
    assign layer_1[2900] = layer_0[2568]; 
    assign layer_1[2901] = ~(layer_0[2486] & layer_0[2505]); 
    assign layer_1[2902] = layer_0[1149] | layer_0[1194]; 
    assign layer_1[2903] = layer_0[2798] & ~layer_0[2739]; 
    assign layer_1[2904] = ~layer_0[933]; 
    assign layer_1[2905] = layer_0[3272] ^ layer_0[3294]; 
    assign layer_1[2906] = layer_0[2327] & layer_0[2356]; 
    assign layer_1[2907] = ~layer_0[1397]; 
    assign layer_1[2908] = ~layer_0[1786] | (layer_0[1786] & layer_0[1904]); 
    assign layer_1[2909] = layer_0[3007] & ~layer_0[3033]; 
    assign layer_1[2910] = layer_0[3315] | layer_0[3308]; 
    assign layer_1[2911] = layer_0[576]; 
    assign layer_1[2912] = layer_0[3955] & layer_0[3993]; 
    assign layer_1[2913] = layer_0[485]; 
    assign layer_1[2914] = ~layer_0[422]; 
    assign layer_1[2915] = ~(layer_0[1827] | layer_0[1833]); 
    assign layer_1[2916] = ~layer_0[3242]; 
    assign layer_1[2917] = ~layer_0[71]; 
    assign layer_1[2918] = ~(layer_0[1170] ^ layer_0[1050]); 
    assign layer_1[2919] = ~layer_0[2647] | (layer_0[2647] & layer_0[2753]); 
    assign layer_1[2920] = ~layer_0[1128]; 
    assign layer_1[2921] = ~layer_0[3270]; 
    assign layer_1[2922] = layer_0[2799] & ~layer_0[2926]; 
    assign layer_1[2923] = ~(layer_0[1571] | layer_0[1559]); 
    assign layer_1[2924] = layer_0[1371] | layer_0[1355]; 
    assign layer_1[2925] = layer_0[84]; 
    assign layer_1[2926] = layer_0[2407]; 
    assign layer_1[2927] = layer_0[3932] ^ layer_0[3826]; 
    assign layer_1[2928] = layer_0[3565]; 
    assign layer_1[2929] = ~layer_0[2871] | (layer_0[2945] & layer_0[2871]); 
    assign layer_1[2930] = layer_0[593] & ~layer_0[561]; 
    assign layer_1[2931] = ~layer_0[3941]; 
    assign layer_1[2932] = ~(layer_0[616] | layer_0[604]); 
    assign layer_1[2933] = layer_0[1347] & layer_0[1286]; 
    assign layer_1[2934] = ~layer_0[1009]; 
    assign layer_1[2935] = layer_0[1191] & ~layer_0[1215]; 
    assign layer_1[2936] = ~(layer_0[3338] & layer_0[3218]); 
    assign layer_1[2937] = layer_0[3467] ^ layer_0[3397]; 
    assign layer_1[2938] = layer_0[388] & ~layer_0[377]; 
    assign layer_1[2939] = layer_0[1350]; 
    assign layer_1[2940] = layer_0[3423] & ~layer_0[3460]; 
    assign layer_1[2941] = layer_0[3170]; 
    assign layer_1[2942] = ~(layer_0[5] ^ layer_0[51]); 
    assign layer_1[2943] = layer_0[571] & ~layer_0[579]; 
    assign layer_1[2944] = ~(layer_0[387] & layer_0[340]); 
    assign layer_1[2945] = layer_0[3367]; 
    assign layer_1[2946] = layer_0[1213] ^ layer_0[1335]; 
    assign layer_1[2947] = layer_0[189] & ~layer_0[253]; 
    assign layer_1[2948] = ~layer_0[2788] | (layer_0[2819] & layer_0[2788]); 
    assign layer_1[2949] = ~layer_0[1556] | (layer_0[1517] & layer_0[1556]); 
    assign layer_1[2950] = layer_0[1761] | layer_0[1818]; 
    assign layer_1[2951] = ~layer_0[3792] | (layer_0[3697] & layer_0[3792]); 
    assign layer_1[2952] = ~(layer_0[2494] | layer_0[2532]); 
    assign layer_1[2953] = ~layer_0[3700]; 
    assign layer_1[2954] = layer_0[955] | layer_0[949]; 
    assign layer_1[2955] = ~layer_0[3374] | (layer_0[3333] & layer_0[3374]); 
    assign layer_1[2956] = ~(layer_0[3303] | layer_0[3183]); 
    assign layer_1[2957] = ~layer_0[616]; 
    assign layer_1[2958] = ~(layer_0[540] | layer_0[501]); 
    assign layer_1[2959] = ~layer_0[999]; 
    assign layer_1[2960] = layer_0[2500] ^ layer_0[2514]; 
    assign layer_1[2961] = layer_0[2523] & layer_0[2553]; 
    assign layer_1[2962] = ~(layer_0[3371] & layer_0[3392]); 
    assign layer_1[2963] = layer_0[260]; 
    assign layer_1[2964] = layer_0[2671] ^ layer_0[2750]; 
    assign layer_1[2965] = layer_0[2260] | layer_0[2273]; 
    assign layer_1[2966] = layer_0[3441] & ~layer_0[3542]; 
    assign layer_1[2967] = layer_0[3458] | layer_0[3501]; 
    assign layer_1[2968] = layer_0[872] & layer_0[838]; 
    assign layer_1[2969] = ~layer_0[789] | (layer_0[870] & layer_0[789]); 
    assign layer_1[2970] = layer_0[2462]; 
    assign layer_1[2971] = ~layer_0[512] | (layer_0[512] & layer_0[426]); 
    assign layer_1[2972] = layer_0[1038] & ~layer_0[957]; 
    assign layer_1[2973] = layer_0[1035] ^ layer_0[957]; 
    assign layer_1[2974] = layer_0[1607] ^ layer_0[1626]; 
    assign layer_1[2975] = layer_0[2496] ^ layer_0[2450]; 
    assign layer_1[2976] = layer_0[411] ^ layer_0[435]; 
    assign layer_1[2977] = ~(layer_0[2874] ^ layer_0[2871]); 
    assign layer_1[2978] = ~layer_0[2793]; 
    assign layer_1[2979] = ~(layer_0[843] | layer_0[819]); 
    assign layer_1[2980] = ~layer_0[2654] | (layer_0[2654] & layer_0[2620]); 
    assign layer_1[2981] = layer_0[3900]; 
    assign layer_1[2982] = layer_0[2045] & layer_0[2151]; 
    assign layer_1[2983] = layer_0[1730] | layer_0[1811]; 
    assign layer_1[2984] = ~layer_0[2108] | (layer_0[2108] & layer_0[2154]); 
    assign layer_1[2985] = ~(layer_0[2690] & layer_0[2684]); 
    assign layer_1[2986] = layer_0[2897] & ~layer_0[2911]; 
    assign layer_1[2987] = layer_0[3487] & layer_0[3604]; 
    assign layer_1[2988] = layer_0[3312] | layer_0[3371]; 
    assign layer_1[2989] = ~layer_0[2906]; 
    assign layer_1[2990] = ~layer_0[3934]; 
    assign layer_1[2991] = ~layer_0[1753]; 
    assign layer_1[2992] = layer_0[794]; 
    assign layer_1[2993] = ~(layer_0[3486] | layer_0[3425]); 
    assign layer_1[2994] = layer_0[3322] ^ layer_0[3281]; 
    assign layer_1[2995] = ~layer_0[1690]; 
    assign layer_1[2996] = layer_0[2392] | layer_0[2291]; 
    assign layer_1[2997] = layer_0[3870] & ~layer_0[3839]; 
    assign layer_1[2998] = ~(layer_0[1649] | layer_0[1677]); 
    assign layer_1[2999] = layer_0[2668] & ~layer_0[2650]; 
    assign layer_1[3000] = layer_0[2187] ^ layer_0[2074]; 
    assign layer_1[3001] = layer_0[1979] & ~layer_0[1955]; 
    assign layer_1[3002] = ~(layer_0[121] & layer_0[134]); 
    assign layer_1[3003] = ~(layer_0[3286] ^ layer_0[3280]); 
    assign layer_1[3004] = layer_0[1427]; 
    assign layer_1[3005] = ~(layer_0[545] & layer_0[632]); 
    assign layer_1[3006] = ~(layer_0[3705] ^ layer_0[3607]); 
    assign layer_1[3007] = layer_0[2454] & ~layer_0[2461]; 
    assign layer_1[3008] = layer_0[520]; 
    assign layer_1[3009] = ~(layer_0[1085] | layer_0[1153]); 
    assign layer_1[3010] = ~layer_0[3619]; 
    assign layer_1[3011] = ~(layer_0[3843] & layer_0[3875]); 
    assign layer_1[3012] = ~layer_0[1276] | (layer_0[1276] & layer_0[1334]); 
    assign layer_1[3013] = ~(layer_0[859] ^ layer_0[842]); 
    assign layer_1[3014] = layer_0[2002] ^ layer_0[1948]; 
    assign layer_1[3015] = ~layer_0[751]; 
    assign layer_1[3016] = layer_0[2127] & ~layer_0[2042]; 
    assign layer_1[3017] = ~(layer_0[1776] | layer_0[1658]); 
    assign layer_1[3018] = ~(layer_0[333] & layer_0[254]); 
    assign layer_1[3019] = ~(layer_0[230] | layer_0[197]); 
    assign layer_1[3020] = layer_0[1979]; 
    assign layer_1[3021] = ~layer_0[3679]; 
    assign layer_1[3022] = ~layer_0[1134]; 
    assign layer_1[3023] = layer_0[222] ^ layer_0[158]; 
    assign layer_1[3024] = layer_0[3743] ^ layer_0[3790]; 
    assign layer_1[3025] = layer_0[2442]; 
    assign layer_1[3026] = layer_0[3624] | layer_0[3534]; 
    assign layer_1[3027] = ~(layer_0[3395] | layer_0[3322]); 
    assign layer_1[3028] = layer_0[2288]; 
    assign layer_1[3029] = layer_0[3973] | layer_0[3866]; 
    assign layer_1[3030] = ~layer_0[933]; 
    assign layer_1[3031] = layer_0[543] & ~layer_0[634]; 
    assign layer_1[3032] = layer_0[321] & ~layer_0[434]; 
    assign layer_1[3033] = layer_0[1900] & layer_0[2010]; 
    assign layer_1[3034] = ~(layer_0[2275] | layer_0[2149]); 
    assign layer_1[3035] = layer_0[194]; 
    assign layer_1[3036] = ~layer_0[1934] | (layer_0[1934] & layer_0[1991]); 
    assign layer_1[3037] = layer_0[1113]; 
    assign layer_1[3038] = layer_0[1165]; 
    assign layer_1[3039] = layer_0[443] & ~layer_0[506]; 
    assign layer_1[3040] = ~(layer_0[2307] | layer_0[2285]); 
    assign layer_1[3041] = layer_0[2355] | layer_0[2478]; 
    assign layer_1[3042] = ~layer_0[3290] | (layer_0[3175] & layer_0[3290]); 
    assign layer_1[3043] = layer_0[1087] | layer_0[1018]; 
    assign layer_1[3044] = layer_0[1953] & ~layer_0[2057]; 
    assign layer_1[3045] = ~(layer_0[2482] & layer_0[2421]); 
    assign layer_1[3046] = ~(layer_0[3188] & layer_0[3195]); 
    assign layer_1[3047] = layer_0[3765] & ~layer_0[3805]; 
    assign layer_1[3048] = ~layer_0[3820]; 
    assign layer_1[3049] = ~layer_0[849] | (layer_0[960] & layer_0[849]); 
    assign layer_1[3050] = layer_0[2730]; 
    assign layer_1[3051] = ~layer_0[88]; 
    assign layer_1[3052] = ~(layer_0[3095] ^ layer_0[3041]); 
    assign layer_1[3053] = layer_0[1966] & layer_0[2084]; 
    assign layer_1[3054] = layer_0[3692] & ~layer_0[3800]; 
    assign layer_1[3055] = ~layer_0[2769] | (layer_0[2850] & layer_0[2769]); 
    assign layer_1[3056] = layer_0[1281] & ~layer_0[1403]; 
    assign layer_1[3057] = layer_0[3017] & ~layer_0[3088]; 
    assign layer_1[3058] = layer_0[2276] & ~layer_0[2290]; 
    assign layer_1[3059] = layer_0[3533]; 
    assign layer_1[3060] = layer_0[3360] & ~layer_0[3302]; 
    assign layer_1[3061] = layer_0[688] & layer_0[808]; 
    assign layer_1[3062] = layer_0[3498] & ~layer_0[3452]; 
    assign layer_1[3063] = ~layer_0[3379]; 
    assign layer_1[3064] = ~layer_0[2962] | (layer_0[2962] & layer_0[3033]); 
    assign layer_1[3065] = ~layer_0[1642] | (layer_0[1576] & layer_0[1642]); 
    assign layer_1[3066] = ~(layer_0[3911] ^ layer_0[3872]); 
    assign layer_1[3067] = ~(layer_0[3806] & layer_0[3840]); 
    assign layer_1[3068] = ~(layer_0[2141] ^ layer_0[2137]); 
    assign layer_1[3069] = ~(layer_0[3177] | layer_0[3117]); 
    assign layer_1[3070] = ~(layer_0[3273] | layer_0[3172]); 
    assign layer_1[3071] = layer_0[713] ^ layer_0[742]; 
    assign layer_1[3072] = layer_0[239] & ~layer_0[277]; 
    assign layer_1[3073] = layer_0[730]; 
    assign layer_1[3074] = ~layer_0[3587] | (layer_0[3713] & layer_0[3587]); 
    assign layer_1[3075] = ~(layer_0[3174] ^ layer_0[3080]); 
    assign layer_1[3076] = layer_0[3100]; 
    assign layer_1[3077] = layer_0[515] & layer_0[623]; 
    assign layer_1[3078] = layer_0[1211] & ~layer_0[1093]; 
    assign layer_1[3079] = layer_0[1392]; 
    assign layer_1[3080] = ~layer_0[3936] | (layer_0[3936] & layer_0[3951]); 
    assign layer_1[3081] = layer_0[3676] ^ layer_0[3560]; 
    assign layer_1[3082] = ~(layer_0[1859] & layer_0[1738]); 
    assign layer_1[3083] = layer_0[771]; 
    assign layer_1[3084] = layer_0[2664] & ~layer_0[2588]; 
    assign layer_1[3085] = layer_0[1051] | layer_0[969]; 
    assign layer_1[3086] = layer_0[1069]; 
    assign layer_1[3087] = ~(layer_0[2976] & layer_0[2861]); 
    assign layer_1[3088] = ~(layer_0[2633] | layer_0[2550]); 
    assign layer_1[3089] = ~layer_0[129] | (layer_0[6] & layer_0[129]); 
    assign layer_1[3090] = ~layer_0[3800]; 
    assign layer_1[3091] = layer_0[453] & ~layer_0[581]; 
    assign layer_1[3092] = ~(layer_0[2031] | layer_0[1940]); 
    assign layer_1[3093] = layer_0[1131] ^ layer_0[1043]; 
    assign layer_1[3094] = ~layer_0[1677]; 
    assign layer_1[3095] = layer_0[737] ^ layer_0[759]; 
    assign layer_1[3096] = layer_0[1163] ^ layer_0[1116]; 
    assign layer_1[3097] = layer_0[825] | layer_0[793]; 
    assign layer_1[3098] = layer_0[3617]; 
    assign layer_1[3099] = ~layer_0[2634] | (layer_0[2706] & layer_0[2634]); 
    assign layer_1[3100] = ~(layer_0[634] | layer_0[554]); 
    assign layer_1[3101] = ~layer_0[2768] | (layer_0[2768] & layer_0[2832]); 
    assign layer_1[3102] = ~(layer_0[3393] ^ layer_0[3265]); 
    assign layer_1[3103] = ~layer_0[2455]; 
    assign layer_1[3104] = layer_0[1819] | layer_0[1888]; 
    assign layer_1[3105] = layer_0[1740]; 
    assign layer_1[3106] = ~layer_0[2845]; 
    assign layer_1[3107] = layer_0[241] | layer_0[165]; 
    assign layer_1[3108] = layer_0[3239]; 
    assign layer_1[3109] = ~(layer_0[2723] | layer_0[2686]); 
    assign layer_1[3110] = layer_0[2324]; 
    assign layer_1[3111] = ~(layer_0[1247] ^ layer_0[1133]); 
    assign layer_1[3112] = layer_0[598] & ~layer_0[668]; 
    assign layer_1[3113] = layer_0[1131] & ~layer_0[1119]; 
    assign layer_1[3114] = layer_0[1791]; 
    assign layer_1[3115] = ~layer_0[303] | (layer_0[303] & layer_0[230]); 
    assign layer_1[3116] = layer_0[1042]; 
    assign layer_1[3117] = ~layer_0[3030] | (layer_0[3030] & layer_0[3116]); 
    assign layer_1[3118] = ~layer_0[3144]; 
    assign layer_1[3119] = ~layer_0[3325]; 
    assign layer_1[3120] = ~(layer_0[2190] & layer_0[2072]); 
    assign layer_1[3121] = layer_0[2461] & layer_0[2337]; 
    assign layer_1[3122] = ~layer_0[1809] | (layer_0[1857] & layer_0[1809]); 
    assign layer_1[3123] = ~layer_0[2438]; 
    assign layer_1[3124] = ~layer_0[2970] | (layer_0[3017] & layer_0[2970]); 
    assign layer_1[3125] = layer_0[633] & layer_0[535]; 
    assign layer_1[3126] = layer_0[503] ^ layer_0[478]; 
    assign layer_1[3127] = ~layer_0[3820]; 
    assign layer_1[3128] = layer_0[2531]; 
    assign layer_1[3129] = ~layer_0[1185] | (layer_0[1185] & layer_0[1163]); 
    assign layer_1[3130] = layer_0[2327] ^ layer_0[2380]; 
    assign layer_1[3131] = ~layer_0[2148]; 
    assign layer_1[3132] = layer_0[102]; 
    assign layer_1[3133] = ~layer_0[249]; 
    assign layer_1[3134] = layer_0[977] & ~layer_0[1103]; 
    assign layer_1[3135] = layer_0[3863] & ~layer_0[3779]; 
    assign layer_1[3136] = layer_0[1308] ^ layer_0[1318]; 
    assign layer_1[3137] = ~(layer_0[2509] ^ layer_0[2636]); 
    assign layer_1[3138] = ~(layer_0[1518] | layer_0[1439]); 
    assign layer_1[3139] = ~(layer_0[1146] ^ layer_0[1181]); 
    assign layer_1[3140] = ~layer_0[3919]; 
    assign layer_1[3141] = layer_0[3120] ^ layer_0[3126]; 
    assign layer_1[3142] = ~(layer_0[3375] ^ layer_0[3252]); 
    assign layer_1[3143] = layer_0[2519] & layer_0[2464]; 
    assign layer_1[3144] = layer_0[2527] ^ layer_0[2446]; 
    assign layer_1[3145] = ~layer_0[3916]; 
    assign layer_1[3146] = ~(layer_0[778] | layer_0[666]); 
    assign layer_1[3147] = layer_0[2924] ^ layer_0[2921]; 
    assign layer_1[3148] = layer_0[1247] | layer_0[1370]; 
    assign layer_1[3149] = ~layer_0[548]; 
    assign layer_1[3150] = ~(layer_0[1447] & layer_0[1543]); 
    assign layer_1[3151] = ~(layer_0[2222] ^ layer_0[2175]); 
    assign layer_1[3152] = layer_0[137] | layer_0[17]; 
    assign layer_1[3153] = ~(layer_0[1354] ^ layer_0[1226]); 
    assign layer_1[3154] = layer_0[2006] ^ layer_0[1991]; 
    assign layer_1[3155] = layer_0[2621] & ~layer_0[2711]; 
    assign layer_1[3156] = ~layer_0[832]; 
    assign layer_1[3157] = layer_0[1756] & ~layer_0[1860]; 
    assign layer_1[3158] = ~layer_0[3714]; 
    assign layer_1[3159] = ~layer_0[1485] | (layer_0[1578] & layer_0[1485]); 
    assign layer_1[3160] = ~layer_0[3525] | (layer_0[3525] & layer_0[3471]); 
    assign layer_1[3161] = ~(layer_0[438] ^ layer_0[424]); 
    assign layer_1[3162] = layer_0[777] & ~layer_0[690]; 
    assign layer_1[3163] = layer_0[2114] & ~layer_0[2135]; 
    assign layer_1[3164] = layer_0[373] ^ layer_0[438]; 
    assign layer_1[3165] = layer_0[1738] & layer_0[1768]; 
    assign layer_1[3166] = layer_0[3637] & ~layer_0[3565]; 
    assign layer_1[3167] = ~(layer_0[2916] & layer_0[2989]); 
    assign layer_1[3168] = layer_0[3778] | layer_0[3790]; 
    assign layer_1[3169] = ~(layer_0[3573] | layer_0[3617]); 
    assign layer_1[3170] = layer_0[1089] & layer_0[1169]; 
    assign layer_1[3171] = ~layer_0[1821] | (layer_0[1719] & layer_0[1821]); 
    assign layer_1[3172] = layer_0[2467]; 
    assign layer_1[3173] = ~layer_0[3085]; 
    assign layer_1[3174] = ~(layer_0[528] ^ layer_0[432]); 
    assign layer_1[3175] = layer_0[1373] ^ layer_0[1333]; 
    assign layer_1[3176] = layer_0[194] | layer_0[168]; 
    assign layer_1[3177] = layer_0[1588] & layer_0[1581]; 
    assign layer_1[3178] = ~layer_0[2497]; 
    assign layer_1[3179] = layer_0[904] & ~layer_0[793]; 
    assign layer_1[3180] = layer_0[2037] ^ layer_0[2143]; 
    assign layer_1[3181] = layer_0[178] & layer_0[172]; 
    assign layer_1[3182] = ~layer_0[3515] | (layer_0[3515] & layer_0[3556]); 
    assign layer_1[3183] = ~layer_0[283] | (layer_0[283] & layer_0[381]); 
    assign layer_1[3184] = ~layer_0[454]; 
    assign layer_1[3185] = layer_0[551]; 
    assign layer_1[3186] = ~(layer_0[2392] & layer_0[2467]); 
    assign layer_1[3187] = layer_0[3644] & layer_0[3737]; 
    assign layer_1[3188] = layer_0[1474] & ~layer_0[1466]; 
    assign layer_1[3189] = ~(layer_0[2901] | layer_0[2955]); 
    assign layer_1[3190] = ~layer_0[1674]; 
    assign layer_1[3191] = ~(layer_0[619] | layer_0[716]); 
    assign layer_1[3192] = layer_0[1480] | layer_0[1356]; 
    assign layer_1[3193] = ~(layer_0[493] | layer_0[480]); 
    assign layer_1[3194] = ~(layer_0[2175] | layer_0[2151]); 
    assign layer_1[3195] = layer_0[798] & layer_0[735]; 
    assign layer_1[3196] = ~layer_0[3949] | (layer_0[3949] & layer_0[3961]); 
    assign layer_1[3197] = layer_0[2470] & ~layer_0[2459]; 
    assign layer_1[3198] = ~(layer_0[2074] ^ layer_0[1983]); 
    assign layer_1[3199] = ~(layer_0[2495] & layer_0[2461]); 
    assign layer_1[3200] = layer_0[300] & layer_0[389]; 
    assign layer_1[3201] = ~(layer_0[2796] | layer_0[2911]); 
    assign layer_1[3202] = ~layer_0[3911]; 
    assign layer_1[3203] = ~layer_0[2008] | (layer_0[2046] & layer_0[2008]); 
    assign layer_1[3204] = layer_0[1353] | layer_0[1426]; 
    assign layer_1[3205] = ~(layer_0[2234] & layer_0[2191]); 
    assign layer_1[3206] = ~layer_0[3029]; 
    assign layer_1[3207] = layer_0[1485] & ~layer_0[1502]; 
    assign layer_1[3208] = layer_0[3748] & ~layer_0[3623]; 
    assign layer_1[3209] = layer_0[2941]; 
    assign layer_1[3210] = layer_0[20] & ~layer_0[9]; 
    assign layer_1[3211] = ~layer_0[696]; 
    assign layer_1[3212] = ~layer_0[263]; 
    assign layer_1[3213] = ~(layer_0[497] ^ layer_0[516]); 
    assign layer_1[3214] = layer_0[1790] ^ layer_0[1811]; 
    assign layer_1[3215] = ~(layer_0[1321] & layer_0[1329]); 
    assign layer_1[3216] = layer_0[1615] & ~layer_0[1680]; 
    assign layer_1[3217] = layer_0[1540] & layer_0[1495]; 
    assign layer_1[3218] = ~(layer_0[2607] | layer_0[2542]); 
    assign layer_1[3219] = layer_0[2247] & layer_0[2250]; 
    assign layer_1[3220] = layer_0[2691]; 
    assign layer_1[3221] = ~(layer_0[3510] | layer_0[3385]); 
    assign layer_1[3222] = layer_0[15] | layer_0[78]; 
    assign layer_1[3223] = ~(layer_0[619] | layer_0[540]); 
    assign layer_1[3224] = ~layer_0[621] | (layer_0[621] & layer_0[652]); 
    assign layer_1[3225] = ~layer_0[582]; 
    assign layer_1[3226] = layer_0[894] & ~layer_0[852]; 
    assign layer_1[3227] = layer_0[2526] ^ layer_0[2613]; 
    assign layer_1[3228] = layer_0[159]; 
    assign layer_1[3229] = layer_0[2841] & layer_0[2854]; 
    assign layer_1[3230] = ~layer_0[3603]; 
    assign layer_1[3231] = layer_0[2702] ^ layer_0[2756]; 
    assign layer_1[3232] = layer_0[3221]; 
    assign layer_1[3233] = ~(layer_0[317] | layer_0[402]); 
    assign layer_1[3234] = ~layer_0[2182] | (layer_0[2197] & layer_0[2182]); 
    assign layer_1[3235] = layer_0[1834] & ~layer_0[1806]; 
    assign layer_1[3236] = ~(layer_0[3222] ^ layer_0[3273]); 
    assign layer_1[3237] = ~layer_0[1626]; 
    assign layer_1[3238] = layer_0[2506] ^ layer_0[2416]; 
    assign layer_1[3239] = ~layer_0[2067]; 
    assign layer_1[3240] = layer_0[3756] & ~layer_0[3826]; 
    assign layer_1[3241] = ~(layer_0[2089] & layer_0[2136]); 
    assign layer_1[3242] = layer_0[2953] ^ layer_0[3007]; 
    assign layer_1[3243] = ~(layer_0[3044] | layer_0[2941]); 
    assign layer_1[3244] = ~layer_0[143]; 
    assign layer_1[3245] = ~layer_0[3584] | (layer_0[3711] & layer_0[3584]); 
    assign layer_1[3246] = layer_0[2344]; 
    assign layer_1[3247] = layer_0[1776] ^ layer_0[1836]; 
    assign layer_1[3248] = ~(layer_0[3098] ^ layer_0[2980]); 
    assign layer_1[3249] = layer_0[501]; 
    assign layer_1[3250] = layer_0[1931]; 
    assign layer_1[3251] = ~layer_0[521] | (layer_0[497] & layer_0[521]); 
    assign layer_1[3252] = layer_0[3824]; 
    assign layer_1[3253] = ~layer_0[1107]; 
    assign layer_1[3254] = layer_0[3859]; 
    assign layer_1[3255] = layer_0[1282] | layer_0[1314]; 
    assign layer_1[3256] = ~layer_0[2969]; 
    assign layer_1[3257] = ~(layer_0[1992] ^ layer_0[1929]); 
    assign layer_1[3258] = layer_0[1362]; 
    assign layer_1[3259] = layer_0[3757]; 
    assign layer_1[3260] = ~layer_0[1347]; 
    assign layer_1[3261] = ~layer_0[2669]; 
    assign layer_1[3262] = layer_0[2631] | layer_0[2621]; 
    assign layer_1[3263] = ~layer_0[484]; 
    assign layer_1[3264] = ~layer_0[110]; 
    assign layer_1[3265] = layer_0[3334]; 
    assign layer_1[3266] = ~layer_0[310]; 
    assign layer_1[3267] = layer_0[3071]; 
    assign layer_1[3268] = ~(layer_0[2761] & layer_0[2873]); 
    assign layer_1[3269] = layer_0[2465]; 
    assign layer_1[3270] = ~layer_0[923] | (layer_0[923] & layer_0[1038]); 
    assign layer_1[3271] = layer_0[1398] ^ layer_0[1328]; 
    assign layer_1[3272] = ~layer_0[3511]; 
    assign layer_1[3273] = ~layer_0[1046]; 
    assign layer_1[3274] = layer_0[1007]; 
    assign layer_1[3275] = ~layer_0[2438]; 
    assign layer_1[3276] = layer_0[3625]; 
    assign layer_1[3277] = layer_0[130]; 
    assign layer_1[3278] = layer_0[1995]; 
    assign layer_1[3279] = ~(layer_0[1616] & layer_0[1614]); 
    assign layer_1[3280] = layer_0[290] | layer_0[390]; 
    assign layer_1[3281] = layer_0[1315]; 
    assign layer_1[3282] = layer_0[2710] | layer_0[2661]; 
    assign layer_1[3283] = layer_0[1246] & ~layer_0[1123]; 
    assign layer_1[3284] = layer_0[2684] | layer_0[2736]; 
    assign layer_1[3285] = layer_0[3201] & ~layer_0[3164]; 
    assign layer_1[3286] = ~layer_0[1798]; 
    assign layer_1[3287] = layer_0[664]; 
    assign layer_1[3288] = ~layer_0[1126]; 
    assign layer_1[3289] = layer_0[1752]; 
    assign layer_1[3290] = layer_0[2645]; 
    assign layer_1[3291] = layer_0[989]; 
    assign layer_1[3292] = layer_0[3297]; 
    assign layer_1[3293] = ~layer_0[3959]; 
    assign layer_1[3294] = ~layer_0[2063] | (layer_0[2063] & layer_0[2025]); 
    assign layer_1[3295] = ~layer_0[3274] | (layer_0[3274] & layer_0[3174]); 
    assign layer_1[3296] = layer_0[596]; 
    assign layer_1[3297] = ~layer_0[2608] | (layer_0[2703] & layer_0[2608]); 
    assign layer_1[3298] = layer_0[2976] ^ layer_0[2925]; 
    assign layer_1[3299] = layer_0[2277] & ~layer_0[2324]; 
    assign layer_1[3300] = ~(layer_0[1097] ^ layer_0[983]); 
    assign layer_1[3301] = layer_0[3197] & layer_0[3173]; 
    assign layer_1[3302] = ~layer_0[1670] | (layer_0[1798] & layer_0[1670]); 
    assign layer_1[3303] = layer_0[419]; 
    assign layer_1[3304] = layer_0[2825]; 
    assign layer_1[3305] = layer_0[2128] & ~layer_0[2093]; 
    assign layer_1[3306] = ~layer_0[3742]; 
    assign layer_1[3307] = layer_0[2531] & layer_0[2484]; 
    assign layer_1[3308] = ~layer_0[430]; 
    assign layer_1[3309] = layer_0[3806]; 
    assign layer_1[3310] = layer_0[1111]; 
    assign layer_1[3311] = layer_0[2110] ^ layer_0[2205]; 
    assign layer_1[3312] = ~(layer_0[1690] | layer_0[1798]); 
    assign layer_1[3313] = layer_0[2972] & layer_0[2868]; 
    assign layer_1[3314] = layer_0[1849] | layer_0[1973]; 
    assign layer_1[3315] = layer_0[1303] ^ layer_0[1293]; 
    assign layer_1[3316] = ~(layer_0[2009] ^ layer_0[1909]); 
    assign layer_1[3317] = ~(layer_0[2150] | layer_0[2246]); 
    assign layer_1[3318] = layer_0[505] | layer_0[417]; 
    assign layer_1[3319] = ~layer_0[1204] | (layer_0[1204] & layer_0[1217]); 
    assign layer_1[3320] = ~(layer_0[1010] | layer_0[1049]); 
    assign layer_1[3321] = layer_0[487] ^ layer_0[394]; 
    assign layer_1[3322] = layer_0[2120] ^ layer_0[2202]; 
    assign layer_1[3323] = ~(layer_0[3148] & layer_0[3234]); 
    assign layer_1[3324] = ~layer_0[1113] | (layer_0[1037] & layer_0[1113]); 
    assign layer_1[3325] = ~layer_0[856]; 
    assign layer_1[3326] = layer_0[371]; 
    assign layer_1[3327] = layer_0[3097] & layer_0[3210]; 
    assign layer_1[3328] = ~layer_0[1838] | (layer_0[1944] & layer_0[1838]); 
    assign layer_1[3329] = layer_0[327] ^ layer_0[246]; 
    assign layer_1[3330] = layer_0[3409] ^ layer_0[3518]; 
    assign layer_1[3331] = layer_0[2695]; 
    assign layer_1[3332] = layer_0[1985] & ~layer_0[1857]; 
    assign layer_1[3333] = ~layer_0[1841]; 
    assign layer_1[3334] = layer_0[614] | layer_0[664]; 
    assign layer_1[3335] = layer_0[720]; 
    assign layer_1[3336] = ~layer_0[3242]; 
    assign layer_1[3337] = layer_0[72] | layer_0[118]; 
    assign layer_1[3338] = layer_0[3976]; 
    assign layer_1[3339] = layer_0[2675] ^ layer_0[2654]; 
    assign layer_1[3340] = ~layer_0[171] | (layer_0[181] & layer_0[171]); 
    assign layer_1[3341] = layer_0[1596]; 
    assign layer_1[3342] = ~(layer_0[3466] ^ layer_0[3425]); 
    assign layer_1[3343] = ~(layer_0[994] ^ layer_0[874]); 
    assign layer_1[3344] = ~layer_0[3692] | (layer_0[3657] & layer_0[3692]); 
    assign layer_1[3345] = ~layer_0[2789] | (layer_0[2789] & layer_0[2911]); 
    assign layer_1[3346] = layer_0[1743] & ~layer_0[1623]; 
    assign layer_1[3347] = layer_0[3483] & ~layer_0[3450]; 
    assign layer_1[3348] = ~layer_0[1206] | (layer_0[1206] & layer_0[1114]); 
    assign layer_1[3349] = layer_0[1988] & layer_0[2063]; 
    assign layer_1[3350] = layer_0[3801] & ~layer_0[3821]; 
    assign layer_1[3351] = layer_0[3068] ^ layer_0[3108]; 
    assign layer_1[3352] = layer_0[2884] & layer_0[2880]; 
    assign layer_1[3353] = ~(layer_0[1721] | layer_0[1772]); 
    assign layer_1[3354] = layer_0[3494] & layer_0[3485]; 
    assign layer_1[3355] = layer_0[2493] & layer_0[2414]; 
    assign layer_1[3356] = layer_0[1386] & ~layer_0[1295]; 
    assign layer_1[3357] = layer_0[837] & ~layer_0[785]; 
    assign layer_1[3358] = ~(layer_0[3213] & layer_0[3196]); 
    assign layer_1[3359] = ~layer_0[658] | (layer_0[702] & layer_0[658]); 
    assign layer_1[3360] = layer_0[3575] | layer_0[3543]; 
    assign layer_1[3361] = layer_0[81]; 
    assign layer_1[3362] = layer_0[493] & ~layer_0[451]; 
    assign layer_1[3363] = layer_0[915]; 
    assign layer_1[3364] = ~layer_0[660] | (layer_0[660] & layer_0[534]); 
    assign layer_1[3365] = ~layer_0[927]; 
    assign layer_1[3366] = layer_0[3618] & ~layer_0[3652]; 
    assign layer_1[3367] = ~layer_0[1775]; 
    assign layer_1[3368] = ~layer_0[1931]; 
    assign layer_1[3369] = ~layer_0[2931] | (layer_0[2967] & layer_0[2931]); 
    assign layer_1[3370] = layer_0[366]; 
    assign layer_1[3371] = ~layer_0[3055] | (layer_0[3079] & layer_0[3055]); 
    assign layer_1[3372] = layer_0[3196]; 
    assign layer_1[3373] = ~(layer_0[2688] | layer_0[2758]); 
    assign layer_1[3374] = ~(layer_0[79] | layer_0[114]); 
    assign layer_1[3375] = layer_0[864] & ~layer_0[827]; 
    assign layer_1[3376] = layer_0[323] | layer_0[330]; 
    assign layer_1[3377] = ~layer_0[3772] | (layer_0[3772] & layer_0[3817]); 
    assign layer_1[3378] = ~(layer_0[2086] & layer_0[2161]); 
    assign layer_1[3379] = layer_0[1129] ^ layer_0[1214]; 
    assign layer_1[3380] = ~layer_0[2634] | (layer_0[2719] & layer_0[2634]); 
    assign layer_1[3381] = ~(layer_0[1708] & layer_0[1683]); 
    assign layer_1[3382] = layer_0[3747] & layer_0[3823]; 
    assign layer_1[3383] = ~layer_0[955]; 
    assign layer_1[3384] = ~layer_0[2005]; 
    assign layer_1[3385] = layer_0[513]; 
    assign layer_1[3386] = layer_0[3638] | layer_0[3681]; 
    assign layer_1[3387] = layer_0[1662] | layer_0[1599]; 
    assign layer_1[3388] = layer_0[1852] & layer_0[1885]; 
    assign layer_1[3389] = ~layer_0[3867]; 
    assign layer_1[3390] = ~(layer_0[1564] ^ layer_0[1496]); 
    assign layer_1[3391] = ~(layer_0[1427] ^ layer_0[1334]); 
    assign layer_1[3392] = layer_0[2915] | layer_0[2791]; 
    assign layer_1[3393] = layer_0[3847] & layer_0[3759]; 
    assign layer_1[3394] = layer_0[3301] | layer_0[3243]; 
    assign layer_1[3395] = ~layer_0[1753] | (layer_0[1798] & layer_0[1753]); 
    assign layer_1[3396] = ~layer_0[2652]; 
    assign layer_1[3397] = ~layer_0[3357] | (layer_0[3357] & layer_0[3230]); 
    assign layer_1[3398] = ~layer_0[3855]; 
    assign layer_1[3399] = ~(layer_0[2899] | layer_0[2989]); 
    assign layer_1[3400] = ~layer_0[1224]; 
    assign layer_1[3401] = ~(layer_0[3831] | layer_0[3761]); 
    assign layer_1[3402] = ~(layer_0[3376] & layer_0[3346]); 
    assign layer_1[3403] = layer_0[3711] | layer_0[3648]; 
    assign layer_1[3404] = ~layer_0[3019] | (layer_0[3019] & layer_0[3099]); 
    assign layer_1[3405] = ~layer_0[3064] | (layer_0[2957] & layer_0[3064]); 
    assign layer_1[3406] = layer_0[2100]; 
    assign layer_1[3407] = ~layer_0[2419] | (layer_0[2419] & layer_0[2522]); 
    assign layer_1[3408] = ~layer_0[2160] | (layer_0[2275] & layer_0[2160]); 
    assign layer_1[3409] = layer_0[2274]; 
    assign layer_1[3410] = ~(layer_0[429] | layer_0[355]); 
    assign layer_1[3411] = ~layer_0[3518] | (layer_0[3518] & layer_0[3613]); 
    assign layer_1[3412] = layer_0[3346]; 
    assign layer_1[3413] = ~layer_0[3520]; 
    assign layer_1[3414] = ~layer_0[673] | (layer_0[673] & layer_0[603]); 
    assign layer_1[3415] = ~layer_0[2442]; 
    assign layer_1[3416] = ~layer_0[3642]; 
    assign layer_1[3417] = ~(layer_0[1767] & layer_0[1751]); 
    assign layer_1[3418] = ~layer_0[1839]; 
    assign layer_1[3419] = ~(layer_0[935] & layer_0[926]); 
    assign layer_1[3420] = layer_0[3828]; 
    assign layer_1[3421] = layer_0[3859] & ~layer_0[3957]; 
    assign layer_1[3422] = layer_0[1453]; 
    assign layer_1[3423] = layer_0[890]; 
    assign layer_1[3424] = layer_0[3578]; 
    assign layer_1[3425] = layer_0[405]; 
    assign layer_1[3426] = layer_0[1813]; 
    assign layer_1[3427] = ~(layer_0[2933] ^ layer_0[2905]); 
    assign layer_1[3428] = ~layer_0[1006]; 
    assign layer_1[3429] = layer_0[917] & layer_0[795]; 
    assign layer_1[3430] = ~(layer_0[2587] | layer_0[2516]); 
    assign layer_1[3431] = layer_0[123] | layer_0[206]; 
    assign layer_1[3432] = ~(layer_0[1799] ^ layer_0[1926]); 
    assign layer_1[3433] = layer_0[2205]; 
    assign layer_1[3434] = ~(layer_0[3594] ^ layer_0[3505]); 
    assign layer_1[3435] = ~layer_0[1925]; 
    assign layer_1[3436] = ~(layer_0[3643] | layer_0[3550]); 
    assign layer_1[3437] = ~layer_0[3347]; 
    assign layer_1[3438] = ~(layer_0[783] & layer_0[680]); 
    assign layer_1[3439] = layer_0[3021] | layer_0[2964]; 
    assign layer_1[3440] = layer_0[1536] & ~layer_0[1413]; 
    assign layer_1[3441] = ~layer_0[2031]; 
    assign layer_1[3442] = layer_0[1016] ^ layer_0[897]; 
    assign layer_1[3443] = ~layer_0[2653]; 
    assign layer_1[3444] = ~layer_0[69]; 
    assign layer_1[3445] = layer_0[1054]; 
    assign layer_1[3446] = layer_0[1661]; 
    assign layer_1[3447] = ~(layer_0[1978] | layer_0[1982]); 
    assign layer_1[3448] = layer_0[2891] | layer_0[2984]; 
    assign layer_1[3449] = ~(layer_0[2646] | layer_0[2618]); 
    assign layer_1[3450] = layer_0[1351]; 
    assign layer_1[3451] = ~layer_0[2836]; 
    assign layer_1[3452] = layer_0[340] | layer_0[421]; 
    assign layer_1[3453] = layer_0[1235] & layer_0[1250]; 
    assign layer_1[3454] = ~(layer_0[2066] | layer_0[2054]); 
    assign layer_1[3455] = ~layer_0[1035] | (layer_0[1154] & layer_0[1035]); 
    assign layer_1[3456] = ~(layer_0[805] | layer_0[889]); 
    assign layer_1[3457] = layer_0[3683] ^ layer_0[3764]; 
    assign layer_1[3458] = ~(layer_0[1686] | layer_0[1765]); 
    assign layer_1[3459] = layer_0[28]; 
    assign layer_1[3460] = layer_0[2039]; 
    assign layer_1[3461] = ~layer_0[1473]; 
    assign layer_1[3462] = ~(layer_0[2838] & layer_0[2746]); 
    assign layer_1[3463] = ~layer_0[2272] | (layer_0[2272] & layer_0[2388]); 
    assign layer_1[3464] = layer_0[130] & ~layer_0[207]; 
    assign layer_1[3465] = layer_0[202] | layer_0[218]; 
    assign layer_1[3466] = layer_0[1142] & ~layer_0[1215]; 
    assign layer_1[3467] = ~(layer_0[240] | layer_0[259]); 
    assign layer_1[3468] = layer_0[1230]; 
    assign layer_1[3469] = ~(layer_0[2986] & layer_0[3076]); 
    assign layer_1[3470] = layer_0[1888] & ~layer_0[1858]; 
    assign layer_1[3471] = layer_0[3509] ^ layer_0[3580]; 
    assign layer_1[3472] = ~layer_0[476] | (layer_0[471] & layer_0[476]); 
    assign layer_1[3473] = ~layer_0[2449] | (layer_0[2547] & layer_0[2449]); 
    assign layer_1[3474] = ~layer_0[530] | (layer_0[530] & layer_0[437]); 
    assign layer_1[3475] = layer_0[2029] | layer_0[2001]; 
    assign layer_1[3476] = ~layer_0[1501]; 
    assign layer_1[3477] = ~(layer_0[2416] | layer_0[2319]); 
    assign layer_1[3478] = ~layer_0[1336] | (layer_0[1336] & layer_0[1242]); 
    assign layer_1[3479] = layer_0[3887] | layer_0[3935]; 
    assign layer_1[3480] = ~layer_0[1236]; 
    assign layer_1[3481] = ~(layer_0[1646] ^ layer_0[1577]); 
    assign layer_1[3482] = layer_0[187] & layer_0[190]; 
    assign layer_1[3483] = ~(layer_0[2972] ^ layer_0[2935]); 
    assign layer_1[3484] = ~layer_0[958]; 
    assign layer_1[3485] = layer_0[3147] ^ layer_0[3239]; 
    assign layer_1[3486] = ~layer_0[3150]; 
    assign layer_1[3487] = ~(layer_0[3080] | layer_0[2959]); 
    assign layer_1[3488] = ~(layer_0[1271] ^ layer_0[1327]); 
    assign layer_1[3489] = layer_0[2574] | layer_0[2462]; 
    assign layer_1[3490] = ~layer_0[2829]; 
    assign layer_1[3491] = layer_0[157] | layer_0[168]; 
    assign layer_1[3492] = layer_0[2001] | layer_0[1949]; 
    assign layer_1[3493] = ~(layer_0[2321] ^ layer_0[2264]); 
    assign layer_1[3494] = layer_0[2348] & ~layer_0[2453]; 
    assign layer_1[3495] = layer_0[2767] & ~layer_0[2674]; 
    assign layer_1[3496] = layer_0[1569]; 
    assign layer_1[3497] = layer_0[2975] | layer_0[2967]; 
    assign layer_1[3498] = ~layer_0[143]; 
    assign layer_1[3499] = layer_0[2494] | layer_0[2373]; 
    assign layer_1[3500] = ~(layer_0[2022] & layer_0[2041]); 
    assign layer_1[3501] = layer_0[3282] & layer_0[3171]; 
    assign layer_1[3502] = layer_0[898] & ~layer_0[968]; 
    assign layer_1[3503] = layer_0[2875] & ~layer_0[2970]; 
    assign layer_1[3504] = ~(layer_0[2520] ^ layer_0[2420]); 
    assign layer_1[3505] = ~(layer_0[629] | layer_0[720]); 
    assign layer_1[3506] = ~(layer_0[300] ^ layer_0[287]); 
    assign layer_1[3507] = layer_0[594]; 
    assign layer_1[3508] = layer_0[195]; 
    assign layer_1[3509] = layer_0[435]; 
    assign layer_1[3510] = layer_0[3626] | layer_0[3510]; 
    assign layer_1[3511] = layer_0[734]; 
    assign layer_1[3512] = ~layer_0[2603]; 
    assign layer_1[3513] = ~(layer_0[249] ^ layer_0[224]); 
    assign layer_1[3514] = ~layer_0[2462]; 
    assign layer_1[3515] = ~(layer_0[835] & layer_0[849]); 
    assign layer_1[3516] = ~layer_0[258]; 
    assign layer_1[3517] = ~(layer_0[3587] & layer_0[3661]); 
    assign layer_1[3518] = ~layer_0[3029]; 
    assign layer_1[3519] = ~layer_0[1352]; 
    assign layer_1[3520] = layer_0[3998]; 
    assign layer_1[3521] = ~(layer_0[601] ^ layer_0[541]); 
    assign layer_1[3522] = layer_0[2545]; 
    assign layer_1[3523] = layer_0[910] & layer_0[887]; 
    assign layer_1[3524] = ~layer_0[1210] | (layer_0[1210] & layer_0[1275]); 
    assign layer_1[3525] = ~(layer_0[1572] | layer_0[1451]); 
    assign layer_1[3526] = layer_0[2472] | layer_0[2489]; 
    assign layer_1[3527] = layer_0[3551]; 
    assign layer_1[3528] = ~(layer_0[904] | layer_0[919]); 
    assign layer_1[3529] = layer_0[2415]; 
    assign layer_1[3530] = ~(layer_0[3049] & layer_0[3047]); 
    assign layer_1[3531] = layer_0[3260]; 
    assign layer_1[3532] = layer_0[3659] ^ layer_0[3583]; 
    assign layer_1[3533] = ~layer_0[2305] | (layer_0[2290] & layer_0[2305]); 
    assign layer_1[3534] = ~layer_0[3067]; 
    assign layer_1[3535] = ~layer_0[3485]; 
    assign layer_1[3536] = layer_0[1305] & ~layer_0[1338]; 
    assign layer_1[3537] = layer_0[808] | layer_0[821]; 
    assign layer_1[3538] = layer_0[1198]; 
    assign layer_1[3539] = ~layer_0[1930]; 
    assign layer_1[3540] = ~layer_0[537]; 
    assign layer_1[3541] = ~layer_0[3701]; 
    assign layer_1[3542] = layer_0[2193] | layer_0[2106]; 
    assign layer_1[3543] = ~layer_0[730] | (layer_0[710] & layer_0[730]); 
    assign layer_1[3544] = ~(layer_0[1866] & layer_0[1782]); 
    assign layer_1[3545] = layer_0[2213]; 
    assign layer_1[3546] = layer_0[2137] & layer_0[2158]; 
    assign layer_1[3547] = layer_0[1815] & ~layer_0[1719]; 
    assign layer_1[3548] = layer_0[1126] & ~layer_0[1032]; 
    assign layer_1[3549] = layer_0[500] | layer_0[528]; 
    assign layer_1[3550] = ~(layer_0[1179] | layer_0[1178]); 
    assign layer_1[3551] = layer_0[2899] ^ layer_0[2894]; 
    assign layer_1[3552] = layer_0[1740] ^ layer_0[1668]; 
    assign layer_1[3553] = ~(layer_0[1999] ^ layer_0[2040]); 
    assign layer_1[3554] = ~layer_0[2022] | (layer_0[1894] & layer_0[2022]); 
    assign layer_1[3555] = ~layer_0[751] | (layer_0[741] & layer_0[751]); 
    assign layer_1[3556] = layer_0[2301]; 
    assign layer_1[3557] = ~(layer_0[1250] | layer_0[1300]); 
    assign layer_1[3558] = ~layer_0[95] | (layer_0[95] & layer_0[115]); 
    assign layer_1[3559] = layer_0[3723] & ~layer_0[3795]; 
    assign layer_1[3560] = layer_0[3367]; 
    assign layer_1[3561] = ~layer_0[223]; 
    assign layer_1[3562] = layer_0[1216]; 
    assign layer_1[3563] = layer_0[3393]; 
    assign layer_1[3564] = ~layer_0[1394]; 
    assign layer_1[3565] = layer_0[495]; 
    assign layer_1[3566] = ~(layer_0[3875] | layer_0[3799]); 
    assign layer_1[3567] = layer_0[62]; 
    assign layer_1[3568] = layer_0[1773] & ~layer_0[1771]; 
    assign layer_1[3569] = ~layer_0[2103]; 
    assign layer_1[3570] = ~layer_0[1413]; 
    assign layer_1[3571] = ~layer_0[827] | (layer_0[818] & layer_0[827]); 
    assign layer_1[3572] = ~layer_0[3242]; 
    assign layer_1[3573] = layer_0[1195] & ~layer_0[1094]; 
    assign layer_1[3574] = layer_0[2918] | layer_0[2838]; 
    assign layer_1[3575] = layer_0[1186]; 
    assign layer_1[3576] = ~(layer_0[352] ^ layer_0[438]); 
    assign layer_1[3577] = ~layer_0[812] | (layer_0[812] & layer_0[896]); 
    assign layer_1[3578] = ~layer_0[2833]; 
    assign layer_1[3579] = layer_0[3150]; 
    assign layer_1[3580] = layer_0[172]; 
    assign layer_1[3581] = ~(layer_0[2611] ^ layer_0[2507]); 
    assign layer_1[3582] = ~layer_0[3911]; 
    assign layer_1[3583] = layer_0[3687] & ~layer_0[3627]; 
    assign layer_1[3584] = ~layer_0[3953]; 
    assign layer_1[3585] = layer_0[1463]; 
    assign layer_1[3586] = ~(layer_0[2433] & layer_0[2335]); 
    assign layer_1[3587] = layer_0[770] | layer_0[868]; 
    assign layer_1[3588] = layer_0[941]; 
    assign layer_1[3589] = layer_0[1090] ^ layer_0[1130]; 
    assign layer_1[3590] = layer_0[739] ^ layer_0[729]; 
    assign layer_1[3591] = layer_0[927]; 
    assign layer_1[3592] = layer_0[760]; 
    assign layer_1[3593] = layer_0[1383] & ~layer_0[1397]; 
    assign layer_1[3594] = layer_0[643]; 
    assign layer_1[3595] = layer_0[1122] & ~layer_0[1068]; 
    assign layer_1[3596] = layer_0[1649]; 
    assign layer_1[3597] = ~(layer_0[1152] ^ layer_0[1245]); 
    assign layer_1[3598] = layer_0[843] & ~layer_0[791]; 
    assign layer_1[3599] = layer_0[2796] | layer_0[2746]; 
    assign layer_1[3600] = layer_0[2898]; 
    assign layer_1[3601] = ~(layer_0[616] | layer_0[628]); 
    assign layer_1[3602] = ~layer_0[29] | (layer_0[106] & layer_0[29]); 
    assign layer_1[3603] = ~(layer_0[2867] | layer_0[2890]); 
    assign layer_1[3604] = layer_0[3598] | layer_0[3620]; 
    assign layer_1[3605] = layer_0[3470] | layer_0[3540]; 
    assign layer_1[3606] = ~layer_0[2147]; 
    assign layer_1[3607] = layer_0[3536] & layer_0[3556]; 
    assign layer_1[3608] = layer_0[3913]; 
    assign layer_1[3609] = layer_0[404] & layer_0[346]; 
    assign layer_1[3610] = layer_0[708] & ~layer_0[726]; 
    assign layer_1[3611] = ~layer_0[3344]; 
    assign layer_1[3612] = layer_0[445]; 
    assign layer_1[3613] = ~layer_0[584] | (layer_0[584] & layer_0[539]); 
    assign layer_1[3614] = layer_0[2256]; 
    assign layer_1[3615] = ~(layer_0[275] ^ layer_0[279]); 
    assign layer_1[3616] = ~(layer_0[1732] | layer_0[1747]); 
    assign layer_1[3617] = ~layer_0[2805] | (layer_0[2805] & layer_0[2803]); 
    assign layer_1[3618] = layer_0[3438] | layer_0[3432]; 
    assign layer_1[3619] = layer_0[2265] & ~layer_0[2351]; 
    assign layer_1[3620] = layer_0[282]; 
    assign layer_1[3621] = layer_0[3428]; 
    assign layer_1[3622] = layer_0[455]; 
    assign layer_1[3623] = ~layer_0[3477] | (layer_0[3477] & layer_0[3448]); 
    assign layer_1[3624] = ~(layer_0[3486] | layer_0[3408]); 
    assign layer_1[3625] = layer_0[324] ^ layer_0[401]; 
    assign layer_1[3626] = layer_0[3078]; 
    assign layer_1[3627] = ~(layer_0[2981] ^ layer_0[2969]); 
    assign layer_1[3628] = ~(layer_0[3393] | layer_0[3340]); 
    assign layer_1[3629] = layer_0[1717] & ~layer_0[1609]; 
    assign layer_1[3630] = layer_0[1679] & layer_0[1646]; 
    assign layer_1[3631] = layer_0[3882]; 
    assign layer_1[3632] = layer_0[3319] | layer_0[3211]; 
    assign layer_1[3633] = ~layer_0[1544] | (layer_0[1442] & layer_0[1544]); 
    assign layer_1[3634] = ~layer_0[260] | (layer_0[260] & layer_0[315]); 
    assign layer_1[3635] = ~(layer_0[2139] | layer_0[2054]); 
    assign layer_1[3636] = layer_0[3252] & layer_0[3137]; 
    assign layer_1[3637] = layer_0[3007] & ~layer_0[3091]; 
    assign layer_1[3638] = ~layer_0[1725]; 
    assign layer_1[3639] = layer_0[662] | layer_0[711]; 
    assign layer_1[3640] = ~layer_0[1236] | (layer_0[1236] & layer_0[1327]); 
    assign layer_1[3641] = layer_0[556] & layer_0[679]; 
    assign layer_1[3642] = ~layer_0[1945]; 
    assign layer_1[3643] = layer_0[1198] & ~layer_0[1303]; 
    assign layer_1[3644] = ~(layer_0[2527] ^ layer_0[2419]); 
    assign layer_1[3645] = layer_0[1849] & layer_0[1925]; 
    assign layer_1[3646] = ~layer_0[2804] | (layer_0[2763] & layer_0[2804]); 
    assign layer_1[3647] = layer_0[1598]; 
    assign layer_1[3648] = ~layer_0[3822]; 
    assign layer_1[3649] = layer_0[1758] | layer_0[1738]; 
    assign layer_1[3650] = ~layer_0[3453]; 
    assign layer_1[3651] = ~(layer_0[3635] ^ layer_0[3510]); 
    assign layer_1[3652] = ~layer_0[2346]; 
    assign layer_1[3653] = ~layer_0[1534] | (layer_0[1534] & layer_0[1456]); 
    assign layer_1[3654] = ~(layer_0[3126] ^ layer_0[3169]); 
    assign layer_1[3655] = ~layer_0[28]; 
    assign layer_1[3656] = layer_0[2022] & ~layer_0[2113]; 
    assign layer_1[3657] = ~layer_0[1975]; 
    assign layer_1[3658] = layer_0[1786] ^ layer_0[1718]; 
    assign layer_1[3659] = layer_0[3134] | layer_0[3058]; 
    assign layer_1[3660] = ~layer_0[3717] | (layer_0[3717] & layer_0[3641]); 
    assign layer_1[3661] = ~(layer_0[448] | layer_0[495]); 
    assign layer_1[3662] = layer_0[724] & ~layer_0[716]; 
    assign layer_1[3663] = ~layer_0[627] | (layer_0[627] & layer_0[673]); 
    assign layer_1[3664] = ~(layer_0[2203] & layer_0[2274]); 
    assign layer_1[3665] = ~layer_0[3164] | (layer_0[3097] & layer_0[3164]); 
    assign layer_1[3666] = ~layer_0[2720]; 
    assign layer_1[3667] = ~layer_0[2594] | (layer_0[2594] & layer_0[2610]); 
    assign layer_1[3668] = ~layer_0[2099] | (layer_0[2099] & layer_0[2079]); 
    assign layer_1[3669] = ~layer_0[1589]; 
    assign layer_1[3670] = ~layer_0[275] | (layer_0[275] & layer_0[202]); 
    assign layer_1[3671] = ~(layer_0[3856] ^ layer_0[3760]); 
    assign layer_1[3672] = ~layer_0[3456] | (layer_0[3456] & layer_0[3465]); 
    assign layer_1[3673] = layer_0[1620] & ~layer_0[1536]; 
    assign layer_1[3674] = ~layer_0[1555]; 
    assign layer_1[3675] = layer_0[1897] & ~layer_0[1876]; 
    assign layer_1[3676] = ~(layer_0[561] | layer_0[490]); 
    assign layer_1[3677] = layer_0[1400] ^ layer_0[1358]; 
    assign layer_1[3678] = ~layer_0[3907]; 
    assign layer_1[3679] = layer_0[3956]; 
    assign layer_1[3680] = layer_0[1335] & ~layer_0[1345]; 
    assign layer_1[3681] = layer_0[5]; 
    assign layer_1[3682] = ~(layer_0[2958] & layer_0[3083]); 
    assign layer_1[3683] = ~layer_0[3202]; 
    assign layer_1[3684] = ~(layer_0[1153] & layer_0[1159]); 
    assign layer_1[3685] = ~layer_0[1932]; 
    assign layer_1[3686] = layer_0[2065]; 
    assign layer_1[3687] = layer_0[1945] | layer_0[1845]; 
    assign layer_1[3688] = ~layer_0[2938]; 
    assign layer_1[3689] = ~layer_0[372]; 
    assign layer_1[3690] = ~layer_0[624] | (layer_0[624] & layer_0[588]); 
    assign layer_1[3691] = layer_0[3983] & ~layer_0[3931]; 
    assign layer_1[3692] = layer_0[1348]; 
    assign layer_1[3693] = layer_0[1800] | layer_0[1849]; 
    assign layer_1[3694] = ~(layer_0[3550] ^ layer_0[3424]); 
    assign layer_1[3695] = layer_0[3231] & ~layer_0[3227]; 
    assign layer_1[3696] = layer_0[903]; 
    assign layer_1[3697] = layer_0[3542] ^ layer_0[3605]; 
    assign layer_1[3698] = layer_0[1277]; 
    assign layer_1[3699] = layer_0[2002] ^ layer_0[2094]; 
    assign layer_1[3700] = ~layer_0[2891]; 
    assign layer_1[3701] = ~layer_0[2358]; 
    assign layer_1[3702] = layer_0[3535] & ~layer_0[3486]; 
    assign layer_1[3703] = layer_0[2912] ^ layer_0[3020]; 
    assign layer_1[3704] = layer_0[1483] ^ layer_0[1557]; 
    assign layer_1[3705] = layer_0[1862] & layer_0[1906]; 
    assign layer_1[3706] = layer_0[2324] ^ layer_0[2387]; 
    assign layer_1[3707] = layer_0[1832] ^ layer_0[1844]; 
    assign layer_1[3708] = layer_0[1295] & layer_0[1176]; 
    assign layer_1[3709] = ~layer_0[2282]; 
    assign layer_1[3710] = ~layer_0[2698]; 
    assign layer_1[3711] = layer_0[1652] & ~layer_0[1778]; 
    assign layer_1[3712] = layer_0[3697]; 
    assign layer_1[3713] = ~(layer_0[2388] ^ layer_0[2478]); 
    assign layer_1[3714] = layer_0[2521] & layer_0[2480]; 
    assign layer_1[3715] = ~(layer_0[2874] & layer_0[2900]); 
    assign layer_1[3716] = layer_0[3788] & layer_0[3751]; 
    assign layer_1[3717] = layer_0[2940]; 
    assign layer_1[3718] = ~layer_0[3842]; 
    assign layer_1[3719] = layer_0[3243] ^ layer_0[3136]; 
    assign layer_1[3720] = ~(layer_0[3037] ^ layer_0[3065]); 
    assign layer_1[3721] = layer_0[382] ^ layer_0[267]; 
    assign layer_1[3722] = ~(layer_0[347] | layer_0[455]); 
    assign layer_1[3723] = ~layer_0[1315] | (layer_0[1295] & layer_0[1315]); 
    assign layer_1[3724] = layer_0[2289] | layer_0[2387]; 
    assign layer_1[3725] = ~layer_0[3086]; 
    assign layer_1[3726] = layer_0[165]; 
    assign layer_1[3727] = ~(layer_0[529] & layer_0[469]); 
    assign layer_1[3728] = layer_0[1381] | layer_0[1410]; 
    assign layer_1[3729] = ~(layer_0[94] ^ layer_0[179]); 
    assign layer_1[3730] = layer_0[1163]; 
    assign layer_1[3731] = ~layer_0[2843] | (layer_0[2843] & layer_0[2789]); 
    assign layer_1[3732] = layer_0[1084]; 
    assign layer_1[3733] = ~layer_0[2172]; 
    assign layer_1[3734] = layer_0[3327]; 
    assign layer_1[3735] = ~(layer_0[3249] ^ layer_0[3350]); 
    assign layer_1[3736] = layer_0[2195]; 
    assign layer_1[3737] = ~layer_0[1486]; 
    assign layer_1[3738] = layer_0[88]; 
    assign layer_1[3739] = ~layer_0[3803] | (layer_0[3803] & layer_0[3920]); 
    assign layer_1[3740] = ~(layer_0[384] ^ layer_0[502]); 
    assign layer_1[3741] = ~layer_0[2956] | (layer_0[3004] & layer_0[2956]); 
    assign layer_1[3742] = ~(layer_0[819] | layer_0[801]); 
    assign layer_1[3743] = layer_0[3888] & ~layer_0[3893]; 
    assign layer_1[3744] = layer_0[722] & ~layer_0[832]; 
    assign layer_1[3745] = ~layer_0[3879]; 
    assign layer_1[3746] = layer_0[2799]; 
    assign layer_1[3747] = ~layer_0[398]; 
    assign layer_1[3748] = layer_0[117]; 
    assign layer_1[3749] = layer_0[200]; 
    assign layer_1[3750] = layer_0[393] & ~layer_0[502]; 
    assign layer_1[3751] = ~(layer_0[2037] ^ layer_0[2026]); 
    assign layer_1[3752] = layer_0[1398]; 
    assign layer_1[3753] = ~layer_0[1487]; 
    assign layer_1[3754] = ~layer_0[1977] | (layer_0[1977] & layer_0[2041]); 
    assign layer_1[3755] = ~(layer_0[1861] ^ layer_0[1775]); 
    assign layer_1[3756] = ~layer_0[3750] | (layer_0[3725] & layer_0[3750]); 
    assign layer_1[3757] = layer_0[2702] | layer_0[2711]; 
    assign layer_1[3758] = layer_0[248] & ~layer_0[333]; 
    assign layer_1[3759] = layer_0[1947]; 
    assign layer_1[3760] = ~(layer_0[2468] | layer_0[2421]); 
    assign layer_1[3761] = layer_0[1302]; 
    assign layer_1[3762] = layer_0[2622]; 
    assign layer_1[3763] = layer_0[7] & layer_0[39]; 
    assign layer_1[3764] = ~layer_0[1410] | (layer_0[1410] & layer_0[1358]); 
    assign layer_1[3765] = ~layer_0[1497]; 
    assign layer_1[3766] = layer_0[3667] | layer_0[3755]; 
    assign layer_1[3767] = layer_0[1886] & ~layer_0[1789]; 
    assign layer_1[3768] = ~layer_0[2877]; 
    assign layer_1[3769] = layer_0[3862] | layer_0[3965]; 
    assign layer_1[3770] = layer_0[18] & ~layer_0[85]; 
    assign layer_1[3771] = layer_0[2878] & ~layer_0[2902]; 
    assign layer_1[3772] = layer_0[3000] & ~layer_0[3040]; 
    assign layer_1[3773] = layer_0[2288] | layer_0[2196]; 
    assign layer_1[3774] = ~(layer_0[2553] | layer_0[2504]); 
    assign layer_1[3775] = ~layer_0[534] | (layer_0[534] & layer_0[505]); 
    assign layer_1[3776] = layer_0[1410]; 
    assign layer_1[3777] = layer_0[3347]; 
    assign layer_1[3778] = ~layer_0[2014]; 
    assign layer_1[3779] = layer_0[138]; 
    assign layer_1[3780] = layer_0[884]; 
    assign layer_1[3781] = layer_0[1579]; 
    assign layer_1[3782] = layer_0[475] ^ layer_0[402]; 
    assign layer_1[3783] = ~layer_0[1101] | (layer_0[1101] & layer_0[1183]); 
    assign layer_1[3784] = layer_0[2875]; 
    assign layer_1[3785] = ~(layer_0[1752] ^ layer_0[1677]); 
    assign layer_1[3786] = ~layer_0[3585]; 
    assign layer_1[3787] = layer_0[2861]; 
    assign layer_1[3788] = ~(layer_0[3961] & layer_0[3936]); 
    assign layer_1[3789] = layer_0[1538] ^ layer_0[1590]; 
    assign layer_1[3790] = layer_0[3926]; 
    assign layer_1[3791] = ~(layer_0[174] ^ layer_0[281]); 
    assign layer_1[3792] = ~layer_0[3297]; 
    assign layer_1[3793] = ~layer_0[1716] | (layer_0[1833] & layer_0[1716]); 
    assign layer_1[3794] = layer_0[442] & ~layer_0[327]; 
    assign layer_1[3795] = layer_0[1925]; 
    assign layer_1[3796] = layer_0[1614] | layer_0[1699]; 
    assign layer_1[3797] = layer_0[1100] & layer_0[1102]; 
    assign layer_1[3798] = layer_0[3811] & ~layer_0[3740]; 
    assign layer_1[3799] = ~layer_0[3479] | (layer_0[3479] & layer_0[3573]); 
    assign layer_1[3800] = ~layer_0[780]; 
    assign layer_1[3801] = ~(layer_0[3935] | layer_0[3877]); 
    assign layer_1[3802] = ~(layer_0[3311] | layer_0[3217]); 
    assign layer_1[3803] = ~(layer_0[2884] ^ layer_0[2901]); 
    assign layer_1[3804] = layer_0[915] & ~layer_0[897]; 
    assign layer_1[3805] = ~layer_0[411]; 
    assign layer_1[3806] = layer_0[2941]; 
    assign layer_1[3807] = ~(layer_0[2508] & layer_0[2421]); 
    assign layer_1[3808] = ~(layer_0[790] ^ layer_0[740]); 
    assign layer_1[3809] = layer_0[3140] ^ layer_0[3033]; 
    assign layer_1[3810] = ~layer_0[2959]; 
    assign layer_1[3811] = layer_0[2712] & ~layer_0[2687]; 
    assign layer_1[3812] = ~(layer_0[1852] | layer_0[1874]); 
    assign layer_1[3813] = layer_0[666]; 
    assign layer_1[3814] = layer_0[3273] | layer_0[3296]; 
    assign layer_1[3815] = layer_0[2288] ^ layer_0[2394]; 
    assign layer_1[3816] = layer_0[412]; 
    assign layer_1[3817] = ~(layer_0[1458] ^ layer_0[1366]); 
    assign layer_1[3818] = ~layer_0[955]; 
    assign layer_1[3819] = ~layer_0[826]; 
    assign layer_1[3820] = ~(layer_0[2341] | layer_0[2229]); 
    assign layer_1[3821] = layer_0[2312] | layer_0[2395]; 
    assign layer_1[3822] = layer_0[1618] ^ layer_0[1638]; 
    assign layer_1[3823] = layer_0[2797] & ~layer_0[2924]; 
    assign layer_1[3824] = layer_0[3807]; 
    assign layer_1[3825] = ~(layer_0[1971] | layer_0[1985]); 
    assign layer_1[3826] = ~(layer_0[3987] ^ layer_0[3962]); 
    assign layer_1[3827] = ~layer_0[180] | (layer_0[180] & layer_0[70]); 
    assign layer_1[3828] = ~layer_0[3824]; 
    assign layer_1[3829] = ~(layer_0[3720] ^ layer_0[3739]); 
    assign layer_1[3830] = layer_0[3894] & ~layer_0[3867]; 
    assign layer_1[3831] = layer_0[1240]; 
    assign layer_1[3832] = ~(layer_0[1787] ^ layer_0[1709]); 
    assign layer_1[3833] = ~(layer_0[2684] ^ layer_0[2762]); 
    assign layer_1[3834] = ~(layer_0[1634] ^ layer_0[1612]); 
    assign layer_1[3835] = layer_0[2006] & ~layer_0[2032]; 
    assign layer_1[3836] = ~(layer_0[3260] & layer_0[3282]); 
    assign layer_1[3837] = ~layer_0[2907]; 
    assign layer_1[3838] = ~layer_0[623]; 
    assign layer_1[3839] = ~layer_0[2619] | (layer_0[2619] & layer_0[2596]); 
    assign layer_1[3840] = layer_0[2470] & layer_0[2371]; 
    assign layer_1[3841] = ~layer_0[1477]; 
    assign layer_1[3842] = ~layer_0[936]; 
    assign layer_1[3843] = ~layer_0[3679]; 
    assign layer_1[3844] = layer_0[3011] & ~layer_0[2984]; 
    assign layer_1[3845] = layer_0[3411] & ~layer_0[3388]; 
    assign layer_1[3846] = layer_0[1224] & ~layer_0[1143]; 
    assign layer_1[3847] = ~layer_0[2861]; 
    assign layer_1[3848] = ~layer_0[87] | (layer_0[87] & layer_0[121]); 
    assign layer_1[3849] = ~layer_0[2808]; 
    assign layer_1[3850] = ~layer_0[3039] | (layer_0[2926] & layer_0[3039]); 
    assign layer_1[3851] = ~layer_0[1048] | (layer_0[1048] & layer_0[1095]); 
    assign layer_1[3852] = ~layer_0[625] | (layer_0[625] & layer_0[729]); 
    assign layer_1[3853] = ~layer_0[3966]; 
    assign layer_1[3854] = ~layer_0[1065]; 
    assign layer_1[3855] = ~layer_0[3148] | (layer_0[3076] & layer_0[3148]); 
    assign layer_1[3856] = ~layer_0[2914]; 
    assign layer_1[3857] = ~(layer_0[3165] ^ layer_0[3242]); 
    assign layer_1[3858] = ~layer_0[1088]; 
    assign layer_1[3859] = layer_0[842] & layer_0[807]; 
    assign layer_1[3860] = ~(layer_0[903] ^ layer_0[825]); 
    assign layer_1[3861] = layer_0[3115] & ~layer_0[3198]; 
    assign layer_1[3862] = layer_0[3001] | layer_0[2963]; 
    assign layer_1[3863] = layer_0[165] | layer_0[233]; 
    assign layer_1[3864] = layer_0[836]; 
    assign layer_1[3865] = ~layer_0[212] | (layer_0[108] & layer_0[212]); 
    assign layer_1[3866] = layer_0[3227] | layer_0[3190]; 
    assign layer_1[3867] = ~layer_0[3172]; 
    assign layer_1[3868] = ~layer_0[3387]; 
    assign layer_1[3869] = ~(layer_0[902] | layer_0[969]); 
    assign layer_1[3870] = ~layer_0[1664] | (layer_0[1575] & layer_0[1664]); 
    assign layer_1[3871] = layer_0[2409] & ~layer_0[2420]; 
    assign layer_1[3872] = layer_0[942] & ~layer_0[895]; 
    assign layer_1[3873] = layer_0[3631] & ~layer_0[3603]; 
    assign layer_1[3874] = ~(layer_0[1306] ^ layer_0[1251]); 
    assign layer_1[3875] = ~layer_0[3672]; 
    assign layer_1[3876] = ~layer_0[2339]; 
    assign layer_1[3877] = ~layer_0[1821]; 
    assign layer_1[3878] = layer_0[2947] & ~layer_0[3048]; 
    assign layer_1[3879] = ~layer_0[2525]; 
    assign layer_1[3880] = layer_0[2696] ^ layer_0[2776]; 
    assign layer_1[3881] = ~layer_0[3191] | (layer_0[3230] & layer_0[3191]); 
    assign layer_1[3882] = ~(layer_0[893] ^ layer_0[844]); 
    assign layer_1[3883] = layer_0[1239] ^ layer_0[1363]; 
    assign layer_1[3884] = ~layer_0[1563]; 
    assign layer_1[3885] = layer_0[2716] & ~layer_0[2645]; 
    assign layer_1[3886] = ~layer_0[146] | (layer_0[147] & layer_0[146]); 
    assign layer_1[3887] = ~layer_0[862]; 
    assign layer_1[3888] = ~layer_0[1066]; 
    assign layer_1[3889] = layer_0[1166]; 
    assign layer_1[3890] = ~layer_0[2492] | (layer_0[2492] & layer_0[2600]); 
    assign layer_1[3891] = ~layer_0[3083]; 
    assign layer_1[3892] = layer_0[447]; 
    assign layer_1[3893] = layer_0[3175] & ~layer_0[3269]; 
    assign layer_1[3894] = layer_0[999]; 
    assign layer_1[3895] = layer_0[125]; 
    assign layer_1[3896] = layer_0[1335]; 
    assign layer_1[3897] = ~(layer_0[676] ^ layer_0[636]); 
    assign layer_1[3898] = layer_0[3914] & ~layer_0[3829]; 
    assign layer_1[3899] = ~layer_0[2811] | (layer_0[2760] & layer_0[2811]); 
    assign layer_1[3900] = ~layer_0[2697]; 
    assign layer_1[3901] = layer_0[1138]; 
    assign layer_1[3902] = layer_0[3970]; 
    assign layer_1[3903] = layer_0[3817] & layer_0[3825]; 
    assign layer_1[3904] = layer_0[2315]; 
    assign layer_1[3905] = layer_0[21]; 
    assign layer_1[3906] = layer_0[2743]; 
    assign layer_1[3907] = layer_0[704]; 
    assign layer_1[3908] = layer_0[3776] & ~layer_0[3702]; 
    assign layer_1[3909] = ~(layer_0[2633] ^ layer_0[2721]); 
    assign layer_1[3910] = ~layer_0[2549]; 
    assign layer_1[3911] = layer_0[1299] & ~layer_0[1230]; 
    assign layer_1[3912] = layer_0[2818]; 
    assign layer_1[3913] = layer_0[1875] ^ layer_0[1944]; 
    assign layer_1[3914] = layer_0[166] & ~layer_0[190]; 
    assign layer_1[3915] = ~layer_0[3273]; 
    assign layer_1[3916] = ~layer_0[95] | (layer_0[91] & layer_0[95]); 
    assign layer_1[3917] = ~(layer_0[1538] & layer_0[1532]); 
    assign layer_1[3918] = layer_0[2309] | layer_0[2209]; 
    assign layer_1[3919] = layer_0[1153] | layer_0[1069]; 
    assign layer_1[3920] = ~layer_0[3922] | (layer_0[3843] & layer_0[3922]); 
    assign layer_1[3921] = layer_0[2665]; 
    assign layer_1[3922] = layer_0[2771]; 
    assign layer_1[3923] = layer_0[1636] & ~layer_0[1738]; 
    assign layer_1[3924] = layer_0[3224] & ~layer_0[3099]; 
    assign layer_1[3925] = layer_0[1605] & layer_0[1544]; 
    assign layer_1[3926] = ~layer_0[1575]; 
    assign layer_1[3927] = ~layer_0[283] | (layer_0[183] & layer_0[283]); 
    assign layer_1[3928] = ~layer_0[213]; 
    assign layer_1[3929] = ~(layer_0[778] ^ layer_0[699]); 
    assign layer_1[3930] = ~(layer_0[2677] & layer_0[2784]); 
    assign layer_1[3931] = layer_0[187]; 
    assign layer_1[3932] = layer_0[949] | layer_0[925]; 
    assign layer_1[3933] = ~layer_0[1837] | (layer_0[1837] & layer_0[1814]); 
    assign layer_1[3934] = layer_0[385] & layer_0[412]; 
    assign layer_1[3935] = layer_0[3417] | layer_0[3410]; 
    assign layer_1[3936] = ~(layer_0[3353] ^ layer_0[3226]); 
    assign layer_1[3937] = layer_0[2858] & ~layer_0[2903]; 
    assign layer_1[3938] = ~(layer_0[1318] | layer_0[1320]); 
    assign layer_1[3939] = ~layer_0[3789]; 
    assign layer_1[3940] = ~(layer_0[2089] ^ layer_0[1967]); 
    assign layer_1[3941] = layer_0[554] & ~layer_0[551]; 
    assign layer_1[3942] = layer_0[1328] & layer_0[1321]; 
    assign layer_1[3943] = ~layer_0[3537]; 
    assign layer_1[3944] = ~layer_0[426] | (layer_0[426] & layer_0[478]); 
    assign layer_1[3945] = ~layer_0[956]; 
    assign layer_1[3946] = ~layer_0[1212]; 
    assign layer_1[3947] = ~layer_0[1228] | (layer_0[1228] & layer_0[1102]); 
    assign layer_1[3948] = layer_0[2175] | layer_0[2116]; 
    assign layer_1[3949] = layer_0[2348] ^ layer_0[2333]; 
    assign layer_1[3950] = layer_0[3568] & ~layer_0[3563]; 
    assign layer_1[3951] = ~layer_0[3258]; 
    assign layer_1[3952] = layer_0[1878] & ~layer_0[1958]; 
    assign layer_1[3953] = layer_0[3911] & ~layer_0[3785]; 
    assign layer_1[3954] = ~layer_0[1978]; 
    assign layer_1[3955] = layer_0[2504]; 
    assign layer_1[3956] = layer_0[1502] | layer_0[1400]; 
    assign layer_1[3957] = ~(layer_0[20] ^ layer_0[44]); 
    assign layer_1[3958] = ~layer_0[3848]; 
    assign layer_1[3959] = ~layer_0[3582]; 
    assign layer_1[3960] = ~layer_0[287] | (layer_0[178] & layer_0[287]); 
    assign layer_1[3961] = layer_0[2028] | layer_0[2128]; 
    assign layer_1[3962] = layer_0[2498] ^ layer_0[2593]; 
    assign layer_1[3963] = ~layer_0[557] | (layer_0[604] & layer_0[557]); 
    assign layer_1[3964] = ~(layer_0[82] & layer_0[9]); 
    assign layer_1[3965] = layer_0[1822] & ~layer_0[1737]; 
    assign layer_1[3966] = layer_0[1433]; 
    assign layer_1[3967] = layer_0[2510] | layer_0[2430]; 
    assign layer_1[3968] = layer_0[1238] & ~layer_0[1305]; 
    assign layer_1[3969] = layer_0[960] & ~layer_0[842]; 
    assign layer_1[3970] = ~(layer_0[103] & layer_0[50]); 
    assign layer_1[3971] = layer_0[1761] ^ layer_0[1879]; 
    assign layer_1[3972] = layer_0[3998] & layer_0[3898]; 
    assign layer_1[3973] = layer_0[1976]; 
    assign layer_1[3974] = layer_0[557] & ~layer_0[541]; 
    assign layer_1[3975] = ~layer_0[2588]; 
    assign layer_1[3976] = layer_0[932] & layer_0[937]; 
    assign layer_1[3977] = layer_0[1326] | layer_0[1224]; 
    assign layer_1[3978] = ~(layer_0[1303] ^ layer_0[1227]); 
    assign layer_1[3979] = ~layer_0[1906]; 
    assign layer_1[3980] = ~layer_0[3638]; 
    assign layer_1[3981] = ~layer_0[2858]; 
    assign layer_1[3982] = ~(layer_0[1366] ^ layer_0[1479]); 
    assign layer_1[3983] = layer_0[3259] & ~layer_0[3136]; 
    assign layer_1[3984] = layer_0[1484] ^ layer_0[1476]; 
    assign layer_1[3985] = layer_0[3879] & ~layer_0[3973]; 
    assign layer_1[3986] = layer_0[2955] & layer_0[2994]; 
    assign layer_1[3987] = layer_0[3190] | layer_0[3198]; 
    assign layer_1[3988] = layer_0[764] ^ layer_0[706]; 
    assign layer_1[3989] = layer_0[2571] & layer_0[2522]; 
    assign layer_1[3990] = ~layer_0[2231]; 
    assign layer_1[3991] = layer_0[2493] & ~layer_0[2379]; 
    assign layer_1[3992] = layer_0[1402]; 
    assign layer_1[3993] = layer_0[296]; 
    assign layer_1[3994] = ~layer_0[827] | (layer_0[827] & layer_0[860]); 
    assign layer_1[3995] = ~(layer_0[2867] ^ layer_0[2830]); 
    assign layer_1[3996] = ~layer_0[1735]; 
    assign layer_1[3997] = layer_0[2829]; 
    assign layer_1[3998] = ~layer_0[1714]; 
    assign layer_1[3999] = layer_0[172] & ~layer_0[59]; 
    // Layer 2 ============================================================
    assign out[0] = layer_1[1290] & ~layer_1[1231]; 
    assign out[1] = layer_1[2480] & layer_1[2459]; 
    assign out[2] = layer_1[531] & ~layer_1[438]; 
    assign out[3] = ~layer_1[1692]; 
    assign out[4] = layer_1[2150]; 
    assign out[5] = layer_1[646] & ~layer_1[755]; 
    assign out[6] = layer_1[978] ^ layer_1[1105]; 
    assign out[7] = ~layer_1[1361]; 
    assign out[8] = ~(layer_1[3726] ^ layer_1[3609]); 
    assign out[9] = layer_1[2202] & layer_1[2254]; 
    assign out[10] = ~layer_1[3761] | (layer_1[3761] & layer_1[3854]); 
    assign out[11] = ~(layer_1[343] | layer_1[413]); 
    assign out[12] = ~(layer_1[2842] ^ layer_1[2775]); 
    assign out[13] = ~layer_1[3922]; 
    assign out[14] = ~layer_1[2834] | (layer_1[2909] & layer_1[2834]); 
    assign out[15] = ~layer_1[2981]; 
    assign out[16] = ~(layer_1[1850] | layer_1[1761]); 
    assign out[17] = layer_1[3687] & ~layer_1[3635]; 
    assign out[18] = layer_1[873] ^ layer_1[954]; 
    assign out[19] = ~(layer_1[1520] & layer_1[1430]); 
    assign out[20] = ~layer_1[1535]; 
    assign out[21] = layer_1[3214] | layer_1[3238]; 
    assign out[22] = layer_1[2511]; 
    assign out[23] = layer_1[461]; 
    assign out[24] = layer_1[3103] & layer_1[3048]; 
    assign out[25] = layer_1[3177] ^ layer_1[3156]; 
    assign out[26] = ~(layer_1[2203] | layer_1[2312]); 
    assign out[27] = ~(layer_1[1296] ^ layer_1[1289]); 
    assign out[28] = layer_1[1256]; 
    assign out[29] = layer_1[2413]; 
    assign out[30] = ~(layer_1[2263] | layer_1[2312]); 
    assign out[31] = ~layer_1[3107]; 
    assign out[32] = layer_1[7] & ~layer_1[110]; 
    assign out[33] = ~layer_1[3657]; 
    assign out[34] = ~(layer_1[420] ^ layer_1[532]); 
    assign out[35] = layer_1[2079] & ~layer_1[2027]; 
    assign out[36] = ~(layer_1[3033] ^ layer_1[2963]); 
    assign out[37] = layer_1[3287]; 
    assign out[38] = ~layer_1[1265] | (layer_1[1265] & layer_1[1168]); 
    assign out[39] = ~layer_1[1200]; 
    assign out[40] = layer_1[175]; 
    assign out[41] = layer_1[2328]; 
    assign out[42] = layer_1[3577] & layer_1[3499]; 
    assign out[43] = layer_1[2578] & ~layer_1[2450]; 
    assign out[44] = ~(layer_1[2080] & layer_1[2061]); 
    assign out[45] = layer_1[2279] | layer_1[2336]; 
    assign out[46] = layer_1[600] & ~layer_1[682]; 
    assign out[47] = layer_1[1552] ^ layer_1[1548]; 
    assign out[48] = ~layer_1[2801]; 
    assign out[49] = layer_1[2577] & layer_1[2705]; 
    assign out[50] = ~layer_1[990] | (layer_1[1082] & layer_1[990]); 
    assign out[51] = ~(layer_1[3799] ^ layer_1[3785]); 
    assign out[52] = ~layer_1[2958]; 
    assign out[53] = layer_1[2513]; 
    assign out[54] = ~(layer_1[3381] | layer_1[3339]); 
    assign out[55] = layer_1[3612] ^ layer_1[3690]; 
    assign out[56] = ~layer_1[386]; 
    assign out[57] = layer_1[1771] & ~layer_1[1850]; 
    assign out[58] = ~layer_1[826] | (layer_1[869] & layer_1[826]); 
    assign out[59] = ~layer_1[1125]; 
    assign out[60] = ~(layer_1[3468] ^ layer_1[3581]); 
    assign out[61] = layer_1[870] & ~layer_1[840]; 
    assign out[62] = layer_1[2164] & layer_1[2209]; 
    assign out[63] = ~layer_1[3489]; 
    assign out[64] = layer_1[27] & ~layer_1[88]; 
    assign out[65] = ~(layer_1[1064] ^ layer_1[1009]); 
    assign out[66] = layer_1[776] & ~layer_1[811]; 
    assign out[67] = ~(layer_1[1064] ^ layer_1[1167]); 
    assign out[68] = ~(layer_1[2401] ^ layer_1[2286]); 
    assign out[69] = layer_1[1823] & layer_1[1709]; 
    assign out[70] = layer_1[2322]; 
    assign out[71] = layer_1[2782]; 
    assign out[72] = ~layer_1[912]; 
    assign out[73] = layer_1[3525] & ~layer_1[3615]; 
    assign out[74] = ~layer_1[3638]; 
    assign out[75] = layer_1[1409]; 
    assign out[76] = ~layer_1[2640]; 
    assign out[77] = ~layer_1[682]; 
    assign out[78] = ~(layer_1[2647] & layer_1[2529]); 
    assign out[79] = layer_1[3221] & ~layer_1[3228]; 
    assign out[80] = ~(layer_1[1659] ^ layer_1[1614]); 
    assign out[81] = layer_1[378]; 
    assign out[82] = ~layer_1[1529]; 
    assign out[83] = layer_1[2118]; 
    assign out[84] = layer_1[2644] ^ layer_1[2741]; 
    assign out[85] = layer_1[502]; 
    assign out[86] = layer_1[1623]; 
    assign out[87] = ~layer_1[1936]; 
    assign out[88] = layer_1[3116] ^ layer_1[3067]; 
    assign out[89] = ~layer_1[3400] | (layer_1[3400] & layer_1[3498]); 
    assign out[90] = ~layer_1[1289]; 
    assign out[91] = ~(layer_1[1689] ^ layer_1[1595]); 
    assign out[92] = ~layer_1[976]; 
    assign out[93] = ~layer_1[1736]; 
    assign out[94] = ~(layer_1[3792] ^ layer_1[3785]); 
    assign out[95] = ~layer_1[2948]; 
    assign out[96] = ~(layer_1[2839] | layer_1[2714]); 
    assign out[97] = ~layer_1[256] | (layer_1[256] & layer_1[376]); 
    assign out[98] = ~(layer_1[1863] ^ layer_1[1910]); 
    assign out[99] = ~(layer_1[539] ^ layer_1[521]); 
    assign out[100] = ~(layer_1[3712] ^ layer_1[3656]); 
    assign out[101] = layer_1[1441]; 
    assign out[102] = ~(layer_1[1108] ^ layer_1[1032]); 
    assign out[103] = layer_1[488] ^ layer_1[402]; 
    assign out[104] = ~layer_1[1315]; 
    assign out[105] = ~(layer_1[2228] ^ layer_1[2316]); 
    assign out[106] = layer_1[2771] & layer_1[2820]; 
    assign out[107] = ~layer_1[3562] | (layer_1[3562] & layer_1[3652]); 
    assign out[108] = layer_1[2234] & layer_1[2331]; 
    assign out[109] = layer_1[2830]; 
    assign out[110] = layer_1[2296]; 
    assign out[111] = ~(layer_1[2194] ^ layer_1[2069]); 
    assign out[112] = layer_1[1016]; 
    assign out[113] = ~(layer_1[2007] ^ layer_1[1954]); 
    assign out[114] = ~layer_1[768]; 
    assign out[115] = layer_1[2190] ^ layer_1[2072]; 
    assign out[116] = ~layer_1[1964]; 
    assign out[117] = ~layer_1[1996]; 
    assign out[118] = ~(layer_1[993] & layer_1[1011]); 
    assign out[119] = layer_1[1411]; 
    assign out[120] = layer_1[510]; 
    assign out[121] = layer_1[1049] & ~layer_1[1047]; 
    assign out[122] = ~layer_1[3121]; 
    assign out[123] = layer_1[702] ^ layer_1[602]; 
    assign out[124] = ~layer_1[2181]; 
    assign out[125] = ~(layer_1[3543] ^ layer_1[3512]); 
    assign out[126] = ~(layer_1[1419] ^ layer_1[1494]); 
    assign out[127] = ~layer_1[712]; 
    assign out[128] = ~(layer_1[992] ^ layer_1[886]); 
    assign out[129] = layer_1[2812] & ~layer_1[2859]; 
    assign out[130] = layer_1[171] & layer_1[212]; 
    assign out[131] = layer_1[3855]; 
    assign out[132] = ~layer_1[627]; 
    assign out[133] = ~layer_1[3489]; 
    assign out[134] = layer_1[282] & ~layer_1[261]; 
    assign out[135] = ~layer_1[836]; 
    assign out[136] = ~layer_1[2545]; 
    assign out[137] = layer_1[3424] & ~layer_1[3338]; 
    assign out[138] = ~(layer_1[3234] & layer_1[3227]); 
    assign out[139] = ~(layer_1[616] | layer_1[505]); 
    assign out[140] = ~(layer_1[922] | layer_1[1048]); 
    assign out[141] = ~(layer_1[2623] ^ layer_1[2692]); 
    assign out[142] = ~layer_1[3779]; 
    assign out[143] = layer_1[2347]; 
    assign out[144] = ~layer_1[428]; 
    assign out[145] = ~layer_1[628]; 
    assign out[146] = layer_1[729] | layer_1[605]; 
    assign out[147] = layer_1[1222] ^ layer_1[1273]; 
    assign out[148] = ~layer_1[1309] | (layer_1[1309] & layer_1[1429]); 
    assign out[149] = ~layer_1[1785] | (layer_1[1666] & layer_1[1785]); 
    assign out[150] = layer_1[2674] & ~layer_1[2565]; 
    assign out[151] = layer_1[2241]; 
    assign out[152] = ~layer_1[2500]; 
    assign out[153] = ~layer_1[2035]; 
    assign out[154] = ~layer_1[3201]; 
    assign out[155] = ~layer_1[544]; 
    assign out[156] = ~layer_1[56]; 
    assign out[157] = layer_1[3770] & ~layer_1[3817]; 
    assign out[158] = ~layer_1[2964]; 
    assign out[159] = ~(layer_1[3551] ^ layer_1[3476]); 
    assign out[160] = ~layer_1[1910]; 
    assign out[161] = layer_1[1798] ^ layer_1[1914]; 
    assign out[162] = layer_1[1059] & ~layer_1[979]; 
    assign out[163] = layer_1[1369] & ~layer_1[1417]; 
    assign out[164] = layer_1[3784] & layer_1[3775]; 
    assign out[165] = ~layer_1[3890]; 
    assign out[166] = layer_1[2883] & ~layer_1[2805]; 
    assign out[167] = layer_1[418]; 
    assign out[168] = ~layer_1[3957] | (layer_1[3957] & layer_1[3979]); 
    assign out[169] = ~layer_1[3631]; 
    assign out[170] = layer_1[3875] ^ layer_1[3976]; 
    assign out[171] = ~(layer_1[1180] ^ layer_1[1073]); 
    assign out[172] = layer_1[2191]; 
    assign out[173] = ~(layer_1[3558] & layer_1[3639]); 
    assign out[174] = ~(layer_1[749] | layer_1[764]); 
    assign out[175] = ~(layer_1[1267] & layer_1[1196]); 
    assign out[176] = ~(layer_1[1996] | layer_1[2066]); 
    assign out[177] = layer_1[2665]; 
    assign out[178] = ~(layer_1[1244] ^ layer_1[1201]); 
    assign out[179] = layer_1[3900] & ~layer_1[3810]; 
    assign out[180] = layer_1[2662]; 
    assign out[181] = ~layer_1[3144] | (layer_1[3164] & layer_1[3144]); 
    assign out[182] = layer_1[116]; 
    assign out[183] = ~(layer_1[1274] | layer_1[1224]); 
    assign out[184] = ~layer_1[620]; 
    assign out[185] = layer_1[2405] | layer_1[2398]; 
    assign out[186] = layer_1[16] & layer_1[137]; 
    assign out[187] = ~layer_1[1928] | (layer_1[1832] & layer_1[1928]); 
    assign out[188] = ~(layer_1[2889] | layer_1[2805]); 
    assign out[189] = layer_1[333] ^ layer_1[285]; 
    assign out[190] = ~layer_1[3832]; 
    assign out[191] = layer_1[884] & ~layer_1[979]; 
    assign out[192] = layer_1[3236] & ~layer_1[3194]; 
    assign out[193] = layer_1[130] & ~layer_1[44]; 
    assign out[194] = layer_1[3938]; 
    assign out[195] = layer_1[2595] | layer_1[2467]; 
    assign out[196] = ~layer_1[3688]; 
    assign out[197] = ~layer_1[290]; 
    assign out[198] = ~layer_1[3111]; 
    assign out[199] = ~(layer_1[51] | layer_1[109]); 
    assign out[200] = layer_1[1980] & layer_1[1861]; 
    assign out[201] = layer_1[3868]; 
    assign out[202] = layer_1[2671]; 
    assign out[203] = ~layer_1[989]; 
    assign out[204] = ~layer_1[460]; 
    assign out[205] = ~(layer_1[2086] & layer_1[2193]); 
    assign out[206] = layer_1[2830]; 
    assign out[207] = ~(layer_1[2962] ^ layer_1[2957]); 
    assign out[208] = ~(layer_1[1364] ^ layer_1[1486]); 
    assign out[209] = layer_1[3305] ^ layer_1[3318]; 
    assign out[210] = ~layer_1[2747]; 
    assign out[211] = ~(layer_1[3709] ^ layer_1[3702]); 
    assign out[212] = ~layer_1[3719]; 
    assign out[213] = ~(layer_1[2367] ^ layer_1[2306]); 
    assign out[214] = layer_1[1643] & ~layer_1[1609]; 
    assign out[215] = layer_1[2011] & ~layer_1[1993]; 
    assign out[216] = layer_1[2289] & layer_1[2324]; 
    assign out[217] = layer_1[3826] & layer_1[3868]; 
    assign out[218] = layer_1[1586]; 
    assign out[219] = layer_1[2578]; 
    assign out[220] = layer_1[3337]; 
    assign out[221] = layer_1[3218] ^ layer_1[3192]; 
    assign out[222] = ~(layer_1[1438] | layer_1[1483]); 
    assign out[223] = ~layer_1[1107]; 
    assign out[224] = ~(layer_1[1882] ^ layer_1[1949]); 
    assign out[225] = ~layer_1[1683]; 
    assign out[226] = ~(layer_1[1539] ^ layer_1[1472]); 
    assign out[227] = ~(layer_1[3425] | layer_1[3507]); 
    assign out[228] = ~(layer_1[923] ^ layer_1[1019]); 
    assign out[229] = layer_1[3769] ^ layer_1[3809]; 
    assign out[230] = ~(layer_1[2080] & layer_1[2108]); 
    assign out[231] = layer_1[1275] & ~layer_1[1157]; 
    assign out[232] = ~(layer_1[3721] ^ layer_1[3679]); 
    assign out[233] = ~layer_1[3905]; 
    assign out[234] = layer_1[3711] ^ layer_1[3747]; 
    assign out[235] = layer_1[489]; 
    assign out[236] = layer_1[945]; 
    assign out[237] = layer_1[2175]; 
    assign out[238] = ~layer_1[3403]; 
    assign out[239] = ~layer_1[3089]; 
    assign out[240] = ~layer_1[1150]; 
    assign out[241] = ~layer_1[2514]; 
    assign out[242] = layer_1[646]; 
    assign out[243] = layer_1[3265] & layer_1[3181]; 
    assign out[244] = ~layer_1[2942]; 
    assign out[245] = ~layer_1[2931]; 
    assign out[246] = ~(layer_1[915] ^ layer_1[868]); 
    assign out[247] = ~layer_1[2009]; 
    assign out[248] = layer_1[2372] & ~layer_1[2381]; 
    assign out[249] = layer_1[1112] ^ layer_1[1022]; 
    assign out[250] = ~layer_1[1985]; 
    assign out[251] = layer_1[3397] ^ layer_1[3517]; 
    assign out[252] = layer_1[687] ^ layer_1[751]; 
    assign out[253] = ~layer_1[499]; 
    assign out[254] = layer_1[2224] & ~layer_1[2168]; 
    assign out[255] = ~(layer_1[2503] ^ layer_1[2435]); 
    assign out[256] = layer_1[2734]; 
    assign out[257] = layer_1[601] & ~layer_1[586]; 
    assign out[258] = ~layer_1[663]; 
    assign out[259] = layer_1[510] & ~layer_1[613]; 
    assign out[260] = ~layer_1[3880] | (layer_1[3891] & layer_1[3880]); 
    assign out[261] = ~(layer_1[487] | layer_1[613]); 
    assign out[262] = layer_1[3974]; 
    assign out[263] = layer_1[1285] ^ layer_1[1187]; 
    assign out[264] = ~layer_1[1853] | (layer_1[1902] & layer_1[1853]); 
    assign out[265] = ~(layer_1[2059] ^ layer_1[2090]); 
    assign out[266] = layer_1[3964] & layer_1[3906]; 
    assign out[267] = ~layer_1[806]; 
    assign out[268] = layer_1[380] ^ layer_1[352]; 
    assign out[269] = ~(layer_1[1765] ^ layer_1[1845]); 
    assign out[270] = ~(layer_1[1157] | layer_1[1269]); 
    assign out[271] = layer_1[2395]; 
    assign out[272] = layer_1[289] ^ layer_1[249]; 
    assign out[273] = layer_1[368]; 
    assign out[274] = ~layer_1[1130]; 
    assign out[275] = layer_1[547]; 
    assign out[276] = layer_1[3184] & ~layer_1[3108]; 
    assign out[277] = ~layer_1[1250]; 
    assign out[278] = ~(layer_1[482] | layer_1[532]); 
    assign out[279] = ~(layer_1[1187] ^ layer_1[1217]); 
    assign out[280] = layer_1[3694] ^ layer_1[3795]; 
    assign out[281] = layer_1[321] ^ layer_1[430]; 
    assign out[282] = layer_1[174]; 
    assign out[283] = ~(layer_1[2244] ^ layer_1[2260]); 
    assign out[284] = layer_1[591] | layer_1[711]; 
    assign out[285] = ~layer_1[1731]; 
    assign out[286] = layer_1[2623]; 
    assign out[287] = layer_1[3610] ^ layer_1[3548]; 
    assign out[288] = ~layer_1[2931]; 
    assign out[289] = layer_1[1503] & layer_1[1449]; 
    assign out[290] = layer_1[721] & ~layer_1[839]; 
    assign out[291] = layer_1[442] & ~layer_1[388]; 
    assign out[292] = layer_1[2414]; 
    assign out[293] = layer_1[3298] ^ layer_1[3357]; 
    assign out[294] = layer_1[3048]; 
    assign out[295] = ~(layer_1[816] ^ layer_1[752]); 
    assign out[296] = ~(layer_1[1163] ^ layer_1[1206]); 
    assign out[297] = layer_1[646]; 
    assign out[298] = layer_1[420] ^ layer_1[425]; 
    assign out[299] = layer_1[1620]; 
    assign out[300] = layer_1[2670] & layer_1[2712]; 
    assign out[301] = layer_1[1445] & layer_1[1370]; 
    assign out[302] = layer_1[1988] | layer_1[1889]; 
    assign out[303] = layer_1[1645] ^ layer_1[1559]; 
    assign out[304] = layer_1[40] ^ layer_1[54]; 
    assign out[305] = layer_1[2536] & layer_1[2581]; 
    assign out[306] = layer_1[694]; 
    assign out[307] = layer_1[1887]; 
    assign out[308] = ~layer_1[3371]; 
    assign out[309] = ~layer_1[953] | (layer_1[964] & layer_1[953]); 
    assign out[310] = layer_1[3023] | layer_1[3081]; 
    assign out[311] = ~layer_1[772]; 
    assign out[312] = layer_1[1824] ^ layer_1[1851]; 
    assign out[313] = layer_1[288] ^ layer_1[192]; 
    assign out[314] = layer_1[3230]; 
    assign out[315] = layer_1[1325]; 
    assign out[316] = ~layer_1[1599]; 
    assign out[317] = layer_1[760] | layer_1[651]; 
    assign out[318] = ~(layer_1[1935] ^ layer_1[2028]); 
    assign out[319] = layer_1[2850] | layer_1[2733]; 
    assign out[320] = ~(layer_1[3554] ^ layer_1[3437]); 
    assign out[321] = layer_1[275] & ~layer_1[359]; 
    assign out[322] = layer_1[1449] & ~layer_1[1555]; 
    assign out[323] = ~layer_1[122]; 
    assign out[324] = layer_1[1698] ^ layer_1[1665]; 
    assign out[325] = layer_1[2788]; 
    assign out[326] = layer_1[1307] ^ layer_1[1403]; 
    assign out[327] = ~layer_1[861]; 
    assign out[328] = ~(layer_1[2805] | layer_1[2900]); 
    assign out[329] = layer_1[780]; 
    assign out[330] = layer_1[2372] ^ layer_1[2378]; 
    assign out[331] = ~layer_1[3890]; 
    assign out[332] = ~layer_1[2093]; 
    assign out[333] = layer_1[1913] & ~layer_1[1975]; 
    assign out[334] = ~layer_1[1428]; 
    assign out[335] = layer_1[733] ^ layer_1[840]; 
    assign out[336] = ~(layer_1[787] ^ layer_1[679]); 
    assign out[337] = layer_1[1704] ^ layer_1[1753]; 
    assign out[338] = ~layer_1[279]; 
    assign out[339] = ~layer_1[1615]; 
    assign out[340] = layer_1[1897]; 
    assign out[341] = ~(layer_1[253] ^ layer_1[354]); 
    assign out[342] = layer_1[3720]; 
    assign out[343] = layer_1[3088]; 
    assign out[344] = layer_1[3492]; 
    assign out[345] = layer_1[3918] & layer_1[3866]; 
    assign out[346] = layer_1[3889] & ~layer_1[3802]; 
    assign out[347] = ~layer_1[3309]; 
    assign out[348] = layer_1[3238]; 
    assign out[349] = layer_1[3642] & layer_1[3527]; 
    assign out[350] = layer_1[149]; 
    assign out[351] = layer_1[1586]; 
    assign out[352] = layer_1[2274] | layer_1[2164]; 
    assign out[353] = layer_1[3190] & ~layer_1[3142]; 
    assign out[354] = layer_1[3090]; 
    assign out[355] = layer_1[13] & ~layer_1[125]; 
    assign out[356] = ~layer_1[763] | (layer_1[675] & layer_1[763]); 
    assign out[357] = layer_1[652]; 
    assign out[358] = ~(layer_1[2124] ^ layer_1[2059]); 
    assign out[359] = ~(layer_1[747] ^ layer_1[719]); 
    assign out[360] = layer_1[3530] & layer_1[3444]; 
    assign out[361] = ~layer_1[1278] | (layer_1[1278] & layer_1[1349]); 
    assign out[362] = layer_1[870]; 
    assign out[363] = layer_1[3832] ^ layer_1[3947]; 
    assign out[364] = layer_1[3643]; 
    assign out[365] = layer_1[1990] & layer_1[2016]; 
    assign out[366] = ~layer_1[3188]; 
    assign out[367] = layer_1[1470] & layer_1[1495]; 
    assign out[368] = ~(layer_1[365] & layer_1[346]); 
    assign out[369] = ~(layer_1[3798] | layer_1[3882]); 
    assign out[370] = layer_1[640]; 
    assign out[371] = layer_1[3342] ^ layer_1[3272]; 
    assign out[372] = ~(layer_1[3737] ^ layer_1[3656]); 
    assign out[373] = ~(layer_1[3011] & layer_1[3050]); 
    assign out[374] = ~layer_1[882] | (layer_1[882] & layer_1[888]); 
    assign out[375] = ~(layer_1[2273] | layer_1[2211]); 
    assign out[376] = layer_1[170] & ~layer_1[44]; 
    assign out[377] = ~layer_1[1078]; 
    assign out[378] = layer_1[2222] ^ layer_1[2258]; 
    assign out[379] = ~(layer_1[3594] & layer_1[3638]); 
    assign out[380] = ~(layer_1[2447] ^ layer_1[2500]); 
    assign out[381] = ~layer_1[3365]; 
    assign out[382] = layer_1[3620]; 
    assign out[383] = ~layer_1[3839] | (layer_1[3934] & layer_1[3839]); 
    assign out[384] = ~(layer_1[3810] | layer_1[3688]); 
    assign out[385] = ~layer_1[850] | (layer_1[850] & layer_1[910]); 
    assign out[386] = layer_1[3348] & layer_1[3351]; 
    assign out[387] = layer_1[1829]; 
    assign out[388] = layer_1[2552]; 
    assign out[389] = layer_1[2100]; 
    assign out[390] = layer_1[2670]; 
    assign out[391] = ~layer_1[2647]; 
    assign out[392] = layer_1[2106] & layer_1[2122]; 
    assign out[393] = ~(layer_1[1145] ^ layer_1[1200]); 
    assign out[394] = layer_1[3598] & ~layer_1[3725]; 
    assign out[395] = layer_1[973]; 
    assign out[396] = layer_1[938] ^ layer_1[923]; 
    assign out[397] = layer_1[2620] & layer_1[2526]; 
    assign out[398] = layer_1[869] & ~layer_1[867]; 
    assign out[399] = ~(layer_1[2437] ^ layer_1[2483]); 
    assign out[400] = layer_1[2563] ^ layer_1[2649]; 
    assign out[401] = layer_1[2575]; 
    assign out[402] = layer_1[5] & ~layer_1[11]; 
    assign out[403] = ~layer_1[1941]; 
    assign out[404] = ~layer_1[3517]; 
    assign out[405] = layer_1[2999]; 
    assign out[406] = layer_1[3843] & layer_1[3966]; 
    assign out[407] = layer_1[2991] ^ layer_1[2922]; 
    assign out[408] = layer_1[2375] & ~layer_1[2466]; 
    assign out[409] = layer_1[2063] ^ layer_1[2186]; 
    assign out[410] = ~layer_1[493] | (layer_1[493] & layer_1[411]); 
    assign out[411] = ~(layer_1[318] ^ layer_1[234]); 
    assign out[412] = layer_1[2756] & ~layer_1[2864]; 
    assign out[413] = ~(layer_1[3163] ^ layer_1[3244]); 
    assign out[414] = ~(layer_1[510] | layer_1[387]); 
    assign out[415] = ~(layer_1[3438] ^ layer_1[3495]); 
    assign out[416] = ~layer_1[735]; 
    assign out[417] = layer_1[2017] & ~layer_1[1970]; 
    assign out[418] = ~layer_1[2520]; 
    assign out[419] = layer_1[1198]; 
    assign out[420] = layer_1[3019] & ~layer_1[3089]; 
    assign out[421] = layer_1[3384]; 
    assign out[422] = ~(layer_1[2620] ^ layer_1[2717]); 
    assign out[423] = ~layer_1[516] | (layer_1[518] & layer_1[516]); 
    assign out[424] = layer_1[2218] & layer_1[2093]; 
    assign out[425] = layer_1[965] ^ layer_1[837]; 
    assign out[426] = ~layer_1[929]; 
    assign out[427] = layer_1[819]; 
    assign out[428] = ~layer_1[2071]; 
    assign out[429] = ~layer_1[542]; 
    assign out[430] = ~layer_1[710]; 
    assign out[431] = ~(layer_1[1730] | layer_1[1694]); 
    assign out[432] = layer_1[2537] & ~layer_1[2418]; 
    assign out[433] = ~layer_1[2332] | (layer_1[2204] & layer_1[2332]); 
    assign out[434] = ~layer_1[3500] | (layer_1[3440] & layer_1[3500]); 
    assign out[435] = ~(layer_1[2828] & layer_1[2875]); 
    assign out[436] = ~layer_1[1912] | (layer_1[1846] & layer_1[1912]); 
    assign out[437] = layer_1[3142] & layer_1[3061]; 
    assign out[438] = ~(layer_1[2066] | layer_1[2056]); 
    assign out[439] = ~layer_1[2316]; 
    assign out[440] = ~layer_1[2473]; 
    assign out[441] = layer_1[2929] & ~layer_1[2947]; 
    assign out[442] = layer_1[36] & ~layer_1[49]; 
    assign out[443] = layer_1[3678] ^ layer_1[3651]; 
    assign out[444] = layer_1[1846] & layer_1[1956]; 
    assign out[445] = layer_1[1304] & ~layer_1[1344]; 
    assign out[446] = layer_1[3444] & ~layer_1[3494]; 
    assign out[447] = layer_1[3293] ^ layer_1[3255]; 
    assign out[448] = ~(layer_1[691] ^ layer_1[784]); 
    assign out[449] = layer_1[3719] & ~layer_1[3734]; 
    assign out[450] = layer_1[2204]; 
    assign out[451] = ~(layer_1[935] | layer_1[893]); 
    assign out[452] = ~layer_1[1006]; 
    assign out[453] = layer_1[1573]; 
    assign out[454] = ~layer_1[3475] | (layer_1[3475] & layer_1[3474]); 
    assign out[455] = layer_1[3927] & layer_1[3990]; 
    assign out[456] = layer_1[3848]; 
    assign out[457] = layer_1[2516] & ~layer_1[2546]; 
    assign out[458] = layer_1[272]; 
    assign out[459] = layer_1[815]; 
    assign out[460] = ~(layer_1[1716] ^ layer_1[1656]); 
    assign out[461] = layer_1[501]; 
    assign out[462] = layer_1[1525] & ~layer_1[1476]; 
    assign out[463] = ~(layer_1[1982] & layer_1[1941]); 
    assign out[464] = layer_1[500]; 
    assign out[465] = ~(layer_1[564] & layer_1[665]); 
    assign out[466] = ~(layer_1[3031] | layer_1[3040]); 
    assign out[467] = layer_1[1263] ^ layer_1[1140]; 
    assign out[468] = layer_1[3753] & ~layer_1[3801]; 
    assign out[469] = ~(layer_1[667] ^ layer_1[688]); 
    assign out[470] = layer_1[159] & ~layer_1[263]; 
    assign out[471] = ~layer_1[246]; 
    assign out[472] = ~(layer_1[1801] ^ layer_1[1928]); 
    assign out[473] = ~(layer_1[1299] | layer_1[1425]); 
    assign out[474] = layer_1[3019]; 
    assign out[475] = ~layer_1[3957]; 
    assign out[476] = layer_1[1629] & ~layer_1[1570]; 
    assign out[477] = ~(layer_1[3790] | layer_1[3794]); 
    assign out[478] = ~(layer_1[1310] ^ layer_1[1419]); 
    assign out[479] = layer_1[3559] & ~layer_1[3586]; 
    assign out[480] = ~layer_1[2832]; 
    assign out[481] = ~(layer_1[1081] | layer_1[974]); 
    assign out[482] = ~layer_1[1636] | (layer_1[1636] & layer_1[1621]); 
    assign out[483] = layer_1[822] & ~layer_1[915]; 
    assign out[484] = layer_1[1480]; 
    assign out[485] = layer_1[3986]; 
    assign out[486] = layer_1[1828]; 
    assign out[487] = ~(layer_1[2565] ^ layer_1[2562]); 
    assign out[488] = layer_1[3912] & layer_1[3929]; 
    assign out[489] = layer_1[3253] & ~layer_1[3245]; 
    assign out[490] = layer_1[818] ^ layer_1[752]; 
    assign out[491] = layer_1[304] ^ layer_1[323]; 
    assign out[492] = ~layer_1[97] | (layer_1[97] & layer_1[175]); 
    assign out[493] = ~layer_1[3453]; 
    assign out[494] = layer_1[3085] & ~layer_1[2973]; 
    assign out[495] = ~(layer_1[611] ^ layer_1[572]); 
    assign out[496] = layer_1[3807]; 
    assign out[497] = ~(layer_1[844] | layer_1[935]); 
    assign out[498] = layer_1[306] ^ layer_1[299]; 
    assign out[499] = ~layer_1[2702]; 
    assign out[500] = layer_1[3864] & ~layer_1[3974]; 
    assign out[501] = layer_1[3629] & ~layer_1[3744]; 
    assign out[502] = layer_1[1723] & layer_1[1827]; 
    assign out[503] = layer_1[1214] ^ layer_1[1207]; 
    assign out[504] = layer_1[3704] & ~layer_1[3663]; 
    assign out[505] = layer_1[1808] & ~layer_1[1707]; 
    assign out[506] = layer_1[31] & ~layer_1[33]; 
    assign out[507] = ~(layer_1[2902] ^ layer_1[2781]); 
    assign out[508] = ~layer_1[3653]; 
    assign out[509] = layer_1[1484] ^ layer_1[1410]; 
    assign out[510] = ~(layer_1[3960] | layer_1[3988]); 
    assign out[511] = layer_1[210] ^ layer_1[201]; 
    assign out[512] = ~layer_1[2413]; 
    assign out[513] = ~(layer_1[2053] | layer_1[1945]); 
    assign out[514] = ~(layer_1[138] ^ layer_1[161]); 
    assign out[515] = layer_1[2710] & layer_1[2636]; 
    assign out[516] = layer_1[946]; 
    assign out[517] = ~layer_1[3202]; 
    assign out[518] = ~layer_1[1336]; 
    assign out[519] = layer_1[1956]; 
    assign out[520] = layer_1[864] | layer_1[771]; 
    assign out[521] = layer_1[2787]; 
    assign out[522] = layer_1[3595] & layer_1[3572]; 
    assign out[523] = ~layer_1[3328] | (layer_1[3328] & layer_1[3216]); 
    assign out[524] = ~(layer_1[493] & layer_1[525]); 
    assign out[525] = ~(layer_1[657] | layer_1[710]); 
    assign out[526] = ~(layer_1[1775] | layer_1[1803]); 
    assign out[527] = ~layer_1[1290] | (layer_1[1290] & layer_1[1228]); 
    assign out[528] = ~(layer_1[2519] ^ layer_1[2451]); 
    assign out[529] = layer_1[3295]; 
    assign out[530] = layer_1[716] ^ layer_1[687]; 
    assign out[531] = layer_1[3160] ^ layer_1[3211]; 
    assign out[532] = layer_1[2429] & layer_1[2356]; 
    assign out[533] = layer_1[2085]; 
    assign out[534] = layer_1[2975] & layer_1[2950]; 
    assign out[535] = layer_1[3705]; 
    assign out[536] = ~(layer_1[2732] | layer_1[2608]); 
    assign out[537] = layer_1[423] & ~layer_1[315]; 
    assign out[538] = ~(layer_1[2421] ^ layer_1[2430]); 
    assign out[539] = layer_1[1864]; 
    assign out[540] = layer_1[1206] & ~layer_1[1171]; 
    assign out[541] = ~(layer_1[1508] & layer_1[1452]); 
    assign out[542] = layer_1[2375] & ~layer_1[2452]; 
    assign out[543] = layer_1[1607] | layer_1[1728]; 
    assign out[544] = layer_1[1230]; 
    assign out[545] = layer_1[345]; 
    assign out[546] = layer_1[2921] & ~layer_1[2942]; 
    assign out[547] = layer_1[2591] & layer_1[2676]; 
    assign out[548] = ~layer_1[2488]; 
    assign out[549] = layer_1[2247] & ~layer_1[2283]; 
    assign out[550] = ~layer_1[2167]; 
    assign out[551] = layer_1[2568]; 
    assign out[552] = ~(layer_1[3349] ^ layer_1[3235]); 
    assign out[553] = layer_1[1917] & ~layer_1[1810]; 
    assign out[554] = ~(layer_1[3369] | layer_1[3399]); 
    assign out[555] = ~layer_1[3781] | (layer_1[3696] & layer_1[3781]); 
    assign out[556] = layer_1[2951] ^ layer_1[2957]; 
    assign out[557] = layer_1[2872] & ~layer_1[2993]; 
    assign out[558] = ~layer_1[1381]; 
    assign out[559] = layer_1[297] & ~layer_1[361]; 
    assign out[560] = ~(layer_1[1579] | layer_1[1561]); 
    assign out[561] = ~layer_1[791] | (layer_1[791] & layer_1[763]); 
    assign out[562] = layer_1[151] & layer_1[55]; 
    assign out[563] = ~(layer_1[2599] ^ layer_1[2474]); 
    assign out[564] = layer_1[1174] & ~layer_1[1244]; 
    assign out[565] = ~(layer_1[126] ^ layer_1[54]); 
    assign out[566] = layer_1[268]; 
    assign out[567] = layer_1[1872] & ~layer_1[1916]; 
    assign out[568] = ~(layer_1[2367] ^ layer_1[2447]); 
    assign out[569] = layer_1[3625] & ~layer_1[3499]; 
    assign out[570] = layer_1[133] & layer_1[105]; 
    assign out[571] = layer_1[3106] & layer_1[3124]; 
    assign out[572] = ~(layer_1[3206] ^ layer_1[3099]); 
    assign out[573] = ~(layer_1[3095] | layer_1[3088]); 
    assign out[574] = layer_1[1814] & layer_1[1784]; 
    assign out[575] = layer_1[1671] & ~layer_1[1698]; 
    assign out[576] = layer_1[3805] & ~layer_1[3801]; 
    assign out[577] = ~layer_1[1697] | (layer_1[1683] & layer_1[1697]); 
    assign out[578] = layer_1[2789]; 
    assign out[579] = layer_1[1934] & ~layer_1[1947]; 
    assign out[580] = layer_1[1308] & ~layer_1[1226]; 
    assign out[581] = ~(layer_1[3560] ^ layer_1[3670]); 
    assign out[582] = layer_1[3216]; 
    assign out[583] = ~(layer_1[1408] | layer_1[1507]); 
    assign out[584] = layer_1[3733] & layer_1[3777]; 
    assign out[585] = layer_1[1062] ^ layer_1[989]; 
    assign out[586] = layer_1[2694] & ~layer_1[2708]; 
    assign out[587] = ~layer_1[3663]; 
    assign out[588] = ~(layer_1[1162] ^ layer_1[1168]); 
    assign out[589] = layer_1[2039] & ~layer_1[1970]; 
    assign out[590] = layer_1[3876]; 
    assign out[591] = layer_1[1143] & layer_1[1246]; 
    assign out[592] = ~layer_1[1725]; 
    assign out[593] = layer_1[1142] & layer_1[1105]; 
    assign out[594] = layer_1[970]; 
    assign out[595] = ~layer_1[3138]; 
    assign out[596] = layer_1[473] & ~layer_1[349]; 
    assign out[597] = layer_1[2375] & ~layer_1[2502]; 
    assign out[598] = ~(layer_1[2825] ^ layer_1[2859]); 
    assign out[599] = ~layer_1[3075]; 
    assign out[600] = ~layer_1[2742]; 
    assign out[601] = layer_1[2690] & layer_1[2601]; 
    assign out[602] = ~(layer_1[431] ^ layer_1[429]); 
    assign out[603] = layer_1[3717] & ~layer_1[3707]; 
    assign out[604] = layer_1[120] & ~layer_1[40]; 
    assign out[605] = layer_1[1759]; 
    assign out[606] = layer_1[825]; 
    assign out[607] = ~(layer_1[3615] ^ layer_1[3699]); 
    assign out[608] = layer_1[2879] & ~layer_1[2797]; 
    assign out[609] = layer_1[294] ^ layer_1[170]; 
    assign out[610] = ~(layer_1[1325] | layer_1[1229]); 
    assign out[611] = layer_1[2406]; 
    assign out[612] = ~layer_1[2604]; 
    assign out[613] = ~layer_1[2157]; 
    assign out[614] = layer_1[3321] & layer_1[3358]; 
    assign out[615] = layer_1[3345]; 
    assign out[616] = layer_1[386] & ~layer_1[480]; 
    assign out[617] = ~(layer_1[479] ^ layer_1[474]); 
    assign out[618] = ~layer_1[575]; 
    assign out[619] = ~layer_1[898]; 
    assign out[620] = layer_1[2204] & ~layer_1[2159]; 
    assign out[621] = layer_1[3382] & layer_1[3354]; 
    assign out[622] = layer_1[2495] & layer_1[2577]; 
    assign out[623] = layer_1[1214] ^ layer_1[1205]; 
    assign out[624] = layer_1[3538] & ~layer_1[3558]; 
    assign out[625] = ~layer_1[2157]; 
    assign out[626] = ~layer_1[3506]; 
    assign out[627] = layer_1[2961]; 
    assign out[628] = layer_1[3393] & ~layer_1[3330]; 
    assign out[629] = ~(layer_1[3406] ^ layer_1[3325]); 
    assign out[630] = layer_1[1640] ^ layer_1[1522]; 
    assign out[631] = ~(layer_1[3532] | layer_1[3413]); 
    assign out[632] = layer_1[2028] & ~layer_1[1909]; 
    assign out[633] = layer_1[509] ^ layer_1[440]; 
    assign out[634] = layer_1[2431] & ~layer_1[2370]; 
    assign out[635] = layer_1[423] & ~layer_1[436]; 
    assign out[636] = layer_1[1412] & layer_1[1456]; 
    assign out[637] = layer_1[3644] ^ layer_1[3516]; 
    assign out[638] = layer_1[3226] & ~layer_1[3309]; 
    assign out[639] = layer_1[533] & ~layer_1[572]; 
    assign out[640] = layer_1[3184] & layer_1[3137]; 
    assign out[641] = ~(layer_1[2951] | layer_1[2838]); 
    assign out[642] = layer_1[2193] & ~layer_1[2183]; 
    assign out[643] = layer_1[2171]; 
    assign out[644] = layer_1[771]; 
    assign out[645] = layer_1[840] & layer_1[871]; 
    assign out[646] = ~layer_1[691]; 
    assign out[647] = ~layer_1[1388]; 
    assign out[648] = layer_1[946]; 
    assign out[649] = layer_1[2672] & layer_1[2661]; 
    assign out[650] = ~(layer_1[2547] ^ layer_1[2528]); 
    assign out[651] = layer_1[2684] & ~layer_1[2797]; 
    assign out[652] = ~layer_1[3751]; 
    assign out[653] = ~layer_1[1893]; 
    assign out[654] = ~(layer_1[2075] ^ layer_1[2137]); 
    assign out[655] = layer_1[1093]; 
    assign out[656] = layer_1[2410] ^ layer_1[2431]; 
    assign out[657] = layer_1[2719] ^ layer_1[2714]; 
    assign out[658] = layer_1[459] & ~layer_1[536]; 
    assign out[659] = layer_1[409] & ~layer_1[435]; 
    assign out[660] = layer_1[1924] & layer_1[1865]; 
    assign out[661] = layer_1[3434] ^ layer_1[3325]; 
    assign out[662] = layer_1[1106] & ~layer_1[1057]; 
    assign out[663] = ~layer_1[1434]; 
    assign out[664] = layer_1[2485]; 
    assign out[665] = ~layer_1[3822]; 
    assign out[666] = layer_1[2665] ^ layer_1[2596]; 
    assign out[667] = layer_1[3789] & ~layer_1[3770]; 
    assign out[668] = ~(layer_1[528] | layer_1[599]); 
    assign out[669] = layer_1[286] & ~layer_1[376]; 
    assign out[670] = ~(layer_1[2751] | layer_1[2714]); 
    assign out[671] = ~layer_1[1869]; 
    assign out[672] = layer_1[2958]; 
    assign out[673] = ~(layer_1[531] | layer_1[651]); 
    assign out[674] = layer_1[3581]; 
    assign out[675] = layer_1[2907] & layer_1[2794]; 
    assign out[676] = layer_1[3027] & layer_1[2980]; 
    assign out[677] = ~layer_1[1989] | (layer_1[2016] & layer_1[1989]); 
    assign out[678] = layer_1[1889] & layer_1[1904]; 
    assign out[679] = layer_1[655] & layer_1[534]; 
    assign out[680] = layer_1[1142] & layer_1[1026]; 
    assign out[681] = layer_1[1083] & ~layer_1[1043]; 
    assign out[682] = layer_1[90] & ~layer_1[181]; 
    assign out[683] = layer_1[120] & ~layer_1[123]; 
    assign out[684] = layer_1[444]; 
    assign out[685] = layer_1[2399] & layer_1[2273]; 
    assign out[686] = layer_1[3273] & layer_1[3393]; 
    assign out[687] = ~(layer_1[924] ^ layer_1[900]); 
    assign out[688] = ~layer_1[700] | (layer_1[700] & layer_1[603]); 
    assign out[689] = ~(layer_1[448] ^ layer_1[568]); 
    assign out[690] = ~(layer_1[306] | layer_1[180]); 
    assign out[691] = layer_1[2899]; 
    assign out[692] = layer_1[193] ^ layer_1[203]; 
    assign out[693] = layer_1[2321]; 
    assign out[694] = layer_1[2684] & ~layer_1[2665]; 
    assign out[695] = layer_1[3009] & ~layer_1[3084]; 
    assign out[696] = layer_1[3653] ^ layer_1[3756]; 
    assign out[697] = layer_1[3862] & layer_1[3930]; 
    assign out[698] = layer_1[1094]; 
    assign out[699] = layer_1[96]; 
    assign out[700] = ~(layer_1[975] ^ layer_1[850]); 
    assign out[701] = ~(layer_1[1163] | layer_1[1085]); 
    assign out[702] = layer_1[1988]; 
    assign out[703] = layer_1[2061] | layer_1[2102]; 
    assign out[704] = ~layer_1[3032]; 
    assign out[705] = layer_1[1266] & layer_1[1220]; 
    assign out[706] = ~(layer_1[3219] ^ layer_1[3286]); 
    assign out[707] = layer_1[2709] ^ layer_1[2630]; 
    assign out[708] = ~(layer_1[3395] ^ layer_1[3425]); 
    assign out[709] = layer_1[744] & layer_1[711]; 
    assign out[710] = ~(layer_1[582] ^ layer_1[553]); 
    assign out[711] = layer_1[3223] ^ layer_1[3329]; 
    assign out[712] = layer_1[1119] & ~layer_1[1241]; 
    assign out[713] = ~(layer_1[625] ^ layer_1[539]); 
    assign out[714] = layer_1[1839]; 
    assign out[715] = ~layer_1[319]; 
    assign out[716] = layer_1[2160] & ~layer_1[2098]; 
    assign out[717] = layer_1[2781] ^ layer_1[2771]; 
    assign out[718] = layer_1[2258] & layer_1[2385]; 
    assign out[719] = layer_1[2222] & ~layer_1[2275]; 
    assign out[720] = ~(layer_1[3371] & layer_1[3372]); 
    assign out[721] = ~layer_1[3390]; 
    assign out[722] = ~(layer_1[3029] ^ layer_1[2970]); 
    assign out[723] = layer_1[3656] & ~layer_1[3724]; 
    assign out[724] = ~(layer_1[1111] | layer_1[1158]); 
    assign out[725] = ~layer_1[2917] | (layer_1[2917] & layer_1[2896]); 
    assign out[726] = ~layer_1[812]; 
    assign out[727] = layer_1[1776] & layer_1[1857]; 
    assign out[728] = ~layer_1[3514]; 
    assign out[729] = ~(layer_1[2340] ^ layer_1[2278]); 
    assign out[730] = layer_1[3562] ^ layer_1[3442]; 
    assign out[731] = layer_1[174]; 
    assign out[732] = layer_1[1917] & ~layer_1[1927]; 
    assign out[733] = layer_1[1225]; 
    assign out[734] = ~layer_1[1608] | (layer_1[1608] & layer_1[1543]); 
    assign out[735] = ~layer_1[830]; 
    assign out[736] = layer_1[3139] & layer_1[3197]; 
    assign out[737] = layer_1[1785]; 
    assign out[738] = ~layer_1[2031]; 
    assign out[739] = layer_1[3216] & ~layer_1[3100]; 
    assign out[740] = layer_1[24] ^ layer_1[70]; 
    assign out[741] = layer_1[597]; 
    assign out[742] = ~(layer_1[3048] ^ layer_1[3030]); 
    assign out[743] = ~(layer_1[225] | layer_1[132]); 
    assign out[744] = layer_1[3856] & layer_1[3953]; 
    assign out[745] = layer_1[119] | layer_1[90]; 
    assign out[746] = layer_1[2759] ^ layer_1[2792]; 
    assign out[747] = ~(layer_1[1567] | layer_1[1641]); 
    assign out[748] = ~(layer_1[2336] & layer_1[2434]); 
    assign out[749] = layer_1[3187] & layer_1[3174]; 
    assign out[750] = ~layer_1[77]; 
    assign out[751] = layer_1[290]; 
    assign out[752] = ~(layer_1[2276] | layer_1[2179]); 
    assign out[753] = ~layer_1[2768]; 
    assign out[754] = ~layer_1[1065] | (layer_1[1104] & layer_1[1065]); 
    assign out[755] = ~(layer_1[1488] & layer_1[1387]); 
    assign out[756] = ~layer_1[2357]; 
    assign out[757] = layer_1[3145] ^ layer_1[3209]; 
    assign out[758] = layer_1[144] ^ layer_1[111]; 
    assign out[759] = ~layer_1[1302]; 
    assign out[760] = layer_1[636]; 
    assign out[761] = layer_1[157] & ~layer_1[258]; 
    assign out[762] = layer_1[3135] ^ layer_1[3208]; 
    assign out[763] = layer_1[892]; 
    assign out[764] = layer_1[416] | layer_1[401]; 
    assign out[765] = layer_1[1658]; 
    assign out[766] = layer_1[3177] & layer_1[3155]; 
    assign out[767] = ~(layer_1[3961] | layer_1[3846]); 
    assign out[768] = ~(layer_1[736] | layer_1[701]); 
    assign out[769] = layer_1[2857]; 
    assign out[770] = layer_1[807]; 
    assign out[771] = ~layer_1[2417]; 
    assign out[772] = ~layer_1[915]; 
    assign out[773] = ~(layer_1[1081] & layer_1[1074]); 
    assign out[774] = ~(layer_1[3460] ^ layer_1[3587]); 
    assign out[775] = ~(layer_1[1528] & layer_1[1549]); 
    assign out[776] = layer_1[1505] & layer_1[1590]; 
    assign out[777] = ~(layer_1[2478] ^ layer_1[2490]); 
    assign out[778] = ~(layer_1[3743] ^ layer_1[3628]); 
    assign out[779] = layer_1[1980] ^ layer_1[1999]; 
    assign out[780] = ~(layer_1[1101] & layer_1[1080]); 
    assign out[781] = ~(layer_1[2466] | layer_1[2408]); 
    assign out[782] = ~layer_1[2955]; 
    assign out[783] = ~(layer_1[2973] | layer_1[3067]); 
    assign out[784] = layer_1[2647] & ~layer_1[2742]; 
    assign out[785] = ~layer_1[6]; 
    assign out[786] = ~(layer_1[733] ^ layer_1[613]); 
    assign out[787] = ~(layer_1[3066] ^ layer_1[3072]); 
    assign out[788] = ~layer_1[3156]; 
    assign out[789] = ~(layer_1[2630] ^ layer_1[2515]); 
    assign out[790] = ~layer_1[1465]; 
    assign out[791] = ~(layer_1[1346] | layer_1[1258]); 
    assign out[792] = ~layer_1[736] | (layer_1[729] & layer_1[736]); 
    assign out[793] = ~(layer_1[952] & layer_1[1032]); 
    assign out[794] = layer_1[2625]; 
    assign out[795] = layer_1[3504] & layer_1[3526]; 
    assign out[796] = ~(layer_1[3937] ^ layer_1[3863]); 
    assign out[797] = ~(layer_1[2618] | layer_1[2707]); 
    assign out[798] = ~layer_1[2942]; 
    assign out[799] = ~layer_1[894]; 
    assign out[800] = layer_1[729] ^ layer_1[616]; 
    assign out[801] = layer_1[465] & ~layer_1[528]; 
    assign out[802] = layer_1[3633]; 
    assign out[803] = ~layer_1[3483]; 
    assign out[804] = layer_1[1036] & ~layer_1[978]; 
    assign out[805] = layer_1[1972]; 
    assign out[806] = ~layer_1[3058]; 
    assign out[807] = ~(layer_1[2420] ^ layer_1[2516]); 
    assign out[808] = layer_1[3030] | layer_1[2958]; 
    assign out[809] = layer_1[2313]; 
    assign out[810] = layer_1[3468] | layer_1[3459]; 
    assign out[811] = ~(layer_1[2839] ^ layer_1[2809]); 
    assign out[812] = layer_1[2884]; 
    assign out[813] = ~(layer_1[3150] & layer_1[3161]); 
    assign out[814] = layer_1[1996] ^ layer_1[2016]; 
    assign out[815] = layer_1[350] ^ layer_1[419]; 
    assign out[816] = ~(layer_1[2642] ^ layer_1[2730]); 
    assign out[817] = ~layer_1[3832] | (layer_1[3808] & layer_1[3832]); 
    assign out[818] = layer_1[1425] ^ layer_1[1398]; 
    assign out[819] = layer_1[3089] ^ layer_1[3150]; 
    assign out[820] = ~layer_1[3035]; 
    assign out[821] = layer_1[1247]; 
    assign out[822] = layer_1[2621] ^ layer_1[2588]; 
    assign out[823] = layer_1[2388]; 
    assign out[824] = ~(layer_1[2149] ^ layer_1[2072]); 
    assign out[825] = layer_1[948] & layer_1[1049]; 
    assign out[826] = ~layer_1[1559]; 
    assign out[827] = ~layer_1[2023]; 
    assign out[828] = ~layer_1[1291] | (layer_1[1392] & layer_1[1291]); 
    assign out[829] = ~layer_1[3448] | (layer_1[3565] & layer_1[3448]); 
    assign out[830] = ~(layer_1[2179] & layer_1[2182]); 
    assign out[831] = layer_1[253] | layer_1[142]; 
    assign out[832] = ~layer_1[2786]; 
    assign out[833] = ~(layer_1[3110] ^ layer_1[3037]); 
    assign out[834] = layer_1[1026] ^ layer_1[1120]; 
    assign out[835] = ~layer_1[2363] | (layer_1[2363] & layer_1[2455]); 
    assign out[836] = ~(layer_1[1727] | layer_1[1704]); 
    assign out[837] = layer_1[1366] & ~layer_1[1494]; 
    assign out[838] = layer_1[3736]; 
    assign out[839] = layer_1[2918] ^ layer_1[2938]; 
    assign out[840] = ~layer_1[1653]; 
    assign out[841] = ~layer_1[407]; 
    assign out[842] = ~(layer_1[1587] & layer_1[1532]); 
    assign out[843] = layer_1[2219]; 
    assign out[844] = ~(layer_1[2205] & layer_1[2160]); 
    assign out[845] = ~(layer_1[331] & layer_1[306]); 
    assign out[846] = layer_1[21]; 
    assign out[847] = ~layer_1[1872] | (layer_1[1872] & layer_1[1945]); 
    assign out[848] = layer_1[3755]; 
    assign out[849] = ~(layer_1[610] ^ layer_1[623]); 
    assign out[850] = ~layer_1[1219]; 
    assign out[851] = layer_1[1211]; 
    assign out[852] = ~layer_1[3259]; 
    assign out[853] = layer_1[2443] ^ layer_1[2395]; 
    assign out[854] = layer_1[345] & ~layer_1[250]; 
    assign out[855] = ~layer_1[1504]; 
    assign out[856] = ~(layer_1[1844] ^ layer_1[1879]); 
    assign out[857] = ~(layer_1[2039] & layer_1[2010]); 
    assign out[858] = ~layer_1[2331]; 
    assign out[859] = layer_1[3624]; 
    assign out[860] = ~(layer_1[2696] ^ layer_1[2590]); 
    assign out[861] = ~layer_1[3896] | (layer_1[3991] & layer_1[3896]); 
    assign out[862] = layer_1[1056] ^ layer_1[1053]; 
    assign out[863] = layer_1[2919]; 
    assign out[864] = ~layer_1[2912]; 
    assign out[865] = layer_1[1146] ^ layer_1[1168]; 
    assign out[866] = ~(layer_1[3723] & layer_1[3694]); 
    assign out[867] = layer_1[2457] & layer_1[2415]; 
    assign out[868] = layer_1[457] | layer_1[518]; 
    assign out[869] = layer_1[3720] & layer_1[3775]; 
    assign out[870] = ~layer_1[2422] | (layer_1[2422] & layer_1[2513]); 
    assign out[871] = ~(layer_1[284] & layer_1[375]); 
    assign out[872] = ~(layer_1[2080] ^ layer_1[1965]); 
    assign out[873] = ~layer_1[1011]; 
    assign out[874] = layer_1[2893]; 
    assign out[875] = ~layer_1[340]; 
    assign out[876] = layer_1[3591] ^ layer_1[3716]; 
    assign out[877] = ~layer_1[1830]; 
    assign out[878] = ~(layer_1[3779] | layer_1[3738]); 
    assign out[879] = ~layer_1[893]; 
    assign out[880] = layer_1[566] ^ layer_1[656]; 
    assign out[881] = ~(layer_1[2258] ^ layer_1[2166]); 
    assign out[882] = ~layer_1[1590] | (layer_1[1590] & layer_1[1513]); 
    assign out[883] = ~layer_1[3404] | (layer_1[3463] & layer_1[3404]); 
    assign out[884] = ~(layer_1[1688] ^ layer_1[1664]); 
    assign out[885] = ~(layer_1[1387] ^ layer_1[1499]); 
    assign out[886] = layer_1[1458] ^ layer_1[1556]; 
    assign out[887] = ~layer_1[926] | (layer_1[926] & layer_1[823]); 
    assign out[888] = layer_1[3571]; 
    assign out[889] = layer_1[194] ^ layer_1[134]; 
    assign out[890] = layer_1[244] & ~layer_1[132]; 
    assign out[891] = layer_1[1848] & ~layer_1[1750]; 
    assign out[892] = ~layer_1[1788]; 
    assign out[893] = ~(layer_1[100] ^ layer_1[69]); 
    assign out[894] = layer_1[3274]; 
    assign out[895] = layer_1[2944] & ~layer_1[2973]; 
    assign out[896] = ~(layer_1[3227] & layer_1[3254]); 
    assign out[897] = ~(layer_1[678] ^ layer_1[654]); 
    assign out[898] = ~(layer_1[922] ^ layer_1[955]); 
    assign out[899] = layer_1[3671]; 
    assign out[900] = ~layer_1[3042]; 
    assign out[901] = ~layer_1[1910] | (layer_1[1910] & layer_1[1817]); 
    assign out[902] = ~layer_1[3491]; 
    assign out[903] = layer_1[976]; 
    assign out[904] = ~layer_1[1673]; 
    assign out[905] = layer_1[491]; 
    assign out[906] = ~(layer_1[831] ^ layer_1[725]); 
    assign out[907] = ~layer_1[2023]; 
    assign out[908] = ~layer_1[2077]; 
    assign out[909] = ~(layer_1[2308] ^ layer_1[2250]); 
    assign out[910] = ~layer_1[3074]; 
    assign out[911] = layer_1[3852] ^ layer_1[3743]; 
    assign out[912] = ~layer_1[1213]; 
    assign out[913] = layer_1[890] ^ layer_1[813]; 
    assign out[914] = ~(layer_1[2934] ^ layer_1[2973]); 
    assign out[915] = layer_1[1145]; 
    assign out[916] = ~layer_1[1987]; 
    assign out[917] = layer_1[2986] ^ layer_1[3048]; 
    assign out[918] = layer_1[3470]; 
    assign out[919] = layer_1[2929]; 
    assign out[920] = layer_1[912]; 
    assign out[921] = layer_1[372] ^ layer_1[276]; 
    assign out[922] = ~layer_1[3091]; 
    assign out[923] = ~layer_1[3393]; 
    assign out[924] = layer_1[2538]; 
    assign out[925] = layer_1[3856] & ~layer_1[3848]; 
    assign out[926] = ~(layer_1[2706] ^ layer_1[2648]); 
    assign out[927] = ~layer_1[3632] | (layer_1[3632] & layer_1[3596]); 
    assign out[928] = ~layer_1[2067]; 
    assign out[929] = ~layer_1[1928] | (layer_1[1928] & layer_1[1919]); 
    assign out[930] = layer_1[458]; 
    assign out[931] = ~(layer_1[1071] ^ layer_1[1037]); 
    assign out[932] = ~layer_1[1689] | (layer_1[1814] & layer_1[1689]); 
    assign out[933] = ~layer_1[1065]; 
    assign out[934] = layer_1[1619]; 
    assign out[935] = ~layer_1[3483]; 
    assign out[936] = ~layer_1[2020] | (layer_1[2125] & layer_1[2020]); 
    assign out[937] = layer_1[256]; 
    assign out[938] = layer_1[1173] & layer_1[1216]; 
    assign out[939] = ~layer_1[431] | (layer_1[372] & layer_1[431]); 
    assign out[940] = layer_1[2383]; 
    assign out[941] = layer_1[3585] ^ layer_1[3461]; 
    assign out[942] = layer_1[3096]; 
    assign out[943] = ~layer_1[1524] | (layer_1[1524] & layer_1[1497]); 
    assign out[944] = ~layer_1[1622] | (layer_1[1622] & layer_1[1568]); 
    assign out[945] = layer_1[3871]; 
    assign out[946] = layer_1[2210] ^ layer_1[2204]; 
    assign out[947] = ~layer_1[610]; 
    assign out[948] = layer_1[2841] | layer_1[2862]; 
    assign out[949] = ~(layer_1[1592] ^ layer_1[1687]); 
    assign out[950] = ~layer_1[2599]; 
    assign out[951] = ~(layer_1[1490] & layer_1[1566]); 
    assign out[952] = layer_1[2643] ^ layer_1[2595]; 
    assign out[953] = ~layer_1[1516] | (layer_1[1593] & layer_1[1516]); 
    assign out[954] = ~(layer_1[2907] | layer_1[2899]); 
    assign out[955] = ~layer_1[2803] | (layer_1[2905] & layer_1[2803]); 
    assign out[956] = layer_1[30] & ~layer_1[98]; 
    assign out[957] = ~layer_1[1102]; 
    assign out[958] = layer_1[530] ^ layer_1[576]; 
    assign out[959] = layer_1[2294] & ~layer_1[2170]; 
    assign out[960] = layer_1[2903]; 
    assign out[961] = ~(layer_1[2963] ^ layer_1[2971]); 
    assign out[962] = layer_1[3096] ^ layer_1[3101]; 
    assign out[963] = layer_1[1581] | layer_1[1582]; 
    assign out[964] = ~(layer_1[2676] ^ layer_1[2675]); 
    assign out[965] = ~layer_1[1136]; 
    assign out[966] = layer_1[2388]; 
    assign out[967] = ~(layer_1[2550] ^ layer_1[2529]); 
    assign out[968] = ~layer_1[1675] | (layer_1[1675] & layer_1[1714]); 
    assign out[969] = ~(layer_1[196] ^ layer_1[221]); 
    assign out[970] = ~layer_1[705]; 
    assign out[971] = ~(layer_1[3445] ^ layer_1[3549]); 
    assign out[972] = ~(layer_1[3077] ^ layer_1[3032]); 
    assign out[973] = layer_1[2255] & ~layer_1[2176]; 
    assign out[974] = ~(layer_1[2591] ^ layer_1[2600]); 
    assign out[975] = layer_1[301] | layer_1[333]; 
    assign out[976] = ~(layer_1[193] & layer_1[194]); 
    assign out[977] = layer_1[2994]; 
    assign out[978] = layer_1[2064] & ~layer_1[2046]; 
    assign out[979] = ~layer_1[396]; 
    assign out[980] = ~layer_1[3349]; 
    assign out[981] = layer_1[2253] & layer_1[2152]; 
    assign out[982] = ~layer_1[3328] | (layer_1[3362] & layer_1[3328]); 
    assign out[983] = ~(layer_1[921] & layer_1[903]); 
    assign out[984] = ~layer_1[3474]; 
    assign out[985] = ~layer_1[2185] | (layer_1[2201] & layer_1[2185]); 
    assign out[986] = layer_1[1666] & ~layer_1[1663]; 
    assign out[987] = layer_1[2709] & ~layer_1[2625]; 
    assign out[988] = ~layer_1[289] | (layer_1[172] & layer_1[289]); 
    assign out[989] = layer_1[1182] & layer_1[1196]; 
    assign out[990] = ~(layer_1[2137] ^ layer_1[2114]); 
    assign out[991] = layer_1[965]; 
    assign out[992] = ~(layer_1[1103] ^ layer_1[1038]); 
    assign out[993] = layer_1[1463] & layer_1[1568]; 
    assign out[994] = layer_1[354] ^ layer_1[437]; 
    assign out[995] = ~(layer_1[1667] ^ layer_1[1664]); 
    assign out[996] = ~layer_1[566]; 
    assign out[997] = ~(layer_1[491] ^ layer_1[399]); 
    assign out[998] = layer_1[3885]; 
    assign out[999] = ~layer_1[763] | (layer_1[763] & layer_1[732]); 
    assign out[1000] = layer_1[3797]; 
    assign out[1001] = ~layer_1[1665]; 
    assign out[1002] = ~(layer_1[192] ^ layer_1[95]); 
    assign out[1003] = ~(layer_1[210] ^ layer_1[266]); 
    assign out[1004] = ~(layer_1[860] ^ layer_1[931]); 
    assign out[1005] = layer_1[1216] & ~layer_1[1254]; 
    assign out[1006] = ~layer_1[1727]; 
    assign out[1007] = ~layer_1[586]; 
    assign out[1008] = ~(layer_1[1888] ^ layer_1[1901]); 
    assign out[1009] = layer_1[2340] & ~layer_1[2298]; 
    assign out[1010] = ~layer_1[3374] | (layer_1[3399] & layer_1[3374]); 
    assign out[1011] = ~(layer_1[1694] ^ layer_1[1767]); 
    assign out[1012] = ~layer_1[455]; 
    assign out[1013] = layer_1[1313] ^ layer_1[1304]; 
    assign out[1014] = layer_1[2414] & ~layer_1[2325]; 
    assign out[1015] = ~(layer_1[1981] ^ layer_1[2106]); 
    assign out[1016] = ~(layer_1[3055] ^ layer_1[3129]); 
    assign out[1017] = layer_1[1911]; 
    assign out[1018] = layer_1[666]; 
    assign out[1019] = ~layer_1[3151]; 
    assign out[1020] = layer_1[247] & layer_1[261]; 
    assign out[1021] = ~(layer_1[2953] & layer_1[3041]); 
    assign out[1022] = layer_1[1176] ^ layer_1[1178]; 
    assign out[1023] = ~layer_1[1989]; 
    assign out[1024] = layer_1[3094] & ~layer_1[3182]; 
    assign out[1025] = ~layer_1[3303]; 
    assign out[1026] = ~(layer_1[3277] & layer_1[3178]); 
    assign out[1027] = ~layer_1[3388]; 
    assign out[1028] = layer_1[1539]; 
    assign out[1029] = layer_1[2844] & ~layer_1[2767]; 
    assign out[1030] = layer_1[3306] & ~layer_1[3260]; 
    assign out[1031] = ~layer_1[3575]; 
    assign out[1032] = layer_1[39]; 
    assign out[1033] = layer_1[996] & layer_1[985]; 
    assign out[1034] = layer_1[229]; 
    assign out[1035] = ~(layer_1[1242] ^ layer_1[1207]); 
    assign out[1036] = ~(layer_1[3265] & layer_1[3314]); 
    assign out[1037] = ~layer_1[2724] | (layer_1[2724] & layer_1[2632]); 
    assign out[1038] = layer_1[2177] & layer_1[2236]; 
    assign out[1039] = ~(layer_1[3167] ^ layer_1[3050]); 
    assign out[1040] = layer_1[314]; 
    assign out[1041] = layer_1[3698] ^ layer_1[3714]; 
    assign out[1042] = layer_1[1643] & ~layer_1[1644]; 
    assign out[1043] = layer_1[495]; 
    assign out[1044] = layer_1[2021] & layer_1[2040]; 
    assign out[1045] = ~layer_1[2323]; 
    assign out[1046] = layer_1[3786]; 
    assign out[1047] = ~layer_1[1768]; 
    assign out[1048] = layer_1[3959] & ~layer_1[3911]; 
    assign out[1049] = ~layer_1[813]; 
    assign out[1050] = layer_1[2988] ^ layer_1[3099]; 
    assign out[1051] = layer_1[1536]; 
    assign out[1052] = ~(layer_1[779] ^ layer_1[845]); 
    assign out[1053] = layer_1[3888] | layer_1[3790]; 
    assign out[1054] = layer_1[795] ^ layer_1[823]; 
    assign out[1055] = layer_1[630] & ~layer_1[599]; 
    assign out[1056] = ~(layer_1[516] ^ layer_1[623]); 
    assign out[1057] = layer_1[2877] & ~layer_1[2926]; 
    assign out[1058] = ~layer_1[1335]; 
    assign out[1059] = ~layer_1[171] | (layer_1[171] & layer_1[92]); 
    assign out[1060] = layer_1[1214] | layer_1[1268]; 
    assign out[1061] = layer_1[2749]; 
    assign out[1062] = ~(layer_1[1427] | layer_1[1406]); 
    assign out[1063] = layer_1[957]; 
    assign out[1064] = ~(layer_1[3582] & layer_1[3485]); 
    assign out[1065] = layer_1[3228] ^ layer_1[3184]; 
    assign out[1066] = ~layer_1[619]; 
    assign out[1067] = ~(layer_1[1160] ^ layer_1[1173]); 
    assign out[1068] = ~layer_1[1245] | (layer_1[1218] & layer_1[1245]); 
    assign out[1069] = layer_1[3368] ^ layer_1[3245]; 
    assign out[1070] = layer_1[985] ^ layer_1[859]; 
    assign out[1071] = ~(layer_1[2740] ^ layer_1[2687]); 
    assign out[1072] = layer_1[163] ^ layer_1[113]; 
    assign out[1073] = ~layer_1[3001] | (layer_1[3001] & layer_1[2939]); 
    assign out[1074] = ~layer_1[3970]; 
    assign out[1075] = layer_1[3006]; 
    assign out[1076] = layer_1[635] & layer_1[738]; 
    assign out[1077] = layer_1[1376] | layer_1[1258]; 
    assign out[1078] = layer_1[317]; 
    assign out[1079] = layer_1[2537] | layer_1[2605]; 
    assign out[1080] = ~layer_1[1086] | (layer_1[1086] & layer_1[1059]); 
    assign out[1081] = layer_1[3266] ^ layer_1[3306]; 
    assign out[1082] = ~(layer_1[3745] ^ layer_1[3654]); 
    assign out[1083] = layer_1[58] & layer_1[78]; 
    assign out[1084] = ~(layer_1[3151] | layer_1[3135]); 
    assign out[1085] = ~layer_1[2692] | (layer_1[2692] & layer_1[2791]); 
    assign out[1086] = ~layer_1[2196]; 
    assign out[1087] = ~layer_1[1922]; 
    assign out[1088] = layer_1[3742]; 
    assign out[1089] = layer_1[614]; 
    assign out[1090] = layer_1[1662] & ~layer_1[1541]; 
    assign out[1091] = layer_1[246] | layer_1[328]; 
    assign out[1092] = ~(layer_1[2189] | layer_1[2276]); 
    assign out[1093] = layer_1[1415] & layer_1[1496]; 
    assign out[1094] = ~(layer_1[3042] & layer_1[2953]); 
    assign out[1095] = ~(layer_1[3686] ^ layer_1[3724]); 
    assign out[1096] = ~layer_1[1347]; 
    assign out[1097] = ~layer_1[1131]; 
    assign out[1098] = layer_1[94]; 
    assign out[1099] = layer_1[2377] & ~layer_1[2298]; 
    assign out[1100] = layer_1[570] ^ layer_1[454]; 
    assign out[1101] = layer_1[911] & ~layer_1[783]; 
    assign out[1102] = layer_1[3400] ^ layer_1[3442]; 
    assign out[1103] = ~(layer_1[3187] & layer_1[3073]); 
    assign out[1104] = ~(layer_1[2466] & layer_1[2374]); 
    assign out[1105] = layer_1[1330] & ~layer_1[1287]; 
    assign out[1106] = ~(layer_1[2663] & layer_1[2581]); 
    assign out[1107] = layer_1[3786] & ~layer_1[3768]; 
    assign out[1108] = ~layer_1[3632]; 
    assign out[1109] = layer_1[2242]; 
    assign out[1110] = ~layer_1[3224]; 
    assign out[1111] = ~(layer_1[276] ^ layer_1[351]); 
    assign out[1112] = ~(layer_1[2878] | layer_1[2802]); 
    assign out[1113] = ~layer_1[794] | (layer_1[850] & layer_1[794]); 
    assign out[1114] = ~(layer_1[3430] | layer_1[3440]); 
    assign out[1115] = ~(layer_1[1401] | layer_1[1356]); 
    assign out[1116] = ~(layer_1[3417] ^ layer_1[3366]); 
    assign out[1117] = ~(layer_1[3812] ^ layer_1[3785]); 
    assign out[1118] = ~layer_1[2661] | (layer_1[2661] & layer_1[2544]); 
    assign out[1119] = ~layer_1[735]; 
    assign out[1120] = ~layer_1[3677]; 
    assign out[1121] = layer_1[235] & ~layer_1[167]; 
    assign out[1122] = layer_1[424] & ~layer_1[477]; 
    assign out[1123] = layer_1[1829]; 
    assign out[1124] = ~layer_1[863] | (layer_1[800] & layer_1[863]); 
    assign out[1125] = layer_1[1743] ^ layer_1[1756]; 
    assign out[1126] = ~(layer_1[3636] | layer_1[3668]); 
    assign out[1127] = layer_1[3840] | layer_1[3944]; 
    assign out[1128] = layer_1[2147] & ~layer_1[2256]; 
    assign out[1129] = layer_1[1376] | layer_1[1327]; 
    assign out[1130] = layer_1[1657] ^ layer_1[1766]; 
    assign out[1131] = ~layer_1[2400] | (layer_1[2400] & layer_1[2492]); 
    assign out[1132] = ~layer_1[1793] | (layer_1[1793] & layer_1[1811]); 
    assign out[1133] = ~layer_1[1980] | (layer_1[1980] & layer_1[2105]); 
    assign out[1134] = ~layer_1[3363]; 
    assign out[1135] = ~(layer_1[2460] & layer_1[2386]); 
    assign out[1136] = ~layer_1[2966] | (layer_1[2838] & layer_1[2966]); 
    assign out[1137] = ~(layer_1[1156] | layer_1[1234]); 
    assign out[1138] = layer_1[1577]; 
    assign out[1139] = layer_1[724]; 
    assign out[1140] = ~layer_1[826] | (layer_1[826] & layer_1[733]); 
    assign out[1141] = ~(layer_1[3525] ^ layer_1[3503]); 
    assign out[1142] = layer_1[894] & ~layer_1[1005]; 
    assign out[1143] = layer_1[2070] & ~layer_1[2107]; 
    assign out[1144] = ~layer_1[3733]; 
    assign out[1145] = ~layer_1[826]; 
    assign out[1146] = layer_1[2255] & layer_1[2367]; 
    assign out[1147] = layer_1[2018] | layer_1[1998]; 
    assign out[1148] = layer_1[3071]; 
    assign out[1149] = layer_1[717]; 
    assign out[1150] = ~(layer_1[273] ^ layer_1[268]); 
    assign out[1151] = layer_1[1389] ^ layer_1[1341]; 
    assign out[1152] = layer_1[3509]; 
    assign out[1153] = layer_1[3923] ^ layer_1[3838]; 
    assign out[1154] = ~layer_1[2746]; 
    assign out[1155] = ~layer_1[3131] | (layer_1[3131] & layer_1[3128]); 
    assign out[1156] = ~layer_1[3137]; 
    assign out[1157] = ~layer_1[2913]; 
    assign out[1158] = ~(layer_1[1136] & layer_1[1021]); 
    assign out[1159] = layer_1[3368] & ~layer_1[3296]; 
    assign out[1160] = ~(layer_1[607] ^ layer_1[568]); 
    assign out[1161] = ~layer_1[2683]; 
    assign out[1162] = ~layer_1[1267] | (layer_1[1267] & layer_1[1368]); 
    assign out[1163] = ~layer_1[3456]; 
    assign out[1164] = layer_1[2228]; 
    assign out[1165] = ~layer_1[277]; 
    assign out[1166] = ~layer_1[3813] | (layer_1[3836] & layer_1[3813]); 
    assign out[1167] = ~layer_1[1563] | (layer_1[1563] & layer_1[1530]); 
    assign out[1168] = layer_1[867] & ~layer_1[914]; 
    assign out[1169] = ~(layer_1[133] ^ layer_1[150]); 
    assign out[1170] = ~(layer_1[3551] ^ layer_1[3535]); 
    assign out[1171] = ~layer_1[567] | (layer_1[567] & layer_1[609]); 
    assign out[1172] = layer_1[1409] | layer_1[1462]; 
    assign out[1173] = ~layer_1[744] | (layer_1[744] & layer_1[724]); 
    assign out[1174] = ~layer_1[2443]; 
    assign out[1175] = layer_1[2439] & ~layer_1[2396]; 
    assign out[1176] = layer_1[1973]; 
    assign out[1177] = layer_1[866]; 
    assign out[1178] = ~(layer_1[2171] ^ layer_1[2159]); 
    assign out[1179] = ~(layer_1[490] & layer_1[411]); 
    assign out[1180] = ~(layer_1[143] ^ layer_1[113]); 
    assign out[1181] = layer_1[2305]; 
    assign out[1182] = layer_1[1493]; 
    assign out[1183] = layer_1[3281] & ~layer_1[3310]; 
    assign out[1184] = ~(layer_1[1498] ^ layer_1[1463]); 
    assign out[1185] = layer_1[2201] | layer_1[2293]; 
    assign out[1186] = layer_1[1116]; 
    assign out[1187] = ~(layer_1[2011] ^ layer_1[2000]); 
    assign out[1188] = ~layer_1[2843]; 
    assign out[1189] = layer_1[452] ^ layer_1[513]; 
    assign out[1190] = ~layer_1[3405] | (layer_1[3405] & layer_1[3397]); 
    assign out[1191] = ~(layer_1[507] ^ layer_1[531]); 
    assign out[1192] = layer_1[1002]; 
    assign out[1193] = layer_1[3986] | layer_1[3919]; 
    assign out[1194] = layer_1[3748] & layer_1[3753]; 
    assign out[1195] = ~layer_1[3156] | (layer_1[3036] & layer_1[3156]); 
    assign out[1196] = layer_1[2837] ^ layer_1[2738]; 
    assign out[1197] = ~(layer_1[1199] & layer_1[1168]); 
    assign out[1198] = ~layer_1[3409] | (layer_1[3409] & layer_1[3511]); 
    assign out[1199] = ~layer_1[3407]; 
    assign out[1200] = layer_1[3294]; 
    assign out[1201] = ~(layer_1[1092] | layer_1[1043]); 
    assign out[1202] = ~layer_1[3149] | (layer_1[3030] & layer_1[3149]); 
    assign out[1203] = ~(layer_1[2731] | layer_1[2621]); 
    assign out[1204] = layer_1[1086] & layer_1[1097]; 
    assign out[1205] = ~layer_1[3219] | (layer_1[3219] & layer_1[3249]); 
    assign out[1206] = ~layer_1[2407]; 
    assign out[1207] = ~layer_1[3589] | (layer_1[3651] & layer_1[3589]); 
    assign out[1208] = layer_1[400]; 
    assign out[1209] = ~layer_1[3427]; 
    assign out[1210] = layer_1[2267] | layer_1[2187]; 
    assign out[1211] = layer_1[2155]; 
    assign out[1212] = layer_1[2765]; 
    assign out[1213] = layer_1[2738] | layer_1[2760]; 
    assign out[1214] = layer_1[3803]; 
    assign out[1215] = ~(layer_1[1707] ^ layer_1[1689]); 
    assign out[1216] = layer_1[20] ^ layer_1[138]; 
    assign out[1217] = layer_1[72]; 
    assign out[1218] = ~layer_1[3368]; 
    assign out[1219] = ~layer_1[3407]; 
    assign out[1220] = ~(layer_1[2745] | layer_1[2647]); 
    assign out[1221] = ~layer_1[152] | (layer_1[99] & layer_1[152]); 
    assign out[1222] = layer_1[1205]; 
    assign out[1223] = layer_1[939] & ~layer_1[978]; 
    assign out[1224] = layer_1[787] ^ layer_1[707]; 
    assign out[1225] = layer_1[3015]; 
    assign out[1226] = ~layer_1[2117] | (layer_1[2117] & layer_1[2002]); 
    assign out[1227] = layer_1[3596]; 
    assign out[1228] = ~layer_1[767]; 
    assign out[1229] = ~layer_1[3041]; 
    assign out[1230] = layer_1[2136] & layer_1[2028]; 
    assign out[1231] = layer_1[2009] ^ layer_1[2089]; 
    assign out[1232] = ~(layer_1[1377] | layer_1[1474]); 
    assign out[1233] = ~(layer_1[3256] ^ layer_1[3178]); 
    assign out[1234] = layer_1[3825] & layer_1[3839]; 
    assign out[1235] = layer_1[301] ^ layer_1[377]; 
    assign out[1236] = layer_1[1871]; 
    assign out[1237] = ~layer_1[769] | (layer_1[769] & layer_1[812]); 
    assign out[1238] = ~(layer_1[3595] ^ layer_1[3476]); 
    assign out[1239] = layer_1[1541] & layer_1[1666]; 
    assign out[1240] = layer_1[1263]; 
    assign out[1241] = ~(layer_1[3705] & layer_1[3737]); 
    assign out[1242] = layer_1[3675]; 
    assign out[1243] = ~layer_1[603]; 
    assign out[1244] = ~(layer_1[2167] ^ layer_1[2108]); 
    assign out[1245] = ~layer_1[3846]; 
    assign out[1246] = layer_1[1419] ^ layer_1[1491]; 
    assign out[1247] = ~layer_1[935] | (layer_1[1057] & layer_1[935]); 
    assign out[1248] = ~layer_1[715] | (layer_1[613] & layer_1[715]); 
    assign out[1249] = layer_1[3341] & ~layer_1[3441]; 
    assign out[1250] = layer_1[1799]; 
    assign out[1251] = ~layer_1[1635]; 
    assign out[1252] = layer_1[210] & layer_1[260]; 
    assign out[1253] = ~(layer_1[2669] ^ layer_1[2761]); 
    assign out[1254] = ~(layer_1[3717] ^ layer_1[3660]); 
    assign out[1255] = layer_1[13]; 
    assign out[1256] = layer_1[2591]; 
    assign out[1257] = layer_1[1789] ^ layer_1[1770]; 
    assign out[1258] = layer_1[3672]; 
    assign out[1259] = ~layer_1[2140] | (layer_1[2140] & layer_1[2106]); 
    assign out[1260] = layer_1[1765]; 
    assign out[1261] = ~layer_1[825]; 
    assign out[1262] = ~layer_1[1239]; 
    assign out[1263] = layer_1[858] & ~layer_1[969]; 
    assign out[1264] = layer_1[3339] ^ layer_1[3221]; 
    assign out[1265] = ~(layer_1[3929] ^ layer_1[3816]); 
    assign out[1266] = layer_1[1566] ^ layer_1[1545]; 
    assign out[1267] = layer_1[1180] | layer_1[1296]; 
    assign out[1268] = ~(layer_1[3101] ^ layer_1[3135]); 
    assign out[1269] = layer_1[1434]; 
    assign out[1270] = layer_1[2921]; 
    assign out[1271] = layer_1[3159] ^ layer_1[3078]; 
    assign out[1272] = ~(layer_1[3009] | layer_1[3031]); 
    assign out[1273] = layer_1[2131] ^ layer_1[2073]; 
    assign out[1274] = ~layer_1[842]; 
    assign out[1275] = ~layer_1[379] | (layer_1[379] & layer_1[423]); 
    assign out[1276] = layer_1[344] & ~layer_1[253]; 
    assign out[1277] = layer_1[2370] & ~layer_1[2466]; 
    assign out[1278] = ~layer_1[200]; 
    assign out[1279] = layer_1[362]; 
    assign out[1280] = layer_1[14] | layer_1[46]; 
    assign out[1281] = layer_1[841]; 
    assign out[1282] = layer_1[2833] | layer_1[2755]; 
    assign out[1283] = layer_1[985] & ~layer_1[1069]; 
    assign out[1284] = layer_1[740] & layer_1[700]; 
    assign out[1285] = layer_1[1102] ^ layer_1[1142]; 
    assign out[1286] = ~(layer_1[3945] ^ layer_1[3940]); 
    assign out[1287] = layer_1[3413] | layer_1[3471]; 
    assign out[1288] = layer_1[911]; 
    assign out[1289] = layer_1[886]; 
    assign out[1290] = ~layer_1[2514] | (layer_1[2443] & layer_1[2514]); 
    assign out[1291] = ~(layer_1[478] ^ layer_1[384]); 
    assign out[1292] = ~(layer_1[127] ^ layer_1[226]); 
    assign out[1293] = ~layer_1[3826] | (layer_1[3826] & layer_1[3884]); 
    assign out[1294] = layer_1[460]; 
    assign out[1295] = ~layer_1[3190]; 
    assign out[1296] = layer_1[2768] | layer_1[2759]; 
    assign out[1297] = layer_1[2499] ^ layer_1[2607]; 
    assign out[1298] = ~(layer_1[3723] | layer_1[3745]); 
    assign out[1299] = ~layer_1[1493]; 
    assign out[1300] = ~layer_1[1133]; 
    assign out[1301] = ~(layer_1[236] | layer_1[224]); 
    assign out[1302] = layer_1[2059]; 
    assign out[1303] = ~(layer_1[2465] | layer_1[2530]); 
    assign out[1304] = ~(layer_1[1636] | layer_1[1756]); 
    assign out[1305] = layer_1[1083] & layer_1[1174]; 
    assign out[1306] = layer_1[541] & ~layer_1[462]; 
    assign out[1307] = ~layer_1[2635]; 
    assign out[1308] = ~layer_1[1687]; 
    assign out[1309] = layer_1[2409] ^ layer_1[2391]; 
    assign out[1310] = layer_1[2938] ^ layer_1[2885]; 
    assign out[1311] = layer_1[324]; 
    assign out[1312] = ~layer_1[2730] | (layer_1[2730] & layer_1[2818]); 
    assign out[1313] = layer_1[757] & ~layer_1[870]; 
    assign out[1314] = ~(layer_1[2074] ^ layer_1[2032]); 
    assign out[1315] = layer_1[2706] & ~layer_1[2592]; 
    assign out[1316] = ~(layer_1[2403] | layer_1[2301]); 
    assign out[1317] = ~(layer_1[2125] ^ layer_1[2011]); 
    assign out[1318] = ~layer_1[2734]; 
    assign out[1319] = ~layer_1[1175]; 
    assign out[1320] = ~(layer_1[1622] ^ layer_1[1542]); 
    assign out[1321] = layer_1[3131] ^ layer_1[3083]; 
    assign out[1322] = layer_1[3037] & layer_1[3023]; 
    assign out[1323] = layer_1[2253] & ~layer_1[2315]; 
    assign out[1324] = ~layer_1[2477]; 
    assign out[1325] = ~layer_1[2403]; 
    assign out[1326] = ~(layer_1[1827] & layer_1[1736]); 
    assign out[1327] = ~layer_1[282] | (layer_1[282] & layer_1[321]); 
    assign out[1328] = ~layer_1[3306]; 
    assign out[1329] = layer_1[1369] & layer_1[1443]; 
    assign out[1330] = ~(layer_1[138] | layer_1[264]); 
    assign out[1331] = ~(layer_1[2208] ^ layer_1[2184]); 
    assign out[1332] = ~layer_1[3289] | (layer_1[3289] & layer_1[3250]); 
    assign out[1333] = layer_1[333] | layer_1[230]; 
    assign out[1334] = layer_1[2147]; 
    assign out[1335] = ~(layer_1[676] ^ layer_1[575]); 
    assign out[1336] = layer_1[3946] ^ layer_1[3992]; 
    assign out[1337] = layer_1[2256]; 
    assign out[1338] = ~layer_1[2156]; 
    assign out[1339] = layer_1[814] ^ layer_1[714]; 
    assign out[1340] = layer_1[1801] & layer_1[1785]; 
    assign out[1341] = layer_1[3239] & ~layer_1[3136]; 
    assign out[1342] = layer_1[1343] & layer_1[1414]; 
    assign out[1343] = layer_1[765] ^ layer_1[736]; 
    assign out[1344] = layer_1[2167]; 
    assign out[1345] = ~layer_1[491]; 
    assign out[1346] = layer_1[479] ^ layer_1[452]; 
    assign out[1347] = layer_1[2365] & layer_1[2272]; 
    assign out[1348] = ~layer_1[2647]; 
    assign out[1349] = layer_1[1304]; 
    assign out[1350] = layer_1[2824] & ~layer_1[2723]; 
    assign out[1351] = layer_1[2854] & ~layer_1[2787]; 
    assign out[1352] = layer_1[192] ^ layer_1[202]; 
    assign out[1353] = ~(layer_1[1954] ^ layer_1[1893]); 
    assign out[1354] = layer_1[3873]; 
    assign out[1355] = ~(layer_1[3907] & layer_1[3966]); 
    assign out[1356] = layer_1[495]; 
    assign out[1357] = layer_1[3503]; 
    assign out[1358] = ~layer_1[769] | (layer_1[769] & layer_1[836]); 
    assign out[1359] = layer_1[2917] & ~layer_1[2973]; 
    assign out[1360] = ~(layer_1[3367] ^ layer_1[3421]); 
    assign out[1361] = layer_1[2549] & layer_1[2639]; 
    assign out[1362] = ~(layer_1[2394] ^ layer_1[2490]); 
    assign out[1363] = ~layer_1[1015] | (layer_1[1015] & layer_1[1141]); 
    assign out[1364] = ~(layer_1[2396] | layer_1[2492]); 
    assign out[1365] = ~(layer_1[1798] ^ layer_1[1702]); 
    assign out[1366] = ~(layer_1[1366] ^ layer_1[1240]); 
    assign out[1367] = ~layer_1[1910]; 
    assign out[1368] = layer_1[1572] | layer_1[1478]; 
    assign out[1369] = ~(layer_1[1507] | layer_1[1457]); 
    assign out[1370] = layer_1[468]; 
    assign out[1371] = layer_1[1187]; 
    assign out[1372] = ~(layer_1[518] ^ layer_1[582]); 
    assign out[1373] = ~(layer_1[3429] | layer_1[3469]); 
    assign out[1374] = layer_1[2124] ^ layer_1[2166]; 
    assign out[1375] = ~layer_1[2031]; 
    assign out[1376] = layer_1[277] ^ layer_1[358]; 
    assign out[1377] = layer_1[2963]; 
    assign out[1378] = ~layer_1[3724]; 
    assign out[1379] = layer_1[3476] | layer_1[3357]; 
    assign out[1380] = ~(layer_1[2362] | layer_1[2396]); 
    assign out[1381] = layer_1[3706] & layer_1[3739]; 
    assign out[1382] = layer_1[3979]; 
    assign out[1383] = ~(layer_1[3786] ^ layer_1[3735]); 
    assign out[1384] = ~(layer_1[392] | layer_1[506]); 
    assign out[1385] = layer_1[2071]; 
    assign out[1386] = layer_1[2561]; 
    assign out[1387] = ~layer_1[57]; 
    assign out[1388] = ~layer_1[2556]; 
    assign out[1389] = ~(layer_1[2192] ^ layer_1[2236]); 
    assign out[1390] = ~(layer_1[1578] & layer_1[1595]); 
    assign out[1391] = layer_1[635] & ~layer_1[606]; 
    assign out[1392] = layer_1[1626] & ~layer_1[1693]; 
    assign out[1393] = layer_1[3994] & ~layer_1[3951]; 
    assign out[1394] = layer_1[2310] & ~layer_1[2259]; 
    assign out[1395] = layer_1[3597]; 
    assign out[1396] = layer_1[3669]; 
    assign out[1397] = layer_1[2050] ^ layer_1[1972]; 
    assign out[1398] = layer_1[2008] ^ layer_1[2023]; 
    assign out[1399] = ~layer_1[2463]; 
    assign out[1400] = ~layer_1[1435] | (layer_1[1435] & layer_1[1465]); 
    assign out[1401] = layer_1[1010]; 
    assign out[1402] = layer_1[3024]; 
    assign out[1403] = ~layer_1[1]; 
    assign out[1404] = ~(layer_1[1277] | layer_1[1246]); 
    assign out[1405] = ~layer_1[2274]; 
    assign out[1406] = layer_1[385] ^ layer_1[443]; 
    assign out[1407] = ~layer_1[2961]; 
    assign out[1408] = layer_1[2912]; 
    assign out[1409] = ~(layer_1[3018] ^ layer_1[3123]); 
    assign out[1410] = layer_1[138] ^ layer_1[112]; 
    assign out[1411] = layer_1[2738]; 
    assign out[1412] = layer_1[993] ^ layer_1[907]; 
    assign out[1413] = ~layer_1[1930] | (layer_1[1930] & layer_1[1880]); 
    assign out[1414] = ~layer_1[3527] | (layer_1[3490] & layer_1[3527]); 
    assign out[1415] = ~layer_1[1]; 
    assign out[1416] = layer_1[330] & layer_1[342]; 
    assign out[1417] = layer_1[1034] ^ layer_1[1071]; 
    assign out[1418] = ~(layer_1[448] | layer_1[354]); 
    assign out[1419] = layer_1[2965] ^ layer_1[3049]; 
    assign out[1420] = layer_1[2387]; 
    assign out[1421] = ~(layer_1[522] | layer_1[501]); 
    assign out[1422] = layer_1[2559]; 
    assign out[1423] = layer_1[3795] & ~layer_1[3712]; 
    assign out[1424] = layer_1[1136] & ~layer_1[1085]; 
    assign out[1425] = layer_1[3022] ^ layer_1[3021]; 
    assign out[1426] = ~layer_1[1550] | (layer_1[1513] & layer_1[1550]); 
    assign out[1427] = ~layer_1[2694]; 
    assign out[1428] = layer_1[1690]; 
    assign out[1429] = ~layer_1[1658]; 
    assign out[1430] = layer_1[2272] ^ layer_1[2364]; 
    assign out[1431] = ~(layer_1[1031] ^ layer_1[1092]); 
    assign out[1432] = ~layer_1[2180]; 
    assign out[1433] = layer_1[520]; 
    assign out[1434] = ~layer_1[2867]; 
    assign out[1435] = layer_1[1664] ^ layer_1[1559]; 
    assign out[1436] = ~(layer_1[1448] & layer_1[1355]); 
    assign out[1437] = ~layer_1[953]; 
    assign out[1438] = ~(layer_1[588] & layer_1[534]); 
    assign out[1439] = layer_1[3618] ^ layer_1[3650]; 
    assign out[1440] = ~layer_1[2432]; 
    assign out[1441] = ~layer_1[1133]; 
    assign out[1442] = layer_1[3201] & layer_1[3211]; 
    assign out[1443] = ~(layer_1[779] ^ layer_1[807]); 
    assign out[1444] = layer_1[1472] & ~layer_1[1401]; 
    assign out[1445] = ~layer_1[1802] | (layer_1[1877] & layer_1[1802]); 
    assign out[1446] = layer_1[2735] ^ layer_1[2698]; 
    assign out[1447] = layer_1[2572] & ~layer_1[2632]; 
    assign out[1448] = layer_1[2310] & layer_1[2224]; 
    assign out[1449] = layer_1[340] & layer_1[227]; 
    assign out[1450] = ~layer_1[2881]; 
    assign out[1451] = ~layer_1[3041] | (layer_1[3041] & layer_1[3023]); 
    assign out[1452] = ~layer_1[1033]; 
    assign out[1453] = layer_1[3957]; 
    assign out[1454] = layer_1[1843] & layer_1[1941]; 
    assign out[1455] = ~layer_1[1082] | (layer_1[982] & layer_1[1082]); 
    assign out[1456] = ~layer_1[1278]; 
    assign out[1457] = ~layer_1[3846]; 
    assign out[1458] = layer_1[2567] | layer_1[2633]; 
    assign out[1459] = layer_1[3336] | layer_1[3447]; 
    assign out[1460] = layer_1[674] & layer_1[591]; 
    assign out[1461] = layer_1[417] ^ layer_1[298]; 
    assign out[1462] = layer_1[2799]; 
    assign out[1463] = ~layer_1[2653] | (layer_1[2653] & layer_1[2605]); 
    assign out[1464] = layer_1[1877] | layer_1[1820]; 
    assign out[1465] = layer_1[2075]; 
    assign out[1466] = layer_1[2024] & layer_1[2078]; 
    assign out[1467] = layer_1[2908] | layer_1[2878]; 
    assign out[1468] = ~layer_1[3744]; 
    assign out[1469] = layer_1[3776] | layer_1[3839]; 
    assign out[1470] = layer_1[3093] & ~layer_1[3191]; 
    assign out[1471] = layer_1[2516] & ~layer_1[2612]; 
    assign out[1472] = ~layer_1[846]; 
    assign out[1473] = ~(layer_1[3082] | layer_1[3191]); 
    assign out[1474] = layer_1[1195]; 
    assign out[1475] = ~(layer_1[2046] ^ layer_1[2119]); 
    assign out[1476] = ~(layer_1[755] | layer_1[690]); 
    assign out[1477] = ~layer_1[2951]; 
    assign out[1478] = layer_1[2397] & ~layer_1[2489]; 
    assign out[1479] = ~(layer_1[3788] & layer_1[3697]); 
    assign out[1480] = layer_1[1048]; 
    assign out[1481] = ~layer_1[620] | (layer_1[620] & layer_1[646]); 
    assign out[1482] = ~layer_1[1838] | (layer_1[1953] & layer_1[1838]); 
    assign out[1483] = layer_1[2908]; 
    assign out[1484] = layer_1[3844]; 
    assign out[1485] = ~layer_1[3018] | (layer_1[2938] & layer_1[3018]); 
    assign out[1486] = layer_1[1007] & ~layer_1[922]; 
    assign out[1487] = layer_1[2799]; 
    assign out[1488] = layer_1[2780]; 
    assign out[1489] = layer_1[34] & layer_1[94]; 
    assign out[1490] = layer_1[317] & ~layer_1[437]; 
    assign out[1491] = ~layer_1[3311] | (layer_1[3311] & layer_1[3194]); 
    assign out[1492] = layer_1[2172] ^ layer_1[2286]; 
    assign out[1493] = ~(layer_1[1787] ^ layer_1[1753]); 
    assign out[1494] = ~layer_1[568] | (layer_1[635] & layer_1[568]); 
    assign out[1495] = layer_1[2243] & layer_1[2252]; 
    assign out[1496] = layer_1[34] & ~layer_1[11]; 
    assign out[1497] = layer_1[3642] & layer_1[3660]; 
    assign out[1498] = layer_1[2984] & ~layer_1[3052]; 
    assign out[1499] = layer_1[2014] | layer_1[1991]; 
    assign out[1500] = layer_1[3881]; 
    assign out[1501] = layer_1[2784]; 
    assign out[1502] = layer_1[1645]; 
    assign out[1503] = ~(layer_1[3275] ^ layer_1[3232]); 
    assign out[1504] = ~layer_1[687]; 
    assign out[1505] = layer_1[1051]; 
    assign out[1506] = layer_1[3896]; 
    assign out[1507] = layer_1[734] & ~layer_1[804]; 
    assign out[1508] = layer_1[2862]; 
    assign out[1509] = layer_1[1729]; 
    assign out[1510] = layer_1[2724] | layer_1[2642]; 
    assign out[1511] = layer_1[3916]; 
    assign out[1512] = ~layer_1[437]; 
    assign out[1513] = ~(layer_1[834] ^ layer_1[741]); 
    assign out[1514] = layer_1[1301] | layer_1[1380]; 
    assign out[1515] = ~layer_1[697]; 
    assign out[1516] = ~layer_1[116]; 
    assign out[1517] = ~(layer_1[1321] ^ layer_1[1344]); 
    assign out[1518] = layer_1[2368]; 
    assign out[1519] = ~(layer_1[1424] ^ layer_1[1524]); 
    assign out[1520] = layer_1[2007]; 
    assign out[1521] = layer_1[1117]; 
    assign out[1522] = layer_1[556]; 
    assign out[1523] = layer_1[2606]; 
    assign out[1524] = layer_1[1645] & layer_1[1615]; 
    assign out[1525] = layer_1[2334]; 
    assign out[1526] = ~layer_1[1239]; 
    assign out[1527] = ~(layer_1[2720] | layer_1[2776]); 
    assign out[1528] = layer_1[1605] & layer_1[1615]; 
    assign out[1529] = layer_1[463]; 
    assign out[1530] = ~layer_1[2876]; 
    assign out[1531] = layer_1[2122] ^ layer_1[2023]; 
    assign out[1532] = ~layer_1[1980] | (layer_1[1980] & layer_1[2018]); 
    assign out[1533] = layer_1[3350]; 
    assign out[1534] = ~(layer_1[1628] ^ layer_1[1647]); 
    assign out[1535] = layer_1[2505] ^ layer_1[2500]; 
    assign out[1536] = layer_1[2451] ^ layer_1[2452]; 
    assign out[1537] = layer_1[1302] & ~layer_1[1395]; 
    assign out[1538] = ~(layer_1[57] ^ layer_1[153]); 
    assign out[1539] = layer_1[1341]; 
    assign out[1540] = layer_1[350]; 
    assign out[1541] = layer_1[6] & layer_1[90]; 
    assign out[1542] = layer_1[2921]; 
    assign out[1543] = ~(layer_1[2314] ^ layer_1[2400]); 
    assign out[1544] = layer_1[2612] ^ layer_1[2609]; 
    assign out[1545] = ~(layer_1[2247] ^ layer_1[2157]); 
    assign out[1546] = ~layer_1[292]; 
    assign out[1547] = ~(layer_1[2400] & layer_1[2354]); 
    assign out[1548] = ~layer_1[748]; 
    assign out[1549] = layer_1[2358] & ~layer_1[2471]; 
    assign out[1550] = layer_1[1285]; 
    assign out[1551] = layer_1[3773]; 
    assign out[1552] = layer_1[1842]; 
    assign out[1553] = ~(layer_1[803] ^ layer_1[739]); 
    assign out[1554] = ~layer_1[2042]; 
    assign out[1555] = ~layer_1[3516] | (layer_1[3503] & layer_1[3516]); 
    assign out[1556] = ~layer_1[2035] | (layer_1[2035] & layer_1[2034]); 
    assign out[1557] = layer_1[2676] & ~layer_1[2652]; 
    assign out[1558] = ~layer_1[1461]; 
    assign out[1559] = ~layer_1[620]; 
    assign out[1560] = layer_1[3000] ^ layer_1[3079]; 
    assign out[1561] = ~(layer_1[970] | layer_1[953]); 
    assign out[1562] = ~layer_1[821]; 
    assign out[1563] = ~layer_1[2452] | (layer_1[2424] & layer_1[2452]); 
    assign out[1564] = ~layer_1[1489] | (layer_1[1489] & layer_1[1368]); 
    assign out[1565] = ~(layer_1[3209] | layer_1[3276]); 
    assign out[1566] = layer_1[1206] | layer_1[1241]; 
    assign out[1567] = layer_1[2713]; 
    assign out[1568] = layer_1[1830] & ~layer_1[1958]; 
    assign out[1569] = layer_1[2990] & ~layer_1[2969]; 
    assign out[1570] = layer_1[3388]; 
    assign out[1571] = ~layer_1[2145]; 
    assign out[1572] = ~(layer_1[2275] & layer_1[2326]); 
    assign out[1573] = ~(layer_1[2125] ^ layer_1[2213]); 
    assign out[1574] = ~layer_1[1838] | (layer_1[1838] & layer_1[1729]); 
    assign out[1575] = ~layer_1[1966]; 
    assign out[1576] = layer_1[107] ^ layer_1[163]; 
    assign out[1577] = layer_1[1283] ^ layer_1[1372]; 
    assign out[1578] = layer_1[260]; 
    assign out[1579] = layer_1[1261] & layer_1[1262]; 
    assign out[1580] = layer_1[3573] ^ layer_1[3665]; 
    assign out[1581] = layer_1[509] ^ layer_1[500]; 
    assign out[1582] = ~(layer_1[2437] ^ layer_1[2412]); 
    assign out[1583] = ~(layer_1[810] | layer_1[736]); 
    assign out[1584] = layer_1[2271] ^ layer_1[2265]; 
    assign out[1585] = ~layer_1[2534]; 
    assign out[1586] = layer_1[1954] & ~layer_1[2074]; 
    assign out[1587] = layer_1[1908] & layer_1[1896]; 
    assign out[1588] = ~(layer_1[881] ^ layer_1[816]); 
    assign out[1589] = ~(layer_1[3964] ^ layer_1[3940]); 
    assign out[1590] = layer_1[1876] & layer_1[2004]; 
    assign out[1591] = ~layer_1[3428]; 
    assign out[1592] = layer_1[2338] & layer_1[2437]; 
    assign out[1593] = layer_1[1137] | layer_1[1141]; 
    assign out[1594] = layer_1[88]; 
    assign out[1595] = layer_1[3259] & ~layer_1[3320]; 
    assign out[1596] = ~(layer_1[3682] & layer_1[3559]); 
    assign out[1597] = ~layer_1[2734]; 
    assign out[1598] = ~(layer_1[3127] ^ layer_1[3038]); 
    assign out[1599] = layer_1[1435] & ~layer_1[1557]; 
    assign out[1600] = layer_1[2927]; 
    assign out[1601] = layer_1[1118] & ~layer_1[992]; 
    assign out[1602] = layer_1[270] & ~layer_1[202]; 
    assign out[1603] = layer_1[2918]; 
    assign out[1604] = layer_1[3826] & ~layer_1[3791]; 
    assign out[1605] = layer_1[2518]; 
    assign out[1606] = ~(layer_1[3291] & layer_1[3366]); 
    assign out[1607] = layer_1[2365] & ~layer_1[2445]; 
    assign out[1608] = ~layer_1[3066]; 
    assign out[1609] = layer_1[3429] & ~layer_1[3544]; 
    assign out[1610] = ~layer_1[2052]; 
    assign out[1611] = layer_1[832] & layer_1[750]; 
    assign out[1612] = ~(layer_1[1314] ^ layer_1[1209]); 
    assign out[1613] = layer_1[3064] ^ layer_1[2995]; 
    assign out[1614] = ~(layer_1[183] | layer_1[202]); 
    assign out[1615] = ~(layer_1[1065] | layer_1[1132]); 
    assign out[1616] = ~layer_1[1042]; 
    assign out[1617] = layer_1[3735] & layer_1[3707]; 
    assign out[1618] = layer_1[1011] & ~layer_1[1023]; 
    assign out[1619] = layer_1[237] & layer_1[289]; 
    assign out[1620] = layer_1[2926]; 
    assign out[1621] = layer_1[3764]; 
    assign out[1622] = layer_1[2933]; 
    assign out[1623] = layer_1[3008] & ~layer_1[2917]; 
    assign out[1624] = ~(layer_1[7] | layer_1[1]); 
    assign out[1625] = layer_1[653] & ~layer_1[652]; 
    assign out[1626] = ~layer_1[3012]; 
    assign out[1627] = ~(layer_1[2659] ^ layer_1[2655]); 
    assign out[1628] = ~layer_1[3944]; 
    assign out[1629] = layer_1[287] & ~layer_1[229]; 
    assign out[1630] = ~layer_1[580]; 
    assign out[1631] = ~(layer_1[531] | layer_1[452]); 
    assign out[1632] = ~(layer_1[1031] ^ layer_1[939]); 
    assign out[1633] = ~layer_1[2072] | (layer_1[2020] & layer_1[2072]); 
    assign out[1634] = layer_1[1911] ^ layer_1[1855]; 
    assign out[1635] = layer_1[1037] ^ layer_1[1144]; 
    assign out[1636] = ~(layer_1[3476] | layer_1[3481]); 
    assign out[1637] = ~(layer_1[3388] | layer_1[3318]); 
    assign out[1638] = layer_1[2262] ^ layer_1[2379]; 
    assign out[1639] = layer_1[3005] ^ layer_1[2996]; 
    assign out[1640] = layer_1[771] & layer_1[820]; 
    assign out[1641] = ~(layer_1[2121] ^ layer_1[2058]); 
    assign out[1642] = layer_1[324] ^ layer_1[406]; 
    assign out[1643] = layer_1[371] & layer_1[401]; 
    assign out[1644] = ~(layer_1[2442] ^ layer_1[2564]); 
    assign out[1645] = ~(layer_1[3860] | layer_1[3979]); 
    assign out[1646] = layer_1[1498] ^ layer_1[1395]; 
    assign out[1647] = layer_1[3360]; 
    assign out[1648] = layer_1[432] & ~layer_1[350]; 
    assign out[1649] = layer_1[3909]; 
    assign out[1650] = layer_1[2448] & layer_1[2489]; 
    assign out[1651] = ~layer_1[1463]; 
    assign out[1652] = layer_1[1352]; 
    assign out[1653] = layer_1[5] & ~layer_1[15]; 
    assign out[1654] = layer_1[3711] & layer_1[3694]; 
    assign out[1655] = ~(layer_1[355] & layer_1[299]); 
    assign out[1656] = layer_1[2551] & ~layer_1[2663]; 
    assign out[1657] = layer_1[1927] & ~layer_1[1805]; 
    assign out[1658] = layer_1[1488] & layer_1[1505]; 
    assign out[1659] = ~(layer_1[3943] ^ layer_1[3970]); 
    assign out[1660] = layer_1[2674] & ~layer_1[2663]; 
    assign out[1661] = ~(layer_1[1728] | layer_1[1702]); 
    assign out[1662] = layer_1[3850] ^ layer_1[3843]; 
    assign out[1663] = layer_1[2982] & ~layer_1[2923]; 
    assign out[1664] = layer_1[1190] ^ layer_1[1295]; 
    assign out[1665] = ~layer_1[3573]; 
    assign out[1666] = ~layer_1[3364] | (layer_1[3486] & layer_1[3364]); 
    assign out[1667] = layer_1[3710] & layer_1[3762]; 
    assign out[1668] = layer_1[2908] | layer_1[2848]; 
    assign out[1669] = ~layer_1[12]; 
    assign out[1670] = ~(layer_1[1779] | layer_1[1894]); 
    assign out[1671] = layer_1[583] ^ layer_1[527]; 
    assign out[1672] = ~layer_1[1968]; 
    assign out[1673] = layer_1[3072] & ~layer_1[3123]; 
    assign out[1674] = layer_1[2275] & ~layer_1[2180]; 
    assign out[1675] = ~layer_1[2749] | (layer_1[2636] & layer_1[2749]); 
    assign out[1676] = ~(layer_1[3286] ^ layer_1[3280]); 
    assign out[1677] = layer_1[2952] & ~layer_1[3063]; 
    assign out[1678] = layer_1[904] ^ layer_1[934]; 
    assign out[1679] = layer_1[1438] & ~layer_1[1511]; 
    assign out[1680] = ~layer_1[3349] | (layer_1[3308] & layer_1[3349]); 
    assign out[1681] = ~(layer_1[3493] | layer_1[3517]); 
    assign out[1682] = layer_1[3761] & ~layer_1[3746]; 
    assign out[1683] = ~layer_1[9]; 
    assign out[1684] = ~(layer_1[1343] & layer_1[1452]); 
    assign out[1685] = layer_1[2117] & ~layer_1[2129]; 
    assign out[1686] = layer_1[41] & layer_1[128]; 
    assign out[1687] = ~layer_1[659]; 
    assign out[1688] = ~(layer_1[1823] ^ layer_1[1809]); 
    assign out[1689] = layer_1[3650] ^ layer_1[3613]; 
    assign out[1690] = layer_1[1631] & ~layer_1[1728]; 
    assign out[1691] = ~layer_1[1177]; 
    assign out[1692] = layer_1[3013]; 
    assign out[1693] = ~(layer_1[3518] ^ layer_1[3469]); 
    assign out[1694] = layer_1[1155]; 
    assign out[1695] = layer_1[1952] ^ layer_1[1982]; 
    assign out[1696] = ~layer_1[3455]; 
    assign out[1697] = layer_1[837]; 
    assign out[1698] = ~(layer_1[992] ^ layer_1[1007]); 
    assign out[1699] = ~(layer_1[2892] ^ layer_1[2962]); 
    assign out[1700] = ~layer_1[530]; 
    assign out[1701] = layer_1[777] & ~layer_1[814]; 
    assign out[1702] = ~layer_1[848]; 
    assign out[1703] = ~(layer_1[961] ^ layer_1[940]); 
    assign out[1704] = layer_1[1902]; 
    assign out[1705] = ~layer_1[3622] | (layer_1[3661] & layer_1[3622]); 
    assign out[1706] = layer_1[887]; 
    assign out[1707] = ~layer_1[2786] | (layer_1[2773] & layer_1[2786]); 
    assign out[1708] = layer_1[865] | layer_1[875]; 
    assign out[1709] = layer_1[3213]; 
    assign out[1710] = ~(layer_1[467] ^ layer_1[507]); 
    assign out[1711] = ~layer_1[3394] | (layer_1[3435] & layer_1[3394]); 
    assign out[1712] = ~layer_1[2879]; 
    assign out[1713] = ~layer_1[3592] | (layer_1[3592] & layer_1[3621]); 
    assign out[1714] = layer_1[1844] & layer_1[1759]; 
    assign out[1715] = ~layer_1[479] | (layer_1[513] & layer_1[479]); 
    assign out[1716] = layer_1[3100] ^ layer_1[3033]; 
    assign out[1717] = layer_1[2980] & ~layer_1[2886]; 
    assign out[1718] = ~(layer_1[2147] ^ layer_1[2211]); 
    assign out[1719] = layer_1[249]; 
    assign out[1720] = ~(layer_1[2798] & layer_1[2705]); 
    assign out[1721] = layer_1[2045]; 
    assign out[1722] = layer_1[922] & ~layer_1[971]; 
    assign out[1723] = ~layer_1[373] | (layer_1[405] & layer_1[373]); 
    assign out[1724] = ~(layer_1[1430] & layer_1[1550]); 
    assign out[1725] = ~(layer_1[2823] ^ layer_1[2817]); 
    assign out[1726] = layer_1[3056] | layer_1[3057]; 
    assign out[1727] = layer_1[1625] & ~layer_1[1541]; 
    assign out[1728] = layer_1[217] ^ layer_1[242]; 
    assign out[1729] = layer_1[1464] & layer_1[1576]; 
    assign out[1730] = ~(layer_1[1127] ^ layer_1[1156]); 
    assign out[1731] = ~layer_1[123]; 
    assign out[1732] = ~layer_1[3831] | (layer_1[3918] & layer_1[3831]); 
    assign out[1733] = ~(layer_1[3219] ^ layer_1[3228]); 
    assign out[1734] = ~(layer_1[2730] & layer_1[2701]); 
    assign out[1735] = ~(layer_1[3519] | layer_1[3591]); 
    assign out[1736] = layer_1[2132] ^ layer_1[2101]; 
    assign out[1737] = ~(layer_1[490] ^ layer_1[531]); 
    assign out[1738] = layer_1[3148] ^ layer_1[3132]; 
    assign out[1739] = ~(layer_1[2682] | layer_1[2774]); 
    assign out[1740] = layer_1[2659] & layer_1[2714]; 
    assign out[1741] = layer_1[834] | layer_1[820]; 
    assign out[1742] = ~layer_1[1268]; 
    assign out[1743] = ~(layer_1[1698] ^ layer_1[1581]); 
    assign out[1744] = ~layer_1[1315]; 
    assign out[1745] = layer_1[292] & layer_1[365]; 
    assign out[1746] = ~(layer_1[3224] | layer_1[3115]); 
    assign out[1747] = layer_1[3479]; 
    assign out[1748] = layer_1[2443] & ~layer_1[2342]; 
    assign out[1749] = layer_1[1813] ^ layer_1[1750]; 
    assign out[1750] = layer_1[2346]; 
    assign out[1751] = layer_1[3820] & ~layer_1[3941]; 
    assign out[1752] = layer_1[1764]; 
    assign out[1753] = layer_1[3158]; 
    assign out[1754] = layer_1[84] ^ layer_1[144]; 
    assign out[1755] = ~layer_1[2736] | (layer_1[2856] & layer_1[2736]); 
    assign out[1756] = layer_1[1785]; 
    assign out[1757] = layer_1[54] ^ layer_1[158]; 
    assign out[1758] = layer_1[3483]; 
    assign out[1759] = ~layer_1[3693]; 
    assign out[1760] = ~layer_1[2824] | (layer_1[2732] & layer_1[2824]); 
    assign out[1761] = ~(layer_1[28] & layer_1[30]); 
    assign out[1762] = layer_1[3313] ^ layer_1[3361]; 
    assign out[1763] = ~(layer_1[1843] ^ layer_1[1797]); 
    assign out[1764] = ~layer_1[3721] | (layer_1[3719] & layer_1[3721]); 
    assign out[1765] = layer_1[3601]; 
    assign out[1766] = ~layer_1[2768]; 
    assign out[1767] = ~layer_1[3498]; 
    assign out[1768] = layer_1[287] & ~layer_1[376]; 
    assign out[1769] = ~(layer_1[3891] ^ layer_1[3773]); 
    assign out[1770] = ~layer_1[3506] | (layer_1[3506] & layer_1[3503]); 
    assign out[1771] = layer_1[2565] & layer_1[2540]; 
    assign out[1772] = layer_1[3480] ^ layer_1[3494]; 
    assign out[1773] = ~(layer_1[1650] ^ layer_1[1706]); 
    assign out[1774] = layer_1[1372] & ~layer_1[1469]; 
    assign out[1775] = ~layer_1[3115]; 
    assign out[1776] = layer_1[1404] & ~layer_1[1377]; 
    assign out[1777] = layer_1[3057]; 
    assign out[1778] = layer_1[3194] & layer_1[3170]; 
    assign out[1779] = ~(layer_1[2735] ^ layer_1[2843]); 
    assign out[1780] = layer_1[1098] ^ layer_1[1093]; 
    assign out[1781] = ~(layer_1[2187] ^ layer_1[2230]); 
    assign out[1782] = layer_1[2046]; 
    assign out[1783] = layer_1[2381] & layer_1[2411]; 
    assign out[1784] = layer_1[3452] & ~layer_1[3526]; 
    assign out[1785] = layer_1[2927]; 
    assign out[1786] = layer_1[797] & ~layer_1[873]; 
    assign out[1787] = ~(layer_1[1399] | layer_1[1278]); 
    assign out[1788] = layer_1[3286] & layer_1[3309]; 
    assign out[1789] = layer_1[2119] & ~layer_1[2058]; 
    assign out[1790] = layer_1[3771]; 
    assign out[1791] = layer_1[2570] & ~layer_1[2471]; 
    assign out[1792] = layer_1[3202]; 
    assign out[1793] = ~(layer_1[1898] | layer_1[1931]); 
    assign out[1794] = layer_1[1821]; 
    assign out[1795] = ~layer_1[2115]; 
    assign out[1796] = layer_1[166]; 
    assign out[1797] = ~layer_1[2057]; 
    assign out[1798] = ~layer_1[564]; 
    assign out[1799] = ~layer_1[159] | (layer_1[159] & layer_1[79]); 
    assign out[1800] = layer_1[2442] & ~layer_1[2536]; 
    assign out[1801] = ~(layer_1[1226] | layer_1[1218]); 
    assign out[1802] = layer_1[1742] & layer_1[1780]; 
    assign out[1803] = layer_1[3169]; 
    assign out[1804] = layer_1[1139]; 
    assign out[1805] = ~(layer_1[826] ^ layer_1[771]); 
    assign out[1806] = layer_1[3820] | layer_1[3697]; 
    assign out[1807] = ~(layer_1[694] ^ layer_1[668]); 
    assign out[1808] = ~layer_1[2209]; 
    assign out[1809] = layer_1[3849] & ~layer_1[3928]; 
    assign out[1810] = layer_1[1865] & ~layer_1[1779]; 
    assign out[1811] = layer_1[1243] & layer_1[1289]; 
    assign out[1812] = ~(layer_1[3897] ^ layer_1[3927]); 
    assign out[1813] = layer_1[2368]; 
    assign out[1814] = ~(layer_1[651] | layer_1[650]); 
    assign out[1815] = layer_1[3588] & layer_1[3469]; 
    assign out[1816] = ~layer_1[1262]; 
    assign out[1817] = layer_1[1912]; 
    assign out[1818] = layer_1[3210] & layer_1[3245]; 
    assign out[1819] = ~layer_1[3241]; 
    assign out[1820] = ~layer_1[1771] | (layer_1[1771] & layer_1[1653]); 
    assign out[1821] = ~layer_1[3793]; 
    assign out[1822] = layer_1[3158]; 
    assign out[1823] = layer_1[3849]; 
    assign out[1824] = layer_1[1819] & ~layer_1[1915]; 
    assign out[1825] = layer_1[3930] & ~layer_1[3819]; 
    assign out[1826] = layer_1[3176] & ~layer_1[3230]; 
    assign out[1827] = ~(layer_1[1779] | layer_1[1880]); 
    assign out[1828] = layer_1[1452] ^ layer_1[1328]; 
    assign out[1829] = ~layer_1[1640]; 
    assign out[1830] = ~layer_1[2656] | (layer_1[2656] & layer_1[2721]); 
    assign out[1831] = ~layer_1[276]; 
    assign out[1832] = layer_1[417] & ~layer_1[318]; 
    assign out[1833] = layer_1[2721] & ~layer_1[2841]; 
    assign out[1834] = ~(layer_1[1975] ^ layer_1[1953]); 
    assign out[1835] = layer_1[3058] & ~layer_1[3132]; 
    assign out[1836] = layer_1[2806] & layer_1[2726]; 
    assign out[1837] = layer_1[169] | layer_1[178]; 
    assign out[1838] = ~(layer_1[76] & layer_1[148]); 
    assign out[1839] = layer_1[2391] & layer_1[2500]; 
    assign out[1840] = layer_1[1683]; 
    assign out[1841] = ~(layer_1[3247] | layer_1[3238]); 
    assign out[1842] = ~layer_1[1612]; 
    assign out[1843] = ~(layer_1[3844] & layer_1[3848]); 
    assign out[1844] = ~(layer_1[634] ^ layer_1[757]); 
    assign out[1845] = ~(layer_1[3291] ^ layer_1[3211]); 
    assign out[1846] = ~(layer_1[2048] | layer_1[2090]); 
    assign out[1847] = layer_1[1091] & ~layer_1[1164]; 
    assign out[1848] = layer_1[3254]; 
    assign out[1849] = ~(layer_1[3460] ^ layer_1[3418]); 
    assign out[1850] = layer_1[3971]; 
    assign out[1851] = layer_1[1207] ^ layer_1[1205]; 
    assign out[1852] = layer_1[3631] & layer_1[3625]; 
    assign out[1853] = ~layer_1[3108]; 
    assign out[1854] = layer_1[1565] & ~layer_1[1536]; 
    assign out[1855] = layer_1[3420] & ~layer_1[3300]; 
    assign out[1856] = ~(layer_1[185] | layer_1[188]); 
    assign out[1857] = layer_1[1531] & ~layer_1[1415]; 
    assign out[1858] = layer_1[2490] ^ layer_1[2429]; 
    assign out[1859] = layer_1[2257] | layer_1[2232]; 
    assign out[1860] = layer_1[3354] | layer_1[3429]; 
    assign out[1861] = ~layer_1[3922]; 
    assign out[1862] = layer_1[3076] ^ layer_1[3177]; 
    assign out[1863] = layer_1[1813] ^ layer_1[1762]; 
    assign out[1864] = layer_1[1650]; 
    assign out[1865] = layer_1[1663]; 
    assign out[1866] = layer_1[1646] ^ layer_1[1761]; 
    assign out[1867] = layer_1[2492] ^ layer_1[2444]; 
    assign out[1868] = ~(layer_1[3997] | layer_1[3907]); 
    assign out[1869] = ~(layer_1[1811] | layer_1[1935]); 
    assign out[1870] = ~layer_1[3389] | (layer_1[3371] & layer_1[3389]); 
    assign out[1871] = ~(layer_1[2070] | layer_1[1942]); 
    assign out[1872] = layer_1[116]; 
    assign out[1873] = layer_1[2710] & ~layer_1[2625]; 
    assign out[1874] = layer_1[462]; 
    assign out[1875] = ~layer_1[1883]; 
    assign out[1876] = ~(layer_1[1883] | layer_1[1817]); 
    assign out[1877] = layer_1[3710]; 
    assign out[1878] = layer_1[3202] & ~layer_1[3325]; 
    assign out[1879] = layer_1[1755] ^ layer_1[1831]; 
    assign out[1880] = ~layer_1[1242]; 
    assign out[1881] = layer_1[2092] ^ layer_1[2211]; 
    assign out[1882] = ~(layer_1[3890] ^ layer_1[3776]); 
    assign out[1883] = layer_1[3045]; 
    assign out[1884] = ~layer_1[2879]; 
    assign out[1885] = ~(layer_1[481] | layer_1[552]); 
    assign out[1886] = layer_1[2952] & layer_1[3008]; 
    assign out[1887] = ~(layer_1[1608] ^ layer_1[1494]); 
    assign out[1888] = ~(layer_1[3517] ^ layer_1[3518]); 
    assign out[1889] = layer_1[476] & ~layer_1[349]; 
    assign out[1890] = ~layer_1[892]; 
    assign out[1891] = layer_1[1317]; 
    assign out[1892] = ~(layer_1[2780] & layer_1[2701]); 
    assign out[1893] = layer_1[3763]; 
    assign out[1894] = layer_1[3824]; 
    assign out[1895] = ~layer_1[60] | (layer_1[60] & layer_1[2]); 
    assign out[1896] = layer_1[3815]; 
    assign out[1897] = ~layer_1[2824] | (layer_1[2791] & layer_1[2824]); 
    assign out[1898] = layer_1[2500]; 
    assign out[1899] = ~layer_1[1080]; 
    assign out[1900] = ~layer_1[3390]; 
    assign out[1901] = layer_1[3154] & ~layer_1[3123]; 
    assign out[1902] = layer_1[3634] & ~layer_1[3725]; 
    assign out[1903] = layer_1[1886]; 
    assign out[1904] = layer_1[1028]; 
    assign out[1905] = layer_1[958]; 
    assign out[1906] = layer_1[3040] & ~layer_1[2941]; 
    assign out[1907] = layer_1[1996] & layer_1[1872]; 
    assign out[1908] = layer_1[3593] ^ layer_1[3467]; 
    assign out[1909] = ~layer_1[1442]; 
    assign out[1910] = ~(layer_1[2859] ^ layer_1[2962]); 
    assign out[1911] = ~(layer_1[3950] | layer_1[3915]); 
    assign out[1912] = ~layer_1[260] | (layer_1[260] & layer_1[175]); 
    assign out[1913] = layer_1[1155]; 
    assign out[1914] = layer_1[3256] & ~layer_1[3260]; 
    assign out[1915] = layer_1[1356]; 
    assign out[1916] = layer_1[1715]; 
    assign out[1917] = ~(layer_1[3344] ^ layer_1[3386]); 
    assign out[1918] = layer_1[355] ^ layer_1[412]; 
    assign out[1919] = layer_1[282] & layer_1[166]; 
    assign out[1920] = layer_1[771]; 
    assign out[1921] = layer_1[2581] & ~layer_1[2603]; 
    assign out[1922] = ~layer_1[3417]; 
    assign out[1923] = layer_1[2800] | layer_1[2703]; 
    assign out[1924] = ~(layer_1[2279] | layer_1[2180]); 
    assign out[1925] = ~(layer_1[17] ^ layer_1[117]); 
    assign out[1926] = layer_1[2970] & ~layer_1[2910]; 
    assign out[1927] = layer_1[3653] & ~layer_1[3590]; 
    assign out[1928] = ~layer_1[1320]; 
    assign out[1929] = layer_1[355] ^ layer_1[412]; 
    assign out[1930] = layer_1[78] & layer_1[149]; 
    assign out[1931] = layer_1[27]; 
    assign out[1932] = layer_1[2205] & layer_1[2216]; 
    assign out[1933] = ~layer_1[2504]; 
    assign out[1934] = layer_1[3749] & ~layer_1[3836]; 
    assign out[1935] = ~(layer_1[1970] ^ layer_1[1990]); 
    assign out[1936] = ~(layer_1[2527] | layer_1[2522]); 
    assign out[1937] = layer_1[1244] ^ layer_1[1293]; 
    assign out[1938] = ~layer_1[1447]; 
    assign out[1939] = ~(layer_1[1099] | layer_1[1102]); 
    assign out[1940] = layer_1[3949]; 
    assign out[1941] = layer_1[1401] & ~layer_1[1365]; 
    assign out[1942] = ~layer_1[2217]; 
    assign out[1943] = layer_1[1385] & ~layer_1[1418]; 
    assign out[1944] = ~(layer_1[601] | layer_1[616]); 
    assign out[1945] = layer_1[58] & ~layer_1[96]; 
    assign out[1946] = ~(layer_1[3426] | layer_1[3390]); 
    assign out[1947] = ~layer_1[2743]; 
    assign out[1948] = layer_1[2062] & layer_1[2122]; 
    assign out[1949] = ~(layer_1[1869] | layer_1[1977]); 
    assign out[1950] = layer_1[2989]; 
    assign out[1951] = layer_1[1466] ^ layer_1[1574]; 
    assign out[1952] = ~(layer_1[771] ^ layer_1[842]); 
    assign out[1953] = ~layer_1[355]; 
    assign out[1954] = layer_1[654]; 
    assign out[1955] = layer_1[2914]; 
    assign out[1956] = ~(layer_1[142] ^ layer_1[136]); 
    assign out[1957] = ~(layer_1[3901] ^ layer_1[3888]); 
    assign out[1958] = ~(layer_1[1052] ^ layer_1[1137]); 
    assign out[1959] = layer_1[1239] & layer_1[1318]; 
    assign out[1960] = ~(layer_1[1025] ^ layer_1[1051]); 
    assign out[1961] = layer_1[3404] & layer_1[3330]; 
    assign out[1962] = layer_1[3582]; 
    assign out[1963] = layer_1[3868]; 
    assign out[1964] = layer_1[3116] ^ layer_1[3215]; 
    assign out[1965] = ~(layer_1[3577] ^ layer_1[3539]); 
    assign out[1966] = layer_1[1200]; 
    assign out[1967] = ~layer_1[3152]; 
    assign out[1968] = layer_1[3676] & ~layer_1[3794]; 
    assign out[1969] = ~(layer_1[531] & layer_1[543]); 
    assign out[1970] = ~layer_1[2060]; 
    assign out[1971] = ~(layer_1[3652] ^ layer_1[3573]); 
    assign out[1972] = layer_1[56]; 
    assign out[1973] = ~layer_1[200]; 
    assign out[1974] = layer_1[236]; 
    assign out[1975] = ~layer_1[982]; 
    assign out[1976] = layer_1[289]; 
    assign out[1977] = layer_1[2332] ^ layer_1[2270]; 
    assign out[1978] = layer_1[3256]; 
    assign out[1979] = layer_1[1767]; 
    assign out[1980] = ~layer_1[229]; 
    assign out[1981] = layer_1[1946] ^ layer_1[2043]; 
    assign out[1982] = layer_1[589] & ~layer_1[693]; 
    assign out[1983] = layer_1[573] ^ layer_1[529]; 
    assign out[1984] = layer_1[3134] | layer_1[3217]; 
    assign out[1985] = layer_1[1888] ^ layer_1[1779]; 
    assign out[1986] = ~(layer_1[2041] | layer_1[2098]); 
    assign out[1987] = ~layer_1[1984] | (layer_1[1989] & layer_1[1984]); 
    assign out[1988] = ~(layer_1[92] ^ layer_1[67]); 
    assign out[1989] = layer_1[3598]; 
    assign out[1990] = ~(layer_1[3577] ^ layer_1[3502]); 
    assign out[1991] = layer_1[2166] ^ layer_1[2051]; 
    assign out[1992] = layer_1[2641] & ~layer_1[2701]; 
    assign out[1993] = layer_1[1197] & ~layer_1[1254]; 
    assign out[1994] = layer_1[2361] & ~layer_1[2279]; 
    assign out[1995] = layer_1[2990] & layer_1[2885]; 
    assign out[1996] = ~(layer_1[3731] | layer_1[3734]); 
    assign out[1997] = ~layer_1[473]; 
    assign out[1998] = layer_1[3719]; 
    assign out[1999] = ~layer_1[491]; 
    assign out[2000] = layer_1[3290]; 
    assign out[2001] = layer_1[819]; 
    assign out[2002] = ~layer_1[3327]; 
    assign out[2003] = ~layer_1[1612]; 
    assign out[2004] = ~layer_1[636]; 
    assign out[2005] = ~(layer_1[1467] | layer_1[1368]); 
    assign out[2006] = layer_1[2152] & layer_1[2247]; 
    assign out[2007] = ~layer_1[791] | (layer_1[877] & layer_1[791]); 
    assign out[2008] = layer_1[3554] ^ layer_1[3540]; 
    assign out[2009] = layer_1[88]; 
    assign out[2010] = layer_1[3416] & layer_1[3418]; 
    assign out[2011] = ~(layer_1[1081] | layer_1[988]); 
    assign out[2012] = layer_1[109]; 
    assign out[2013] = ~layer_1[1033]; 
    assign out[2014] = ~(layer_1[3825] ^ layer_1[3823]); 
    assign out[2015] = layer_1[555] | layer_1[551]; 
    assign out[2016] = layer_1[514]; 
    assign out[2017] = layer_1[3721]; 
    assign out[2018] = layer_1[2213] & ~layer_1[2317]; 
    assign out[2019] = ~layer_1[2962]; 
    assign out[2020] = ~layer_1[513] | (layer_1[513] & layer_1[502]); 
    assign out[2021] = ~(layer_1[2023] | layer_1[1910]); 
    assign out[2022] = layer_1[3291] ^ layer_1[3287]; 
    assign out[2023] = layer_1[3481]; 
    assign out[2024] = ~layer_1[627]; 
    assign out[2025] = layer_1[2040] ^ layer_1[2078]; 
    assign out[2026] = layer_1[1596] & layer_1[1474]; 
    assign out[2027] = layer_1[1701]; 
    assign out[2028] = layer_1[3003] ^ layer_1[3100]; 
    assign out[2029] = ~layer_1[1630] | (layer_1[1604] & layer_1[1630]); 
    assign out[2030] = ~layer_1[907]; 
    assign out[2031] = layer_1[3021]; 
    assign out[2032] = ~layer_1[2209] | (layer_1[2271] & layer_1[2209]); 
    assign out[2033] = layer_1[3251]; 
    assign out[2034] = ~(layer_1[3844] ^ layer_1[3764]); 
    assign out[2035] = ~(layer_1[1771] ^ layer_1[1699]); 
    assign out[2036] = ~layer_1[3541]; 
    assign out[2037] = ~layer_1[2193]; 
    assign out[2038] = ~(layer_1[2576] ^ layer_1[2486]); 
    assign out[2039] = ~(layer_1[525] ^ layer_1[618]); 
    assign out[2040] = ~layer_1[940] | (layer_1[940] & layer_1[1062]); 
    assign out[2041] = layer_1[1193]; 
    assign out[2042] = layer_1[3138] ^ layer_1[3022]; 
    assign out[2043] = ~layer_1[2329]; 
    assign out[2044] = layer_1[3402] ^ layer_1[3377]; 
    assign out[2045] = ~(layer_1[2497] | layer_1[2467]); 
    assign out[2046] = ~layer_1[1312]; 
    assign out[2047] = layer_1[1284]; 
    assign out[2048] = layer_1[2525]; 
    assign out[2049] = layer_1[2179]; 
    assign out[2050] = ~layer_1[152]; 
    assign out[2051] = ~layer_1[1801]; 
    assign out[2052] = ~(layer_1[2109] & layer_1[2002]); 
    assign out[2053] = layer_1[195] & ~layer_1[183]; 
    assign out[2054] = layer_1[482]; 
    assign out[2055] = ~layer_1[143]; 
    assign out[2056] = ~layer_1[3427]; 
    assign out[2057] = ~layer_1[2864]; 
    assign out[2058] = ~layer_1[965]; 
    assign out[2059] = layer_1[2006] ^ layer_1[2032]; 
    assign out[2060] = ~(layer_1[776] | layer_1[743]); 
    assign out[2061] = ~layer_1[2745]; 
    assign out[2062] = ~layer_1[617]; 
    assign out[2063] = ~layer_1[2552] | (layer_1[2552] & layer_1[2494]); 
    assign out[2064] = layer_1[1406]; 
    assign out[2065] = ~(layer_1[1465] ^ layer_1[1575]); 
    assign out[2066] = ~(layer_1[3004] ^ layer_1[2917]); 
    assign out[2067] = ~layer_1[224]; 
    assign out[2068] = ~layer_1[2065]; 
    assign out[2069] = layer_1[275]; 
    assign out[2070] = ~(layer_1[3491] ^ layer_1[3538]); 
    assign out[2071] = layer_1[334]; 
    assign out[2072] = layer_1[2494] & ~layer_1[2428]; 
    assign out[2073] = ~(layer_1[2850] ^ layer_1[2820]); 
    assign out[2074] = layer_1[1295] ^ layer_1[1335]; 
    assign out[2075] = layer_1[3411] ^ layer_1[3318]; 
    assign out[2076] = ~layer_1[56]; 
    assign out[2077] = layer_1[3619]; 
    assign out[2078] = layer_1[3338]; 
    assign out[2079] = ~layer_1[2535]; 
    assign out[2080] = layer_1[3688] ^ layer_1[3730]; 
    assign out[2081] = layer_1[543]; 
    assign out[2082] = ~(layer_1[2050] ^ layer_1[1991]); 
    assign out[2083] = layer_1[1739] & layer_1[1632]; 
    assign out[2084] = layer_1[1609]; 
    assign out[2085] = layer_1[311] & ~layer_1[363]; 
    assign out[2086] = ~layer_1[1583]; 
    assign out[2087] = layer_1[3563] | layer_1[3582]; 
    assign out[2088] = layer_1[1641] & ~layer_1[1580]; 
    assign out[2089] = ~(layer_1[2029] ^ layer_1[2129]); 
    assign out[2090] = layer_1[3588] | layer_1[3551]; 
    assign out[2091] = ~(layer_1[290] ^ layer_1[172]); 
    assign out[2092] = layer_1[2638]; 
    assign out[2093] = layer_1[3927]; 
    assign out[2094] = ~(layer_1[394] ^ layer_1[425]); 
    assign out[2095] = layer_1[3793]; 
    assign out[2096] = layer_1[3414] | layer_1[3352]; 
    assign out[2097] = layer_1[3662] & ~layer_1[3536]; 
    assign out[2098] = ~layer_1[1828]; 
    assign out[2099] = ~layer_1[1141] | (layer_1[1141] & layer_1[1092]); 
    assign out[2100] = layer_1[3206] & ~layer_1[3205]; 
    assign out[2101] = ~(layer_1[2783] | layer_1[2817]); 
    assign out[2102] = layer_1[551] | layer_1[550]; 
    assign out[2103] = ~layer_1[1443] | (layer_1[1491] & layer_1[1443]); 
    assign out[2104] = ~(layer_1[3260] ^ layer_1[3350]); 
    assign out[2105] = layer_1[2518] ^ layer_1[2434]; 
    assign out[2106] = layer_1[1866] ^ layer_1[1962]; 
    assign out[2107] = ~(layer_1[1048] & layer_1[1027]); 
    assign out[2108] = ~layer_1[1877] | (layer_1[1877] & layer_1[1977]); 
    assign out[2109] = layer_1[2863] ^ layer_1[2919]; 
    assign out[2110] = ~layer_1[808]; 
    assign out[2111] = ~layer_1[169]; 
    assign out[2112] = ~layer_1[2745]; 
    assign out[2113] = ~layer_1[3599] | (layer_1[3599] & layer_1[3509]); 
    assign out[2114] = ~(layer_1[3962] ^ layer_1[3988]); 
    assign out[2115] = layer_1[2523] ^ layer_1[2444]; 
    assign out[2116] = layer_1[1994] | layer_1[2012]; 
    assign out[2117] = layer_1[3636]; 
    assign out[2118] = layer_1[3882] ^ layer_1[3970]; 
    assign out[2119] = layer_1[2994]; 
    assign out[2120] = layer_1[3969] | layer_1[3957]; 
    assign out[2121] = ~(layer_1[2864] ^ layer_1[2870]); 
    assign out[2122] = layer_1[1585] & ~layer_1[1569]; 
    assign out[2123] = ~layer_1[3174] | (layer_1[3174] & layer_1[3188]); 
    assign out[2124] = ~(layer_1[2513] ^ layer_1[2409]); 
    assign out[2125] = layer_1[1270] ^ layer_1[1147]; 
    assign out[2126] = layer_1[286] & layer_1[399]; 
    assign out[2127] = layer_1[1709] & ~layer_1[1758]; 
    assign out[2128] = ~(layer_1[594] ^ layer_1[627]); 
    assign out[2129] = ~layer_1[3403] | (layer_1[3389] & layer_1[3403]); 
    assign out[2130] = ~(layer_1[2416] ^ layer_1[2468]); 
    assign out[2131] = layer_1[3662] ^ layer_1[3651]; 
    assign out[2132] = layer_1[1200] ^ layer_1[1298]; 
    assign out[2133] = ~(layer_1[2312] | layer_1[2191]); 
    assign out[2134] = ~layer_1[2696]; 
    assign out[2135] = ~layer_1[1573]; 
    assign out[2136] = layer_1[984] & ~layer_1[1059]; 
    assign out[2137] = ~layer_1[2270] | (layer_1[2270] & layer_1[2149]); 
    assign out[2138] = layer_1[2823] ^ layer_1[2820]; 
    assign out[2139] = ~(layer_1[2468] ^ layer_1[2573]); 
    assign out[2140] = layer_1[2182] ^ layer_1[2115]; 
    assign out[2141] = layer_1[928] ^ layer_1[844]; 
    assign out[2142] = ~(layer_1[1421] ^ layer_1[1438]); 
    assign out[2143] = ~(layer_1[3907] ^ layer_1[3831]); 
    assign out[2144] = layer_1[505] | layer_1[493]; 
    assign out[2145] = layer_1[2349]; 
    assign out[2146] = ~(layer_1[452] ^ layer_1[446]); 
    assign out[2147] = layer_1[3681] | layer_1[3710]; 
    assign out[2148] = ~(layer_1[2698] ^ layer_1[2627]); 
    assign out[2149] = layer_1[3409] & ~layer_1[3490]; 
    assign out[2150] = layer_1[533] & layer_1[432]; 
    assign out[2151] = ~(layer_1[1318] ^ layer_1[1226]); 
    assign out[2152] = layer_1[655] | layer_1[584]; 
    assign out[2153] = ~layer_1[2293] | (layer_1[2325] & layer_1[2293]); 
    assign out[2154] = ~layer_1[2872]; 
    assign out[2155] = ~(layer_1[3177] ^ layer_1[3059]); 
    assign out[2156] = ~layer_1[3958]; 
    assign out[2157] = layer_1[3997]; 
    assign out[2158] = layer_1[1456] & ~layer_1[1459]; 
    assign out[2159] = layer_1[2209] ^ layer_1[2155]; 
    assign out[2160] = layer_1[119] & ~layer_1[223]; 
    assign out[2161] = ~(layer_1[913] ^ layer_1[824]); 
    assign out[2162] = layer_1[3476] ^ layer_1[3456]; 
    assign out[2163] = ~layer_1[3580]; 
    assign out[2164] = layer_1[2837] | layer_1[2720]; 
    assign out[2165] = ~layer_1[2939]; 
    assign out[2166] = layer_1[958] ^ layer_1[878]; 
    assign out[2167] = layer_1[3420]; 
    assign out[2168] = layer_1[1022]; 
    assign out[2169] = ~(layer_1[2775] ^ layer_1[2833]); 
    assign out[2170] = ~layer_1[1637]; 
    assign out[2171] = layer_1[3517] & layer_1[3562]; 
    assign out[2172] = layer_1[2480]; 
    assign out[2173] = layer_1[2724]; 
    assign out[2174] = ~layer_1[2583]; 
    assign out[2175] = ~layer_1[157] | (layer_1[157] & layer_1[73]); 
    assign out[2176] = layer_1[2986] ^ layer_1[3006]; 
    assign out[2177] = ~layer_1[2651]; 
    assign out[2178] = layer_1[3544]; 
    assign out[2179] = ~layer_1[1174]; 
    assign out[2180] = layer_1[1594] & ~layer_1[1628]; 
    assign out[2181] = layer_1[3090]; 
    assign out[2182] = ~layer_1[2762]; 
    assign out[2183] = ~layer_1[573] | (layer_1[573] & layer_1[631]); 
    assign out[2184] = ~layer_1[310]; 
    assign out[2185] = layer_1[3934] | layer_1[3927]; 
    assign out[2186] = ~layer_1[1115] | (layer_1[1168] & layer_1[1115]); 
    assign out[2187] = layer_1[2874] ^ layer_1[2953]; 
    assign out[2188] = layer_1[3239]; 
    assign out[2189] = ~(layer_1[1537] & layer_1[1650]); 
    assign out[2190] = layer_1[1567] ^ layer_1[1506]; 
    assign out[2191] = layer_1[591]; 
    assign out[2192] = ~(layer_1[3656] ^ layer_1[3695]); 
    assign out[2193] = ~(layer_1[3923] | layer_1[3802]); 
    assign out[2194] = ~layer_1[3580] | (layer_1[3524] & layer_1[3580]); 
    assign out[2195] = ~layer_1[2376]; 
    assign out[2196] = ~layer_1[659]; 
    assign out[2197] = layer_1[290] & layer_1[199]; 
    assign out[2198] = ~(layer_1[1048] ^ layer_1[1029]); 
    assign out[2199] = layer_1[801]; 
    assign out[2200] = ~layer_1[2780]; 
    assign out[2201] = layer_1[2462]; 
    assign out[2202] = layer_1[2484] | layer_1[2399]; 
    assign out[2203] = ~(layer_1[3928] & layer_1[3916]); 
    assign out[2204] = ~layer_1[1487]; 
    assign out[2205] = ~(layer_1[2066] | layer_1[2144]); 
    assign out[2206] = layer_1[2725]; 
    assign out[2207] = layer_1[1389] & ~layer_1[1376]; 
    assign out[2208] = ~layer_1[3327]; 
    assign out[2209] = layer_1[2553]; 
    assign out[2210] = layer_1[1821]; 
    assign out[2211] = ~layer_1[3691] | (layer_1[3636] & layer_1[3691]); 
    assign out[2212] = layer_1[1609] & ~layer_1[1500]; 
    assign out[2213] = layer_1[2728]; 
    assign out[2214] = ~(layer_1[2479] ^ layer_1[2413]); 
    assign out[2215] = ~(layer_1[1539] ^ layer_1[1468]); 
    assign out[2216] = ~(layer_1[1824] & layer_1[1832]); 
    assign out[2217] = layer_1[1749] ^ layer_1[1761]; 
    assign out[2218] = ~(layer_1[2863] & layer_1[2798]); 
    assign out[2219] = ~layer_1[1755]; 
    assign out[2220] = ~(layer_1[169] & layer_1[237]); 
    assign out[2221] = layer_1[1068]; 
    assign out[2222] = layer_1[2802] & ~layer_1[2721]; 
    assign out[2223] = layer_1[155] ^ layer_1[30]; 
    assign out[2224] = ~layer_1[2376]; 
    assign out[2225] = layer_1[874] ^ layer_1[925]; 
    assign out[2226] = ~layer_1[1442] | (layer_1[1442] & layer_1[1429]); 
    assign out[2227] = layer_1[219] ^ layer_1[207]; 
    assign out[2228] = ~layer_1[2921]; 
    assign out[2229] = ~layer_1[2521]; 
    assign out[2230] = ~(layer_1[279] ^ layer_1[391]); 
    assign out[2231] = layer_1[1414]; 
    assign out[2232] = ~layer_1[24] | (layer_1[24] & layer_1[18]); 
    assign out[2233] = layer_1[2859]; 
    assign out[2234] = layer_1[2118]; 
    assign out[2235] = layer_1[1374] ^ layer_1[1387]; 
    assign out[2236] = ~(layer_1[2555] ^ layer_1[2671]); 
    assign out[2237] = layer_1[621] ^ layer_1[692]; 
    assign out[2238] = ~layer_1[345]; 
    assign out[2239] = ~(layer_1[698] ^ layer_1[795]); 
    assign out[2240] = layer_1[3389] | layer_1[3339]; 
    assign out[2241] = layer_1[2882]; 
    assign out[2242] = layer_1[3748] & ~layer_1[3741]; 
    assign out[2243] = ~layer_1[1955]; 
    assign out[2244] = ~layer_1[1446]; 
    assign out[2245] = ~(layer_1[1925] & layer_1[1951]); 
    assign out[2246] = ~(layer_1[2271] ^ layer_1[2320]); 
    assign out[2247] = ~(layer_1[920] ^ layer_1[875]); 
    assign out[2248] = layer_1[1903] ^ layer_1[1991]; 
    assign out[2249] = ~(layer_1[3657] & layer_1[3612]); 
    assign out[2250] = layer_1[3421] ^ layer_1[3479]; 
    assign out[2251] = layer_1[1074]; 
    assign out[2252] = layer_1[167]; 
    assign out[2253] = ~layer_1[648]; 
    assign out[2254] = layer_1[210] & layer_1[294]; 
    assign out[2255] = ~(layer_1[2534] ^ layer_1[2541]); 
    assign out[2256] = ~layer_1[2814]; 
    assign out[2257] = layer_1[1137]; 
    assign out[2258] = layer_1[1296]; 
    assign out[2259] = layer_1[230]; 
    assign out[2260] = layer_1[2512] | layer_1[2456]; 
    assign out[2261] = layer_1[3604] & ~layer_1[3722]; 
    assign out[2262] = layer_1[3422]; 
    assign out[2263] = ~(layer_1[915] ^ layer_1[899]); 
    assign out[2264] = layer_1[3311]; 
    assign out[2265] = layer_1[608] ^ layer_1[651]; 
    assign out[2266] = ~(layer_1[941] | layer_1[962]); 
    assign out[2267] = layer_1[1074]; 
    assign out[2268] = layer_1[1161] ^ layer_1[1241]; 
    assign out[2269] = ~layer_1[1599]; 
    assign out[2270] = layer_1[639] & ~layer_1[699]; 
    assign out[2271] = layer_1[3815]; 
    assign out[2272] = layer_1[3389]; 
    assign out[2273] = ~layer_1[2015]; 
    assign out[2274] = layer_1[3856] ^ layer_1[3935]; 
    assign out[2275] = layer_1[622] ^ layer_1[561]; 
    assign out[2276] = layer_1[493]; 
    assign out[2277] = ~(layer_1[1133] & layer_1[1039]); 
    assign out[2278] = layer_1[1837]; 
    assign out[2279] = layer_1[3346]; 
    assign out[2280] = ~(layer_1[3110] & layer_1[3002]); 
    assign out[2281] = layer_1[1800] ^ layer_1[1814]; 
    assign out[2282] = ~layer_1[3472]; 
    assign out[2283] = ~layer_1[1833] | (layer_1[1833] & layer_1[1914]); 
    assign out[2284] = ~layer_1[968]; 
    assign out[2285] = ~layer_1[2308]; 
    assign out[2286] = ~(layer_1[3977] ^ layer_1[3874]); 
    assign out[2287] = ~(layer_1[2969] ^ layer_1[3006]); 
    assign out[2288] = ~(layer_1[1127] & layer_1[1095]); 
    assign out[2289] = ~layer_1[2467] | (layer_1[2362] & layer_1[2467]); 
    assign out[2290] = layer_1[2805] ^ layer_1[2850]; 
    assign out[2291] = ~(layer_1[561] | layer_1[573]); 
    assign out[2292] = layer_1[1182] & ~layer_1[1298]; 
    assign out[2293] = ~(layer_1[3395] ^ layer_1[3301]); 
    assign out[2294] = layer_1[2292] ^ layer_1[2261]; 
    assign out[2295] = layer_1[1753]; 
    assign out[2296] = ~layer_1[1412] | (layer_1[1412] & layer_1[1337]); 
    assign out[2297] = ~(layer_1[3497] | layer_1[3578]); 
    assign out[2298] = layer_1[670] ^ layer_1[576]; 
    assign out[2299] = ~layer_1[2125]; 
    assign out[2300] = ~(layer_1[1955] ^ layer_1[1879]); 
    assign out[2301] = ~(layer_1[3659] ^ layer_1[3623]); 
    assign out[2302] = ~layer_1[3226]; 
    assign out[2303] = layer_1[2142] | layer_1[2199]; 
    assign out[2304] = layer_1[1488] & ~layer_1[1380]; 
    assign out[2305] = layer_1[2162]; 
    assign out[2306] = ~(layer_1[3802] | layer_1[3734]); 
    assign out[2307] = layer_1[1635] ^ layer_1[1714]; 
    assign out[2308] = layer_1[3984]; 
    assign out[2309] = layer_1[1999] & ~layer_1[1986]; 
    assign out[2310] = layer_1[3682]; 
    assign out[2311] = ~(layer_1[857] ^ layer_1[850]); 
    assign out[2312] = layer_1[3064]; 
    assign out[2313] = layer_1[228] ^ layer_1[351]; 
    assign out[2314] = layer_1[466] & ~layer_1[561]; 
    assign out[2315] = ~(layer_1[953] & layer_1[1034]); 
    assign out[2316] = layer_1[2516] | layer_1[2514]; 
    assign out[2317] = layer_1[1540] & layer_1[1452]; 
    assign out[2318] = layer_1[3407] | layer_1[3477]; 
    assign out[2319] = layer_1[2025]; 
    assign out[2320] = layer_1[2040] ^ layer_1[2063]; 
    assign out[2321] = ~layer_1[100]; 
    assign out[2322] = layer_1[842]; 
    assign out[2323] = layer_1[2931] ^ layer_1[2839]; 
    assign out[2324] = layer_1[1425] & layer_1[1427]; 
    assign out[2325] = layer_1[482]; 
    assign out[2326] = layer_1[2207]; 
    assign out[2327] = layer_1[1151] & layer_1[1234]; 
    assign out[2328] = layer_1[101] & ~layer_1[71]; 
    assign out[2329] = layer_1[3685] ^ layer_1[3710]; 
    assign out[2330] = layer_1[1960] & ~layer_1[2034]; 
    assign out[2331] = layer_1[1710]; 
    assign out[2332] = ~layer_1[1617]; 
    assign out[2333] = layer_1[3306] | layer_1[3405]; 
    assign out[2334] = ~(layer_1[1778] ^ layer_1[1692]); 
    assign out[2335] = layer_1[2902]; 
    assign out[2336] = layer_1[3054]; 
    assign out[2337] = layer_1[1273] ^ layer_1[1313]; 
    assign out[2338] = layer_1[3041] & layer_1[3165]; 
    assign out[2339] = ~(layer_1[2472] ^ layer_1[2429]); 
    assign out[2340] = layer_1[1387] & ~layer_1[1334]; 
    assign out[2341] = ~layer_1[56]; 
    assign out[2342] = layer_1[1332] ^ layer_1[1363]; 
    assign out[2343] = ~(layer_1[377] ^ layer_1[322]); 
    assign out[2344] = ~layer_1[3606] | (layer_1[3517] & layer_1[3606]); 
    assign out[2345] = layer_1[1444] | layer_1[1572]; 
    assign out[2346] = ~layer_1[3883]; 
    assign out[2347] = ~layer_1[3057]; 
    assign out[2348] = layer_1[588] ^ layer_1[541]; 
    assign out[2349] = ~layer_1[487]; 
    assign out[2350] = ~layer_1[794]; 
    assign out[2351] = ~(layer_1[524] & layer_1[408]); 
    assign out[2352] = layer_1[2080]; 
    assign out[2353] = ~layer_1[1514]; 
    assign out[2354] = ~layer_1[3124] | (layer_1[3083] & layer_1[3124]); 
    assign out[2355] = ~layer_1[413] | (layer_1[406] & layer_1[413]); 
    assign out[2356] = ~layer_1[461] | (layer_1[402] & layer_1[461]); 
    assign out[2357] = ~(layer_1[3347] ^ layer_1[3437]); 
    assign out[2358] = layer_1[1082] ^ layer_1[1170]; 
    assign out[2359] = ~(layer_1[2339] ^ layer_1[2211]); 
    assign out[2360] = ~layer_1[204]; 
    assign out[2361] = layer_1[2223]; 
    assign out[2362] = ~(layer_1[1363] ^ layer_1[1433]); 
    assign out[2363] = layer_1[2217] & layer_1[2331]; 
    assign out[2364] = layer_1[3594] & layer_1[3538]; 
    assign out[2365] = ~(layer_1[1640] ^ layer_1[1734]); 
    assign out[2366] = layer_1[375] | layer_1[459]; 
    assign out[2367] = ~(layer_1[573] | layer_1[648]); 
    assign out[2368] = ~(layer_1[934] ^ layer_1[1014]); 
    assign out[2369] = layer_1[909]; 
    assign out[2370] = ~(layer_1[476] ^ layer_1[353]); 
    assign out[2371] = layer_1[1806]; 
    assign out[2372] = ~(layer_1[1997] & layer_1[2084]); 
    assign out[2373] = ~layer_1[1968] | (layer_1[1968] & layer_1[2010]); 
    assign out[2374] = layer_1[1540] & ~layer_1[1513]; 
    assign out[2375] = layer_1[2385]; 
    assign out[2376] = layer_1[106]; 
    assign out[2377] = layer_1[1486] ^ layer_1[1575]; 
    assign out[2378] = layer_1[2123]; 
    assign out[2379] = layer_1[3785]; 
    assign out[2380] = ~layer_1[1507] | (layer_1[1507] & layer_1[1633]); 
    assign out[2381] = layer_1[3020]; 
    assign out[2382] = layer_1[576]; 
    assign out[2383] = layer_1[1895] ^ layer_1[1954]; 
    assign out[2384] = layer_1[556] & ~layer_1[538]; 
    assign out[2385] = ~(layer_1[3959] ^ layer_1[3910]); 
    assign out[2386] = layer_1[114] ^ layer_1[82]; 
    assign out[2387] = ~layer_1[2195]; 
    assign out[2388] = layer_1[1779]; 
    assign out[2389] = layer_1[109]; 
    assign out[2390] = ~layer_1[968]; 
    assign out[2391] = layer_1[239] & ~layer_1[175]; 
    assign out[2392] = ~layer_1[3981]; 
    assign out[2393] = ~(layer_1[974] ^ layer_1[1076]); 
    assign out[2394] = layer_1[3481]; 
    assign out[2395] = layer_1[1166]; 
    assign out[2396] = layer_1[1144]; 
    assign out[2397] = ~layer_1[1081]; 
    assign out[2398] = layer_1[738] & ~layer_1[785]; 
    assign out[2399] = layer_1[1502] & ~layer_1[1513]; 
    assign out[2400] = layer_1[1777]; 
    assign out[2401] = ~layer_1[1959]; 
    assign out[2402] = layer_1[2099] & ~layer_1[2103]; 
    assign out[2403] = ~(layer_1[2937] ^ layer_1[2839]); 
    assign out[2404] = layer_1[1331] & ~layer_1[1227]; 
    assign out[2405] = ~(layer_1[2106] | layer_1[1990]); 
    assign out[2406] = layer_1[334] & ~layer_1[403]; 
    assign out[2407] = layer_1[1189] & ~layer_1[1102]; 
    assign out[2408] = ~(layer_1[2067] | layer_1[1972]); 
    assign out[2409] = layer_1[3949]; 
    assign out[2410] = ~layer_1[3364]; 
    assign out[2411] = ~(layer_1[1794] ^ layer_1[1686]); 
    assign out[2412] = ~(layer_1[1708] ^ layer_1[1726]); 
    assign out[2413] = layer_1[1929] & ~layer_1[1931]; 
    assign out[2414] = ~layer_1[2613]; 
    assign out[2415] = ~layer_1[2390]; 
    assign out[2416] = ~layer_1[2495]; 
    assign out[2417] = ~(layer_1[1554] | layer_1[1577]); 
    assign out[2418] = ~(layer_1[1103] ^ layer_1[975]); 
    assign out[2419] = layer_1[742] & ~layer_1[722]; 
    assign out[2420] = layer_1[2453]; 
    assign out[2421] = layer_1[2848] & ~layer_1[2851]; 
    assign out[2422] = ~(layer_1[2359] ^ layer_1[2266]); 
    assign out[2423] = layer_1[2292] & ~layer_1[2408]; 
    assign out[2424] = layer_1[2367]; 
    assign out[2425] = layer_1[3727]; 
    assign out[2426] = ~layer_1[1419] | (layer_1[1419] & layer_1[1447]); 
    assign out[2427] = ~layer_1[2224] | (layer_1[2300] & layer_1[2224]); 
    assign out[2428] = layer_1[1975] ^ layer_1[1888]; 
    assign out[2429] = ~layer_1[55]; 
    assign out[2430] = ~(layer_1[618] & layer_1[590]); 
    assign out[2431] = layer_1[3621]; 
    assign out[2432] = ~layer_1[1506]; 
    assign out[2433] = layer_1[1689]; 
    assign out[2434] = ~layer_1[2907]; 
    assign out[2435] = layer_1[429] & ~layer_1[306]; 
    assign out[2436] = ~layer_1[3060]; 
    assign out[2437] = ~(layer_1[2534] & layer_1[2501]); 
    assign out[2438] = layer_1[3488]; 
    assign out[2439] = layer_1[2333] ^ layer_1[2379]; 
    assign out[2440] = layer_1[1060] ^ layer_1[1085]; 
    assign out[2441] = layer_1[2584] & ~layer_1[2506]; 
    assign out[2442] = ~(layer_1[342] & layer_1[408]); 
    assign out[2443] = layer_1[2531]; 
    assign out[2444] = ~(layer_1[2590] | layer_1[2676]); 
    assign out[2445] = ~(layer_1[3122] & layer_1[3196]); 
    assign out[2446] = ~layer_1[1419] | (layer_1[1419] & layer_1[1400]); 
    assign out[2447] = layer_1[1397] | layer_1[1404]; 
    assign out[2448] = ~(layer_1[1361] ^ layer_1[1249]); 
    assign out[2449] = layer_1[1037] & ~layer_1[1151]; 
    assign out[2450] = ~layer_1[3935]; 
    assign out[2451] = layer_1[331] & ~layer_1[443]; 
    assign out[2452] = ~layer_1[1451]; 
    assign out[2453] = layer_1[1739] ^ layer_1[1645]; 
    assign out[2454] = layer_1[3951] & layer_1[3830]; 
    assign out[2455] = ~layer_1[765]; 
    assign out[2456] = layer_1[3396] ^ layer_1[3485]; 
    assign out[2457] = ~(layer_1[1364] | layer_1[1287]); 
    assign out[2458] = layer_1[3138]; 
    assign out[2459] = ~layer_1[923]; 
    assign out[2460] = ~layer_1[3762] | (layer_1[3846] & layer_1[3762]); 
    assign out[2461] = layer_1[2655] ^ layer_1[2650]; 
    assign out[2462] = layer_1[267]; 
    assign out[2463] = ~(layer_1[9] | layer_1[130]); 
    assign out[2464] = layer_1[137]; 
    assign out[2465] = ~(layer_1[2855] ^ layer_1[2829]); 
    assign out[2466] = ~(layer_1[2437] & layer_1[2401]); 
    assign out[2467] = layer_1[1885] & ~layer_1[1805]; 
    assign out[2468] = layer_1[1723] ^ layer_1[1655]; 
    assign out[2469] = layer_1[193] & layer_1[200]; 
    assign out[2470] = ~layer_1[2743]; 
    assign out[2471] = layer_1[3949]; 
    assign out[2472] = layer_1[207] & layer_1[190]; 
    assign out[2473] = layer_1[2335] & layer_1[2268]; 
    assign out[2474] = layer_1[1766] & ~layer_1[1881]; 
    assign out[2475] = layer_1[3009] | layer_1[2921]; 
    assign out[2476] = layer_1[2598] | layer_1[2569]; 
    assign out[2477] = layer_1[836] ^ layer_1[790]; 
    assign out[2478] = ~layer_1[2516]; 
    assign out[2479] = layer_1[1983] & ~layer_1[1943]; 
    assign out[2480] = ~layer_1[2992]; 
    assign out[2481] = layer_1[773] ^ layer_1[772]; 
    assign out[2482] = layer_1[1141] | layer_1[1039]; 
    assign out[2483] = ~(layer_1[176] ^ layer_1[99]); 
    assign out[2484] = layer_1[2176]; 
    assign out[2485] = ~layer_1[3348]; 
    assign out[2486] = ~(layer_1[2992] | layer_1[2909]); 
    assign out[2487] = ~(layer_1[3592] ^ layer_1[3691]); 
    assign out[2488] = layer_1[2422] & layer_1[2308]; 
    assign out[2489] = layer_1[1676]; 
    assign out[2490] = ~(layer_1[3104] & layer_1[3132]); 
    assign out[2491] = layer_1[1835]; 
    assign out[2492] = layer_1[3553]; 
    assign out[2493] = layer_1[3263] & ~layer_1[3365]; 
    assign out[2494] = ~(layer_1[1839] | layer_1[1812]); 
    assign out[2495] = ~(layer_1[1957] | layer_1[1979]); 
    assign out[2496] = ~(layer_1[384] ^ layer_1[325]); 
    assign out[2497] = ~layer_1[863]; 
    assign out[2498] = layer_1[3289] & ~layer_1[3329]; 
    assign out[2499] = layer_1[1536] & ~layer_1[1506]; 
    assign out[2500] = layer_1[566] ^ layer_1[673]; 
    assign out[2501] = ~(layer_1[214] ^ layer_1[170]); 
    assign out[2502] = layer_1[1303]; 
    assign out[2503] = layer_1[2723]; 
    assign out[2504] = ~layer_1[3081]; 
    assign out[2505] = ~layer_1[1496]; 
    assign out[2506] = layer_1[862] & ~layer_1[856]; 
    assign out[2507] = layer_1[2001]; 
    assign out[2508] = layer_1[2214] & ~layer_1[2220]; 
    assign out[2509] = ~layer_1[1639]; 
    assign out[2510] = ~(layer_1[2162] | layer_1[2131]); 
    assign out[2511] = ~layer_1[823]; 
    assign out[2512] = ~(layer_1[1726] ^ layer_1[1630]); 
    assign out[2513] = layer_1[3478] & ~layer_1[3474]; 
    assign out[2514] = layer_1[3634] & layer_1[3641]; 
    assign out[2515] = layer_1[6] & ~layer_1[125]; 
    assign out[2516] = layer_1[1870]; 
    assign out[2517] = layer_1[3533] & ~layer_1[3589]; 
    assign out[2518] = layer_1[670] & layer_1[600]; 
    assign out[2519] = layer_1[2915]; 
    assign out[2520] = ~layer_1[3231]; 
    assign out[2521] = ~(layer_1[91] | layer_1[131]); 
    assign out[2522] = layer_1[2079]; 
    assign out[2523] = layer_1[3469] ^ layer_1[3458]; 
    assign out[2524] = ~layer_1[1439]; 
    assign out[2525] = layer_1[165] ^ layer_1[214]; 
    assign out[2526] = layer_1[1369] & ~layer_1[1432]; 
    assign out[2527] = layer_1[3048] & layer_1[3156]; 
    assign out[2528] = layer_1[1153] & ~layer_1[1066]; 
    assign out[2529] = ~(layer_1[3600] & layer_1[3647]); 
    assign out[2530] = ~layer_1[3765]; 
    assign out[2531] = layer_1[1546] & layer_1[1592]; 
    assign out[2532] = layer_1[2911]; 
    assign out[2533] = ~(layer_1[1351] ^ layer_1[1367]); 
    assign out[2534] = layer_1[918] & layer_1[820]; 
    assign out[2535] = layer_1[999] & ~layer_1[1001]; 
    assign out[2536] = ~layer_1[1801]; 
    assign out[2537] = ~layer_1[3045]; 
    assign out[2538] = layer_1[3553]; 
    assign out[2539] = ~layer_1[3873] | (layer_1[3873] & layer_1[3850]); 
    assign out[2540] = ~layer_1[1745]; 
    assign out[2541] = ~(layer_1[1182] ^ layer_1[1225]); 
    assign out[2542] = ~(layer_1[672] | layer_1[775]); 
    assign out[2543] = layer_1[86] ^ layer_1[147]; 
    assign out[2544] = layer_1[3907] ^ layer_1[3894]; 
    assign out[2545] = layer_1[3276] ^ layer_1[3152]; 
    assign out[2546] = ~(layer_1[989] | layer_1[885]); 
    assign out[2547] = ~layer_1[2753] | (layer_1[2680] & layer_1[2753]); 
    assign out[2548] = layer_1[3466] & ~layer_1[3555]; 
    assign out[2549] = layer_1[1774]; 
    assign out[2550] = layer_1[1476]; 
    assign out[2551] = layer_1[3004] & layer_1[2898]; 
    assign out[2552] = ~layer_1[3932] | (layer_1[3943] & layer_1[3932]); 
    assign out[2553] = layer_1[2244]; 
    assign out[2554] = layer_1[3780] ^ layer_1[3859]; 
    assign out[2555] = layer_1[2794] & layer_1[2896]; 
    assign out[2556] = layer_1[1701] ^ layer_1[1649]; 
    assign out[2557] = layer_1[2459] & ~layer_1[2567]; 
    assign out[2558] = ~(layer_1[255] & layer_1[351]); 
    assign out[2559] = layer_1[3141]; 
    assign out[2560] = ~(layer_1[3833] ^ layer_1[3828]); 
    assign out[2561] = ~layer_1[305]; 
    assign out[2562] = layer_1[1760] & ~layer_1[1818]; 
    assign out[2563] = layer_1[3360]; 
    assign out[2564] = ~layer_1[1262]; 
    assign out[2565] = ~(layer_1[2109] | layer_1[2093]); 
    assign out[2566] = ~(layer_1[1427] ^ layer_1[1415]); 
    assign out[2567] = layer_1[908] & ~layer_1[803]; 
    assign out[2568] = layer_1[3192] ^ layer_1[3078]; 
    assign out[2569] = layer_1[2363]; 
    assign out[2570] = ~layer_1[2436] | (layer_1[2446] & layer_1[2436]); 
    assign out[2571] = ~(layer_1[819] & layer_1[843]); 
    assign out[2572] = layer_1[1881] ^ layer_1[1813]; 
    assign out[2573] = ~(layer_1[3813] ^ layer_1[3834]); 
    assign out[2574] = ~(layer_1[901] & layer_1[1005]); 
    assign out[2575] = ~(layer_1[1497] ^ layer_1[1418]); 
    assign out[2576] = layer_1[1148] & ~layer_1[1120]; 
    assign out[2577] = layer_1[1180] & ~layer_1[1227]; 
    assign out[2578] = layer_1[2204] & ~layer_1[2267]; 
    assign out[2579] = layer_1[2083] & ~layer_1[1974]; 
    assign out[2580] = layer_1[2712] & ~layer_1[2785]; 
    assign out[2581] = layer_1[904] & layer_1[818]; 
    assign out[2582] = layer_1[3800]; 
    assign out[2583] = layer_1[2987] | layer_1[2875]; 
    assign out[2584] = layer_1[1266]; 
    assign out[2585] = ~(layer_1[3879] | layer_1[3790]); 
    assign out[2586] = layer_1[2238] & layer_1[2168]; 
    assign out[2587] = ~layer_1[3154]; 
    assign out[2588] = layer_1[3603]; 
    assign out[2589] = layer_1[1132] & ~layer_1[1254]; 
    assign out[2590] = ~layer_1[302]; 
    assign out[2591] = layer_1[3269] & layer_1[3171]; 
    assign out[2592] = layer_1[3635] ^ layer_1[3705]; 
    assign out[2593] = ~layer_1[1379] | (layer_1[1374] & layer_1[1379]); 
    assign out[2594] = ~layer_1[3735] | (layer_1[3735] & layer_1[3703]); 
    assign out[2595] = ~(layer_1[3490] ^ layer_1[3469]); 
    assign out[2596] = ~(layer_1[3288] | layer_1[3356]); 
    assign out[2597] = ~(layer_1[3854] | layer_1[3742]); 
    assign out[2598] = ~(layer_1[1808] | layer_1[1717]); 
    assign out[2599] = layer_1[2690] | layer_1[2757]; 
    assign out[2600] = ~layer_1[1514]; 
    assign out[2601] = layer_1[3032]; 
    assign out[2602] = ~layer_1[1877]; 
    assign out[2603] = layer_1[644] & ~layer_1[609]; 
    assign out[2604] = ~(layer_1[2977] ^ layer_1[2854]); 
    assign out[2605] = ~(layer_1[2200] | layer_1[2126]); 
    assign out[2606] = ~(layer_1[1219] | layer_1[1214]); 
    assign out[2607] = ~layer_1[2288]; 
    assign out[2608] = ~(layer_1[175] ^ layer_1[199]); 
    assign out[2609] = layer_1[2105]; 
    assign out[2610] = ~layer_1[1999]; 
    assign out[2611] = layer_1[761] & ~layer_1[639]; 
    assign out[2612] = ~layer_1[916]; 
    assign out[2613] = ~(layer_1[3890] | layer_1[3991]); 
    assign out[2614] = layer_1[771]; 
    assign out[2615] = ~(layer_1[3711] & layer_1[3749]); 
    assign out[2616] = ~(layer_1[1162] ^ layer_1[1249]); 
    assign out[2617] = layer_1[231] | layer_1[332]; 
    assign out[2618] = layer_1[3516] & ~layer_1[3429]; 
    assign out[2619] = layer_1[1597] ^ layer_1[1606]; 
    assign out[2620] = ~layer_1[3211]; 
    assign out[2621] = layer_1[1966] & layer_1[1901]; 
    assign out[2622] = layer_1[3314] & layer_1[3389]; 
    assign out[2623] = ~layer_1[2358]; 
    assign out[2624] = layer_1[2086] ^ layer_1[2035]; 
    assign out[2625] = layer_1[631] & ~layer_1[530]; 
    assign out[2626] = layer_1[1150]; 
    assign out[2627] = layer_1[335] & ~layer_1[268]; 
    assign out[2628] = ~layer_1[3672]; 
    assign out[2629] = ~layer_1[1056]; 
    assign out[2630] = ~(layer_1[3486] ^ layer_1[3473]); 
    assign out[2631] = layer_1[3877] & ~layer_1[3928]; 
    assign out[2632] = ~(layer_1[264] & layer_1[305]); 
    assign out[2633] = ~layer_1[2154] | (layer_1[2154] & layer_1[2214]); 
    assign out[2634] = layer_1[1878] & ~layer_1[2006]; 
    assign out[2635] = ~(layer_1[26] | layer_1[93]); 
    assign out[2636] = layer_1[1814] & ~layer_1[1784]; 
    assign out[2637] = layer_1[3602] & layer_1[3581]; 
    assign out[2638] = layer_1[1778]; 
    assign out[2639] = ~layer_1[3538]; 
    assign out[2640] = layer_1[2937]; 
    assign out[2641] = ~layer_1[1419] | (layer_1[1419] & layer_1[1297]); 
    assign out[2642] = ~(layer_1[2142] | layer_1[2057]); 
    assign out[2643] = layer_1[449] & ~layer_1[525]; 
    assign out[2644] = layer_1[1892] ^ layer_1[2012]; 
    assign out[2645] = layer_1[365] & ~layer_1[477]; 
    assign out[2646] = layer_1[3220] | layer_1[3228]; 
    assign out[2647] = layer_1[1905]; 
    assign out[2648] = layer_1[3358]; 
    assign out[2649] = ~(layer_1[2595] & layer_1[2619]); 
    assign out[2650] = ~(layer_1[3087] ^ layer_1[3201]); 
    assign out[2651] = layer_1[1761] ^ layer_1[1855]; 
    assign out[2652] = ~layer_1[104]; 
    assign out[2653] = layer_1[2793]; 
    assign out[2654] = layer_1[3255] ^ layer_1[3242]; 
    assign out[2655] = ~(layer_1[1384] | layer_1[1466]); 
    assign out[2656] = ~layer_1[3960]; 
    assign out[2657] = layer_1[2210]; 
    assign out[2658] = layer_1[2738] & ~layer_1[2816]; 
    assign out[2659] = layer_1[2918] & layer_1[2828]; 
    assign out[2660] = layer_1[2894] ^ layer_1[2945]; 
    assign out[2661] = ~layer_1[2693]; 
    assign out[2662] = layer_1[3985] & ~layer_1[3993]; 
    assign out[2663] = ~layer_1[3020]; 
    assign out[2664] = layer_1[761]; 
    assign out[2665] = layer_1[2280]; 
    assign out[2666] = layer_1[3676] & layer_1[3635]; 
    assign out[2667] = layer_1[315] & layer_1[352]; 
    assign out[2668] = ~layer_1[460]; 
    assign out[2669] = ~(layer_1[2806] ^ layer_1[2903]); 
    assign out[2670] = layer_1[2898] & layer_1[2980]; 
    assign out[2671] = layer_1[917] & ~layer_1[885]; 
    assign out[2672] = ~layer_1[108]; 
    assign out[2673] = ~(layer_1[484] | layer_1[468]); 
    assign out[2674] = layer_1[2967] & layer_1[2949]; 
    assign out[2675] = ~(layer_1[3705] ^ layer_1[3776]); 
    assign out[2676] = layer_1[607]; 
    assign out[2677] = ~(layer_1[1124] ^ layer_1[1157]); 
    assign out[2678] = layer_1[874] & ~layer_1[929]; 
    assign out[2679] = ~(layer_1[3205] ^ layer_1[3304]); 
    assign out[2680] = ~(layer_1[1823] ^ layer_1[1768]); 
    assign out[2681] = ~(layer_1[2883] ^ layer_1[2817]); 
    assign out[2682] = layer_1[2152] & ~layer_1[2067]; 
    assign out[2683] = layer_1[768]; 
    assign out[2684] = layer_1[1163] & ~layer_1[1199]; 
    assign out[2685] = ~(layer_1[1149] & layer_1[1062]); 
    assign out[2686] = ~layer_1[1036]; 
    assign out[2687] = layer_1[326] | layer_1[210]; 
    assign out[2688] = layer_1[3209] & ~layer_1[3085]; 
    assign out[2689] = layer_1[3625] & layer_1[3513]; 
    assign out[2690] = layer_1[932]; 
    assign out[2691] = ~layer_1[901] | (layer_1[810] & layer_1[901]); 
    assign out[2692] = layer_1[1053] & ~layer_1[1124]; 
    assign out[2693] = ~(layer_1[898] | layer_1[929]); 
    assign out[2694] = layer_1[3298] & ~layer_1[3399]; 
    assign out[2695] = ~(layer_1[2325] ^ layer_1[2396]); 
    assign out[2696] = ~(layer_1[3638] | layer_1[3673]); 
    assign out[2697] = ~layer_1[2682]; 
    assign out[2698] = ~(layer_1[1803] ^ layer_1[1785]); 
    assign out[2699] = layer_1[675]; 
    assign out[2700] = layer_1[1537]; 
    assign out[2701] = ~layer_1[785]; 
    assign out[2702] = layer_1[2314]; 
    assign out[2703] = ~layer_1[1718]; 
    assign out[2704] = ~(layer_1[3778] & layer_1[3769]); 
    assign out[2705] = ~layer_1[1451]; 
    assign out[2706] = layer_1[2719] & ~layer_1[2668]; 
    assign out[2707] = ~(layer_1[3075] & layer_1[3167]); 
    assign out[2708] = layer_1[2373] | layer_1[2301]; 
    assign out[2709] = layer_1[3006] & ~layer_1[2883]; 
    assign out[2710] = ~(layer_1[572] | layer_1[490]); 
    assign out[2711] = layer_1[320]; 
    assign out[2712] = ~(layer_1[1765] | layer_1[1750]); 
    assign out[2713] = layer_1[659] & ~layer_1[566]; 
    assign out[2714] = layer_1[3705] ^ layer_1[3631]; 
    assign out[2715] = layer_1[3016]; 
    assign out[2716] = ~layer_1[1598]; 
    assign out[2717] = ~(layer_1[2345] ^ layer_1[2234]); 
    assign out[2718] = layer_1[1096]; 
    assign out[2719] = ~layer_1[1936]; 
    assign out[2720] = layer_1[2232] | layer_1[2245]; 
    assign out[2721] = layer_1[3764] ^ layer_1[3636]; 
    assign out[2722] = layer_1[694] ^ layer_1[795]; 
    assign out[2723] = layer_1[3646] | layer_1[3681]; 
    assign out[2724] = layer_1[2560]; 
    assign out[2725] = ~layer_1[3626]; 
    assign out[2726] = ~layer_1[3261] | (layer_1[3261] & layer_1[3263]); 
    assign out[2727] = layer_1[845]; 
    assign out[2728] = ~layer_1[1064] | (layer_1[1166] & layer_1[1064]); 
    assign out[2729] = ~layer_1[3474]; 
    assign out[2730] = ~layer_1[3956]; 
    assign out[2731] = layer_1[1580]; 
    assign out[2732] = ~layer_1[1633]; 
    assign out[2733] = ~layer_1[3355]; 
    assign out[2734] = layer_1[2110] & ~layer_1[2068]; 
    assign out[2735] = layer_1[2094] ^ layer_1[2096]; 
    assign out[2736] = layer_1[1550]; 
    assign out[2737] = layer_1[267] & ~layer_1[201]; 
    assign out[2738] = ~(layer_1[3745] | layer_1[3697]); 
    assign out[2739] = ~(layer_1[1999] & layer_1[2113]); 
    assign out[2740] = ~(layer_1[3252] ^ layer_1[3325]); 
    assign out[2741] = ~layer_1[901] | (layer_1[901] & layer_1[966]); 
    assign out[2742] = layer_1[243]; 
    assign out[2743] = ~(layer_1[2878] | layer_1[2978]); 
    assign out[2744] = ~layer_1[197]; 
    assign out[2745] = ~(layer_1[3652] ^ layer_1[3619]); 
    assign out[2746] = layer_1[2351]; 
    assign out[2747] = layer_1[1695] | layer_1[1822]; 
    assign out[2748] = ~layer_1[1891]; 
    assign out[2749] = layer_1[1607] ^ layer_1[1563]; 
    assign out[2750] = ~layer_1[1808]; 
    assign out[2751] = ~layer_1[2668]; 
    assign out[2752] = ~(layer_1[1957] ^ layer_1[1919]); 
    assign out[2753] = layer_1[3073] | layer_1[3148]; 
    assign out[2754] = ~layer_1[2822]; 
    assign out[2755] = layer_1[712]; 
    assign out[2756] = layer_1[986] & ~layer_1[1001]; 
    assign out[2757] = layer_1[2018] ^ layer_1[2135]; 
    assign out[2758] = ~layer_1[658] | (layer_1[716] & layer_1[658]); 
    assign out[2759] = ~layer_1[554]; 
    assign out[2760] = layer_1[2673] ^ layer_1[2705]; 
    assign out[2761] = layer_1[2807] & layer_1[2694]; 
    assign out[2762] = layer_1[2238] & ~layer_1[2321]; 
    assign out[2763] = ~(layer_1[2798] | layer_1[2804]); 
    assign out[2764] = ~(layer_1[3051] ^ layer_1[2970]); 
    assign out[2765] = layer_1[2618] ^ layer_1[2523]; 
    assign out[2766] = layer_1[3886] & layer_1[3997]; 
    assign out[2767] = layer_1[833] & ~layer_1[936]; 
    assign out[2768] = ~layer_1[422]; 
    assign out[2769] = ~(layer_1[1784] ^ layer_1[1731]); 
    assign out[2770] = ~(layer_1[503] ^ layer_1[430]); 
    assign out[2771] = ~layer_1[2622]; 
    assign out[2772] = layer_1[917] & layer_1[857]; 
    assign out[2773] = ~(layer_1[2161] ^ layer_1[2199]); 
    assign out[2774] = layer_1[1271] & layer_1[1300]; 
    assign out[2775] = ~layer_1[2103]; 
    assign out[2776] = layer_1[3000] | layer_1[3004]; 
    assign out[2777] = ~layer_1[3050]; 
    assign out[2778] = ~layer_1[3892]; 
    assign out[2779] = layer_1[377] & ~layer_1[252]; 
    assign out[2780] = ~(layer_1[1394] | layer_1[1494]); 
    assign out[2781] = layer_1[281]; 
    assign out[2782] = ~(layer_1[3552] ^ layer_1[3534]); 
    assign out[2783] = ~(layer_1[2822] ^ layer_1[2922]); 
    assign out[2784] = layer_1[146] & layer_1[160]; 
    assign out[2785] = layer_1[1294] | layer_1[1290]; 
    assign out[2786] = layer_1[1602]; 
    assign out[2787] = layer_1[562] | layer_1[666]; 
    assign out[2788] = ~(layer_1[2498] | layer_1[2565]); 
    assign out[2789] = layer_1[1377]; 
    assign out[2790] = layer_1[2363]; 
    assign out[2791] = layer_1[1376] & ~layer_1[1465]; 
    assign out[2792] = ~(layer_1[777] ^ layer_1[695]); 
    assign out[2793] = ~(layer_1[2002] | layer_1[1893]); 
    assign out[2794] = layer_1[3955] & ~layer_1[3944]; 
    assign out[2795] = ~(layer_1[839] ^ layer_1[810]); 
    assign out[2796] = layer_1[1531]; 
    assign out[2797] = ~layer_1[1824]; 
    assign out[2798] = ~layer_1[3394] | (layer_1[3394] & layer_1[3280]); 
    assign out[2799] = layer_1[2973] ^ layer_1[2887]; 
    assign out[2800] = ~layer_1[321] | (layer_1[321] & layer_1[277]); 
    assign out[2801] = layer_1[1939] & layer_1[1951]; 
    assign out[2802] = layer_1[3600] | layer_1[3507]; 
    assign out[2803] = layer_1[1128]; 
    assign out[2804] = ~layer_1[220]; 
    assign out[2805] = layer_1[3174]; 
    assign out[2806] = layer_1[2000]; 
    assign out[2807] = layer_1[792] ^ layer_1[735]; 
    assign out[2808] = layer_1[1682] | layer_1[1670]; 
    assign out[2809] = ~layer_1[2544]; 
    assign out[2810] = ~(layer_1[3345] ^ layer_1[3242]); 
    assign out[2811] = ~(layer_1[3054] & layer_1[3015]); 
    assign out[2812] = layer_1[931] & layer_1[971]; 
    assign out[2813] = ~layer_1[990]; 
    assign out[2814] = ~layer_1[2074] | (layer_1[2074] & layer_1[2050]); 
    assign out[2815] = layer_1[3383]; 
    assign out[2816] = ~(layer_1[35] & layer_1[42]); 
    assign out[2817] = ~(layer_1[1706] & layer_1[1692]); 
    assign out[2818] = layer_1[3205] & ~layer_1[3291]; 
    assign out[2819] = ~(layer_1[804] | layer_1[921]); 
    assign out[2820] = ~(layer_1[1284] ^ layer_1[1360]); 
    assign out[2821] = layer_1[3432] & layer_1[3487]; 
    assign out[2822] = ~(layer_1[3211] ^ layer_1[3272]); 
    assign out[2823] = layer_1[3670]; 
    assign out[2824] = layer_1[846] ^ layer_1[957]; 
    assign out[2825] = layer_1[1867] & layer_1[1769]; 
    assign out[2826] = ~(layer_1[1845] ^ layer_1[1837]); 
    assign out[2827] = layer_1[1007] | layer_1[1025]; 
    assign out[2828] = layer_1[3769] | layer_1[3849]; 
    assign out[2829] = layer_1[1687]; 
    assign out[2830] = ~(layer_1[560] ^ layer_1[540]); 
    assign out[2831] = ~(layer_1[3422] ^ layer_1[3375]); 
    assign out[2832] = layer_1[1194] ^ layer_1[1305]; 
    assign out[2833] = ~layer_1[352]; 
    assign out[2834] = layer_1[2682] ^ layer_1[2554]; 
    assign out[2835] = ~(layer_1[3048] ^ layer_1[3097]); 
    assign out[2836] = ~layer_1[368]; 
    assign out[2837] = layer_1[1063] ^ layer_1[1014]; 
    assign out[2838] = ~(layer_1[3072] ^ layer_1[2963]); 
    assign out[2839] = ~(layer_1[3696] ^ layer_1[3785]); 
    assign out[2840] = layer_1[3336]; 
    assign out[2841] = ~layer_1[2660]; 
    assign out[2842] = ~(layer_1[791] ^ layer_1[723]); 
    assign out[2843] = layer_1[1313]; 
    assign out[2844] = layer_1[1171]; 
    assign out[2845] = layer_1[937] ^ layer_1[932]; 
    assign out[2846] = layer_1[1617] & layer_1[1592]; 
    assign out[2847] = ~layer_1[379]; 
    assign out[2848] = layer_1[3916] ^ layer_1[3930]; 
    assign out[2849] = layer_1[2443] & ~layer_1[2350]; 
    assign out[2850] = layer_1[1867]; 
    assign out[2851] = layer_1[513] | layer_1[394]; 
    assign out[2852] = ~layer_1[1819] | (layer_1[1750] & layer_1[1819]); 
    assign out[2853] = ~(layer_1[119] | layer_1[76]); 
    assign out[2854] = ~(layer_1[450] ^ layer_1[382]); 
    assign out[2855] = layer_1[2366]; 
    assign out[2856] = ~layer_1[3311] | (layer_1[3401] & layer_1[3311]); 
    assign out[2857] = layer_1[1254]; 
    assign out[2858] = layer_1[3756] ^ layer_1[3750]; 
    assign out[2859] = ~(layer_1[2045] | layer_1[1969]); 
    assign out[2860] = ~(layer_1[1624] | layer_1[1579]); 
    assign out[2861] = ~layer_1[3944]; 
    assign out[2862] = layer_1[2872] & layer_1[2966]; 
    assign out[2863] = layer_1[539] & ~layer_1[580]; 
    assign out[2864] = ~layer_1[3595]; 
    assign out[2865] = ~layer_1[3649]; 
    assign out[2866] = layer_1[546]; 
    assign out[2867] = ~layer_1[3553]; 
    assign out[2868] = ~layer_1[1847]; 
    assign out[2869] = ~(layer_1[3711] ^ layer_1[3692]); 
    assign out[2870] = ~layer_1[266]; 
    assign out[2871] = layer_1[93]; 
    assign out[2872] = layer_1[2059]; 
    assign out[2873] = ~(layer_1[352] | layer_1[321]); 
    assign out[2874] = layer_1[755]; 
    assign out[2875] = layer_1[285] | layer_1[224]; 
    assign out[2876] = ~layer_1[3925]; 
    assign out[2877] = ~(layer_1[2393] ^ layer_1[2429]); 
    assign out[2878] = layer_1[255] & layer_1[225]; 
    assign out[2879] = ~layer_1[3569]; 
    assign out[2880] = layer_1[636]; 
    assign out[2881] = layer_1[3886] ^ layer_1[3777]; 
    assign out[2882] = ~layer_1[251]; 
    assign out[2883] = ~(layer_1[3566] ^ layer_1[3571]); 
    assign out[2884] = layer_1[1641] & layer_1[1601]; 
    assign out[2885] = layer_1[2490] ^ layer_1[2564]; 
    assign out[2886] = layer_1[2753] & ~layer_1[2654]; 
    assign out[2887] = layer_1[152]; 
    assign out[2888] = layer_1[546]; 
    assign out[2889] = layer_1[2066] | layer_1[2181]; 
    assign out[2890] = ~layer_1[2630]; 
    assign out[2891] = layer_1[2664] ^ layer_1[2633]; 
    assign out[2892] = layer_1[689]; 
    assign out[2893] = ~layer_1[3521]; 
    assign out[2894] = ~(layer_1[452] | layer_1[424]); 
    assign out[2895] = ~(layer_1[1166] | layer_1[1087]); 
    assign out[2896] = ~layer_1[3546]; 
    assign out[2897] = ~layer_1[422] | (layer_1[413] & layer_1[422]); 
    assign out[2898] = layer_1[312] & ~layer_1[370]; 
    assign out[2899] = ~(layer_1[2370] ^ layer_1[2414]); 
    assign out[2900] = layer_1[3027]; 
    assign out[2901] = layer_1[3086]; 
    assign out[2902] = ~(layer_1[2815] | layer_1[2921]); 
    assign out[2903] = layer_1[1114]; 
    assign out[2904] = layer_1[3316]; 
    assign out[2905] = ~layer_1[2353]; 
    assign out[2906] = layer_1[2144] & ~layer_1[2135]; 
    assign out[2907] = ~layer_1[3435]; 
    assign out[2908] = layer_1[862]; 
    assign out[2909] = layer_1[1769] & ~layer_1[1817]; 
    assign out[2910] = layer_1[3566] | layer_1[3613]; 
    assign out[2911] = layer_1[2308] ^ layer_1[2370]; 
    assign out[2912] = ~(layer_1[1268] ^ layer_1[1153]); 
    assign out[2913] = layer_1[3589] & ~layer_1[3520]; 
    assign out[2914] = layer_1[1895] & ~layer_1[1835]; 
    assign out[2915] = ~(layer_1[2940] | layer_1[2854]); 
    assign out[2916] = ~layer_1[2755]; 
    assign out[2917] = ~layer_1[2632]; 
    assign out[2918] = layer_1[3741] & ~layer_1[3695]; 
    assign out[2919] = ~(layer_1[111] & layer_1[222]); 
    assign out[2920] = ~layer_1[2572]; 
    assign out[2921] = layer_1[2700]; 
    assign out[2922] = layer_1[122] & layer_1[38]; 
    assign out[2923] = layer_1[897] ^ layer_1[832]; 
    assign out[2924] = ~(layer_1[3191] ^ layer_1[3225]); 
    assign out[2925] = ~layer_1[2415]; 
    assign out[2926] = ~layer_1[806] | (layer_1[695] & layer_1[806]); 
    assign out[2927] = layer_1[3589] | layer_1[3636]; 
    assign out[2928] = ~(layer_1[1965] ^ layer_1[2045]); 
    assign out[2929] = layer_1[147] | layer_1[200]; 
    assign out[2930] = layer_1[897] ^ layer_1[864]; 
    assign out[2931] = layer_1[1302] ^ layer_1[1284]; 
    assign out[2932] = ~layer_1[2374] | (layer_1[2354] & layer_1[2374]); 
    assign out[2933] = layer_1[319] & ~layer_1[395]; 
    assign out[2934] = ~(layer_1[872] ^ layer_1[891]); 
    assign out[2935] = ~(layer_1[429] & layer_1[548]); 
    assign out[2936] = layer_1[1648] & ~layer_1[1610]; 
    assign out[2937] = ~layer_1[1124]; 
    assign out[2938] = layer_1[2778] & ~layer_1[2688]; 
    assign out[2939] = ~layer_1[2533]; 
    assign out[2940] = ~layer_1[2255]; 
    assign out[2941] = layer_1[1101]; 
    assign out[2942] = layer_1[206]; 
    assign out[2943] = layer_1[827] & layer_1[714]; 
    assign out[2944] = layer_1[3784] ^ layer_1[3832]; 
    assign out[2945] = ~(layer_1[2933] ^ layer_1[3043]); 
    assign out[2946] = layer_1[3028]; 
    assign out[2947] = layer_1[644]; 
    assign out[2948] = ~(layer_1[3776] ^ layer_1[3802]); 
    assign out[2949] = ~layer_1[3857]; 
    assign out[2950] = ~layer_1[3569]; 
    assign out[2951] = layer_1[709]; 
    assign out[2952] = ~(layer_1[3158] ^ layer_1[3064]); 
    assign out[2953] = ~(layer_1[1375] ^ layer_1[1253]); 
    assign out[2954] = ~(layer_1[132] ^ layer_1[175]); 
    assign out[2955] = layer_1[2615] | layer_1[2539]; 
    assign out[2956] = layer_1[3741] | layer_1[3761]; 
    assign out[2957] = ~(layer_1[382] | layer_1[314]); 
    assign out[2958] = layer_1[3752]; 
    assign out[2959] = ~layer_1[1503]; 
    assign out[2960] = ~(layer_1[3998] ^ layer_1[3938]); 
    assign out[2961] = ~layer_1[248]; 
    assign out[2962] = layer_1[2736] | layer_1[2695]; 
    assign out[2963] = layer_1[32]; 
    assign out[2964] = layer_1[2482]; 
    assign out[2965] = layer_1[2220] ^ layer_1[2342]; 
    assign out[2966] = layer_1[2099] | layer_1[2013]; 
    assign out[2967] = layer_1[618] & ~layer_1[688]; 
    assign out[2968] = layer_1[2007]; 
    assign out[2969] = ~(layer_1[984] ^ layer_1[1008]); 
    assign out[2970] = layer_1[2372] ^ layer_1[2361]; 
    assign out[2971] = ~(layer_1[1047] ^ layer_1[954]); 
    assign out[2972] = layer_1[1577] | layer_1[1620]; 
    assign out[2973] = ~layer_1[672] | (layer_1[697] & layer_1[672]); 
    assign out[2974] = layer_1[3713]; 
    assign out[2975] = ~(layer_1[1676] | layer_1[1643]); 
    assign out[2976] = ~(layer_1[3386] & layer_1[3273]); 
    assign out[2977] = ~(layer_1[657] ^ layer_1[651]); 
    assign out[2978] = layer_1[3628]; 
    assign out[2979] = layer_1[3434] | layer_1[3507]; 
    assign out[2980] = ~(layer_1[2207] & layer_1[2100]); 
    assign out[2981] = ~(layer_1[2312] & layer_1[2197]); 
    assign out[2982] = layer_1[1571] & layer_1[1622]; 
    assign out[2983] = ~layer_1[3933] | (layer_1[3933] & layer_1[3915]); 
    assign out[2984] = layer_1[2910] | layer_1[2917]; 
    assign out[2985] = ~layer_1[2520]; 
    assign out[2986] = ~layer_1[745]; 
    assign out[2987] = layer_1[868] ^ layer_1[987]; 
    assign out[2988] = layer_1[1959] & ~layer_1[1956]; 
    assign out[2989] = ~(layer_1[1452] ^ layer_1[1457]); 
    assign out[2990] = layer_1[1657]; 
    assign out[2991] = layer_1[951]; 
    assign out[2992] = layer_1[3110] & ~layer_1[3165]; 
    assign out[2993] = ~(layer_1[2680] & layer_1[2747]); 
    assign out[2994] = ~layer_1[2519]; 
    assign out[2995] = ~layer_1[3363]; 
    assign out[2996] = layer_1[2054]; 
    assign out[2997] = ~layer_1[2979]; 
    assign out[2998] = layer_1[3961]; 
    assign out[2999] = ~layer_1[3222] | (layer_1[3222] & layer_1[3098]); 
    assign out[3000] = layer_1[1675]; 
    assign out[3001] = layer_1[2866]; 
    assign out[3002] = ~layer_1[849] | (layer_1[971] & layer_1[849]); 
    assign out[3003] = layer_1[1789] & layer_1[1715]; 
    assign out[3004] = ~layer_1[462]; 
    assign out[3005] = layer_1[2058] & ~layer_1[1952]; 
    assign out[3006] = layer_1[878] & ~layer_1[840]; 
    assign out[3007] = ~layer_1[1387]; 
    assign out[3008] = ~layer_1[1357]; 
    assign out[3009] = layer_1[152] & ~layer_1[252]; 
    assign out[3010] = ~layer_1[142] | (layer_1[142] & layer_1[177]); 
    assign out[3011] = layer_1[2015] & ~layer_1[1934]; 
    assign out[3012] = ~layer_1[1096]; 
    assign out[3013] = ~(layer_1[2887] ^ layer_1[2765]); 
    assign out[3014] = ~layer_1[3727] | (layer_1[3606] & layer_1[3727]); 
    assign out[3015] = layer_1[1232]; 
    assign out[3016] = layer_1[3393]; 
    assign out[3017] = ~layer_1[154]; 
    assign out[3018] = layer_1[259]; 
    assign out[3019] = ~layer_1[324] | (layer_1[274] & layer_1[324]); 
    assign out[3020] = layer_1[1151] ^ layer_1[1099]; 
    assign out[3021] = ~(layer_1[57] ^ layer_1[162]); 
    assign out[3022] = ~layer_1[251]; 
    assign out[3023] = ~layer_1[3120] | (layer_1[3120] & layer_1[3039]); 
    assign out[3024] = ~layer_1[1354]; 
    assign out[3025] = layer_1[523]; 
    assign out[3026] = layer_1[2716]; 
    assign out[3027] = ~(layer_1[2342] ^ layer_1[2250]); 
    assign out[3028] = layer_1[3346]; 
    assign out[3029] = layer_1[2124] | layer_1[2211]; 
    assign out[3030] = ~layer_1[1542]; 
    assign out[3031] = layer_1[2984]; 
    assign out[3032] = layer_1[2811]; 
    assign out[3033] = layer_1[3349]; 
    assign out[3034] = ~layer_1[1118]; 
    assign out[3035] = ~layer_1[904]; 
    assign out[3036] = ~(layer_1[2316] | layer_1[2369]); 
    assign out[3037] = ~layer_1[1018]; 
    assign out[3038] = layer_1[1899] & layer_1[1920]; 
    assign out[3039] = ~layer_1[854]; 
    assign out[3040] = ~(layer_1[2121] & layer_1[2125]); 
    assign out[3041] = layer_1[3846] & ~layer_1[3828]; 
    assign out[3042] = ~layer_1[1297]; 
    assign out[3043] = layer_1[1367]; 
    assign out[3044] = ~layer_1[1038] | (layer_1[1038] & layer_1[992]); 
    assign out[3045] = ~layer_1[2594]; 
    assign out[3046] = ~layer_1[1286]; 
    assign out[3047] = layer_1[940] & ~layer_1[889]; 
    assign out[3048] = ~(layer_1[209] | layer_1[133]); 
    assign out[3049] = layer_1[3214] & ~layer_1[3209]; 
    assign out[3050] = layer_1[2036] & ~layer_1[1952]; 
    assign out[3051] = ~(layer_1[1330] | layer_1[1433]); 
    assign out[3052] = layer_1[3424]; 
    assign out[3053] = ~(layer_1[3865] | layer_1[3884]); 
    assign out[3054] = ~(layer_1[1227] ^ layer_1[1103]); 
    assign out[3055] = ~layer_1[334]; 
    assign out[3056] = ~(layer_1[3033] | layer_1[2933]); 
    assign out[3057] = layer_1[2611] ^ layer_1[2600]; 
    assign out[3058] = layer_1[2159]; 
    assign out[3059] = layer_1[144] & ~layer_1[183]; 
    assign out[3060] = layer_1[192] & ~layer_1[237]; 
    assign out[3061] = ~layer_1[1990]; 
    assign out[3062] = layer_1[2169] & ~layer_1[2069]; 
    assign out[3063] = layer_1[371] & ~layer_1[425]; 
    assign out[3064] = layer_1[953] & layer_1[871]; 
    assign out[3065] = ~(layer_1[429] & layer_1[462]); 
    assign out[3066] = ~layer_1[253]; 
    assign out[3067] = layer_1[775] ^ layer_1[834]; 
    assign out[3068] = ~layer_1[460] | (layer_1[387] & layer_1[460]); 
    assign out[3069] = layer_1[1060] & ~layer_1[1088]; 
    assign out[3070] = layer_1[1765]; 
    assign out[3071] = ~layer_1[1164] | (layer_1[1164] & layer_1[1273]); 
    assign out[3072] = layer_1[3128] & layer_1[3194]; 
    assign out[3073] = ~layer_1[3865]; 
    assign out[3074] = layer_1[262] | layer_1[316]; 
    assign out[3075] = ~layer_1[2173]; 
    assign out[3076] = ~(layer_1[2017] ^ layer_1[2014]); 
    assign out[3077] = ~(layer_1[1734] ^ layer_1[1804]); 
    assign out[3078] = layer_1[2513] & layer_1[2474]; 
    assign out[3079] = ~layer_1[739]; 
    assign out[3080] = layer_1[576]; 
    assign out[3081] = layer_1[1042]; 
    assign out[3082] = layer_1[2421] ^ layer_1[2388]; 
    assign out[3083] = layer_1[541] ^ layer_1[455]; 
    assign out[3084] = ~(layer_1[2757] | layer_1[2660]); 
    assign out[3085] = ~layer_1[3564]; 
    assign out[3086] = ~layer_1[570]; 
    assign out[3087] = layer_1[99] ^ layer_1[3]; 
    assign out[3088] = layer_1[548] ^ layer_1[665]; 
    assign out[3089] = ~(layer_1[1723] | layer_1[1829]); 
    assign out[3090] = layer_1[1890] & layer_1[1765]; 
    assign out[3091] = layer_1[2832] ^ layer_1[2756]; 
    assign out[3092] = ~layer_1[75]; 
    assign out[3093] = layer_1[1648]; 
    assign out[3094] = ~layer_1[3678]; 
    assign out[3095] = layer_1[933]; 
    assign out[3096] = ~layer_1[299]; 
    assign out[3097] = layer_1[2771]; 
    assign out[3098] = ~layer_1[1138] | (layer_1[1138] & layer_1[1201]); 
    assign out[3099] = layer_1[380]; 
    assign out[3100] = ~layer_1[3852]; 
    assign out[3101] = ~layer_1[3857]; 
    assign out[3102] = layer_1[3370]; 
    assign out[3103] = ~(layer_1[3928] ^ layer_1[3940]); 
    assign out[3104] = ~layer_1[1950]; 
    assign out[3105] = ~layer_1[472]; 
    assign out[3106] = layer_1[2496] & ~layer_1[2439]; 
    assign out[3107] = layer_1[1802] ^ layer_1[1846]; 
    assign out[3108] = ~layer_1[1538] | (layer_1[1620] & layer_1[1538]); 
    assign out[3109] = ~layer_1[2704] | (layer_1[2704] & layer_1[2790]); 
    assign out[3110] = layer_1[289] ^ layer_1[347]; 
    assign out[3111] = ~(layer_1[2012] | layer_1[2017]); 
    assign out[3112] = layer_1[1592] & ~layer_1[1707]; 
    assign out[3113] = layer_1[1218] & ~layer_1[1272]; 
    assign out[3114] = ~(layer_1[1517] | layer_1[1562]); 
    assign out[3115] = ~layer_1[467]; 
    assign out[3116] = ~layer_1[1960] | (layer_1[1960] & layer_1[2066]); 
    assign out[3117] = ~layer_1[679] | (layer_1[679] & layer_1[701]); 
    assign out[3118] = layer_1[1282] ^ layer_1[1227]; 
    assign out[3119] = ~layer_1[350]; 
    assign out[3120] = layer_1[580] ^ layer_1[674]; 
    assign out[3121] = ~(layer_1[2595] ^ layer_1[2675]); 
    assign out[3122] = layer_1[2592] & layer_1[2511]; 
    assign out[3123] = layer_1[3157] ^ layer_1[3266]; 
    assign out[3124] = ~layer_1[1458] | (layer_1[1458] & layer_1[1439]); 
    assign out[3125] = ~(layer_1[1926] ^ layer_1[1962]); 
    assign out[3126] = layer_1[2198] | layer_1[2302]; 
    assign out[3127] = layer_1[755]; 
    assign out[3128] = ~(layer_1[3897] ^ layer_1[3975]); 
    assign out[3129] = ~(layer_1[8] | layer_1[132]); 
    assign out[3130] = layer_1[2960]; 
    assign out[3131] = layer_1[2248]; 
    assign out[3132] = ~(layer_1[1782] | layer_1[1829]); 
    assign out[3133] = layer_1[1566]; 
    assign out[3134] = ~layer_1[1116]; 
    assign out[3135] = ~layer_1[3754]; 
    assign out[3136] = layer_1[1238] & ~layer_1[1139]; 
    assign out[3137] = layer_1[1729] ^ layer_1[1767]; 
    assign out[3138] = ~layer_1[2309]; 
    assign out[3139] = ~layer_1[2019] | (layer_1[2019] & layer_1[1968]); 
    assign out[3140] = layer_1[3077] & ~layer_1[2954]; 
    assign out[3141] = ~layer_1[2453]; 
    assign out[3142] = layer_1[2201] ^ layer_1[2077]; 
    assign out[3143] = layer_1[1402]; 
    assign out[3144] = layer_1[3047] & ~layer_1[3166]; 
    assign out[3145] = ~layer_1[3320]; 
    assign out[3146] = ~layer_1[1930]; 
    assign out[3147] = layer_1[152]; 
    assign out[3148] = layer_1[2779]; 
    assign out[3149] = ~layer_1[3067]; 
    assign out[3150] = ~layer_1[3629]; 
    assign out[3151] = layer_1[1278]; 
    assign out[3152] = layer_1[673] & ~layer_1[663]; 
    assign out[3153] = layer_1[3788] ^ layer_1[3676]; 
    assign out[3154] = layer_1[2248]; 
    assign out[3155] = layer_1[1100]; 
    assign out[3156] = ~layer_1[742]; 
    assign out[3157] = ~(layer_1[683] ^ layer_1[694]); 
    assign out[3158] = ~(layer_1[3891] & layer_1[3848]); 
    assign out[3159] = layer_1[3680]; 
    assign out[3160] = layer_1[1182] ^ layer_1[1164]; 
    assign out[3161] = layer_1[3836]; 
    assign out[3162] = layer_1[384] & ~layer_1[332]; 
    assign out[3163] = layer_1[454] | layer_1[445]; 
    assign out[3164] = ~layer_1[3974]; 
    assign out[3165] = layer_1[1738]; 
    assign out[3166] = ~(layer_1[470] ^ layer_1[371]); 
    assign out[3167] = layer_1[38] | layer_1[83]; 
    assign out[3168] = ~(layer_1[3102] & layer_1[3072]); 
    assign out[3169] = layer_1[2474] & ~layer_1[2577]; 
    assign out[3170] = layer_1[371] & layer_1[384]; 
    assign out[3171] = ~layer_1[1718] | (layer_1[1634] & layer_1[1718]); 
    assign out[3172] = layer_1[909] & ~layer_1[1027]; 
    assign out[3173] = ~layer_1[1903]; 
    assign out[3174] = layer_1[1830] ^ layer_1[1704]; 
    assign out[3175] = ~layer_1[2879]; 
    assign out[3176] = ~layer_1[686]; 
    assign out[3177] = ~layer_1[2445]; 
    assign out[3178] = ~(layer_1[3856] & layer_1[3932]); 
    assign out[3179] = layer_1[3035] & layer_1[2978]; 
    assign out[3180] = layer_1[2596] & layer_1[2648]; 
    assign out[3181] = layer_1[1333] | layer_1[1310]; 
    assign out[3182] = layer_1[2634] ^ layer_1[2515]; 
    assign out[3183] = ~(layer_1[1058] ^ layer_1[938]); 
    assign out[3184] = ~layer_1[1542]; 
    assign out[3185] = ~(layer_1[3841] ^ layer_1[3756]); 
    assign out[3186] = ~layer_1[3873]; 
    assign out[3187] = layer_1[1842]; 
    assign out[3188] = ~layer_1[3123]; 
    assign out[3189] = ~(layer_1[2448] & layer_1[2426]); 
    assign out[3190] = ~layer_1[1369] | (layer_1[1418] & layer_1[1369]); 
    assign out[3191] = ~(layer_1[1579] | layer_1[1491]); 
    assign out[3192] = layer_1[1084]; 
    assign out[3193] = ~layer_1[408]; 
    assign out[3194] = ~layer_1[1322]; 
    assign out[3195] = layer_1[909] & ~layer_1[813]; 
    assign out[3196] = ~layer_1[2999]; 
    assign out[3197] = layer_1[3392]; 
    assign out[3198] = layer_1[3575] ^ layer_1[3521]; 
    assign out[3199] = layer_1[3039]; 
    assign out[3200] = layer_1[2733] | layer_1[2671]; 
    assign out[3201] = ~(layer_1[2092] | layer_1[2214]); 
    assign out[3202] = layer_1[2986] & layer_1[3104]; 
    assign out[3203] = layer_1[2974]; 
    assign out[3204] = layer_1[3778]; 
    assign out[3205] = ~(layer_1[2691] ^ layer_1[2683]); 
    assign out[3206] = layer_1[3253] & ~layer_1[3263]; 
    assign out[3207] = ~(layer_1[1195] ^ layer_1[1180]); 
    assign out[3208] = ~(layer_1[2973] | layer_1[3046]); 
    assign out[3209] = layer_1[2959] & ~layer_1[2949]; 
    assign out[3210] = ~(layer_1[795] & layer_1[867]); 
    assign out[3211] = layer_1[1527] & ~layer_1[1589]; 
    assign out[3212] = layer_1[3712]; 
    assign out[3213] = layer_1[465] | layer_1[525]; 
    assign out[3214] = layer_1[1106] & layer_1[1097]; 
    assign out[3215] = layer_1[2031] ^ layer_1[2139]; 
    assign out[3216] = layer_1[45] & ~layer_1[22]; 
    assign out[3217] = ~layer_1[2433]; 
    assign out[3218] = ~layer_1[1618]; 
    assign out[3219] = layer_1[1936] ^ layer_1[2059]; 
    assign out[3220] = layer_1[2855] | layer_1[2758]; 
    assign out[3221] = layer_1[1072] & ~layer_1[1132]; 
    assign out[3222] = layer_1[2305] & ~layer_1[2183]; 
    assign out[3223] = layer_1[1116]; 
    assign out[3224] = layer_1[353] ^ layer_1[252]; 
    assign out[3225] = layer_1[1934] & ~layer_1[2017]; 
    assign out[3226] = layer_1[3942] ^ layer_1[3984]; 
    assign out[3227] = ~(layer_1[2750] | layer_1[2723]); 
    assign out[3228] = ~layer_1[1735]; 
    assign out[3229] = ~(layer_1[2441] ^ layer_1[2408]); 
    assign out[3230] = ~layer_1[1317] | (layer_1[1317] & layer_1[1425]); 
    assign out[3231] = layer_1[3229] ^ layer_1[3267]; 
    assign out[3232] = ~layer_1[173]; 
    assign out[3233] = ~layer_1[718]; 
    assign out[3234] = ~(layer_1[120] ^ layer_1[246]); 
    assign out[3235] = layer_1[2646] ^ layer_1[2535]; 
    assign out[3236] = ~layer_1[589] | (layer_1[589] & layer_1[481]); 
    assign out[3237] = layer_1[1697]; 
    assign out[3238] = ~layer_1[331]; 
    assign out[3239] = layer_1[73] & ~layer_1[135]; 
    assign out[3240] = layer_1[354]; 
    assign out[3241] = layer_1[1449] & layer_1[1361]; 
    assign out[3242] = ~layer_1[3963]; 
    assign out[3243] = ~layer_1[3726]; 
    assign out[3244] = ~(layer_1[2947] ^ layer_1[2958]); 
    assign out[3245] = ~(layer_1[3962] ^ layer_1[3880]); 
    assign out[3246] = ~(layer_1[1159] & layer_1[1161]); 
    assign out[3247] = layer_1[1182] & ~layer_1[1141]; 
    assign out[3248] = ~(layer_1[1343] ^ layer_1[1366]); 
    assign out[3249] = ~(layer_1[992] | layer_1[956]); 
    assign out[3250] = ~(layer_1[3663] ^ layer_1[3575]); 
    assign out[3251] = ~(layer_1[636] & layer_1[682]); 
    assign out[3252] = layer_1[280] | layer_1[281]; 
    assign out[3253] = layer_1[1533] & ~layer_1[1501]; 
    assign out[3254] = layer_1[1449]; 
    assign out[3255] = ~(layer_1[1192] | layer_1[1227]); 
    assign out[3256] = ~(layer_1[444] & layer_1[412]); 
    assign out[3257] = ~(layer_1[853] ^ layer_1[797]); 
    assign out[3258] = layer_1[3778] & ~layer_1[3899]; 
    assign out[3259] = ~(layer_1[1591] | layer_1[1589]); 
    assign out[3260] = layer_1[731] & layer_1[715]; 
    assign out[3261] = layer_1[3626] & layer_1[3674]; 
    assign out[3262] = ~layer_1[1016]; 
    assign out[3263] = ~(layer_1[571] ^ layer_1[456]); 
    assign out[3264] = ~layer_1[2936]; 
    assign out[3265] = layer_1[1201] | layer_1[1223]; 
    assign out[3266] = layer_1[349] | layer_1[408]; 
    assign out[3267] = ~(layer_1[545] ^ layer_1[422]); 
    assign out[3268] = layer_1[2045] ^ layer_1[1968]; 
    assign out[3269] = ~layer_1[3143] | (layer_1[3143] & layer_1[3205]); 
    assign out[3270] = ~(layer_1[723] & layer_1[824]); 
    assign out[3271] = layer_1[3223] ^ layer_1[3206]; 
    assign out[3272] = layer_1[2704]; 
    assign out[3273] = ~layer_1[702]; 
    assign out[3274] = ~(layer_1[1016] | layer_1[1053]); 
    assign out[3275] = ~(layer_1[1274] | layer_1[1256]); 
    assign out[3276] = ~layer_1[153]; 
    assign out[3277] = ~(layer_1[3959] ^ layer_1[3975]); 
    assign out[3278] = layer_1[1738] ^ layer_1[1660]; 
    assign out[3279] = layer_1[2718] & ~layer_1[2796]; 
    assign out[3280] = ~(layer_1[1330] ^ layer_1[1366]); 
    assign out[3281] = ~(layer_1[285] ^ layer_1[265]); 
    assign out[3282] = ~layer_1[2343]; 
    assign out[3283] = ~(layer_1[2714] ^ layer_1[2690]); 
    assign out[3284] = ~layer_1[555]; 
    assign out[3285] = ~layer_1[706] | (layer_1[706] & layer_1[820]); 
    assign out[3286] = ~(layer_1[1123] ^ layer_1[1030]); 
    assign out[3287] = layer_1[3258]; 
    assign out[3288] = ~layer_1[3137] | (layer_1[3182] & layer_1[3137]); 
    assign out[3289] = ~layer_1[671] | (layer_1[671] & layer_1[566]); 
    assign out[3290] = ~(layer_1[915] & layer_1[951]); 
    assign out[3291] = ~(layer_1[208] | layer_1[331]); 
    assign out[3292] = layer_1[1855] & layer_1[1836]; 
    assign out[3293] = layer_1[1547] ^ layer_1[1624]; 
    assign out[3294] = layer_1[127] & ~layer_1[215]; 
    assign out[3295] = ~layer_1[3478]; 
    assign out[3296] = layer_1[1857] & layer_1[1818]; 
    assign out[3297] = layer_1[851] & ~layer_1[880]; 
    assign out[3298] = layer_1[2130] & ~layer_1[2079]; 
    assign out[3299] = layer_1[3889] ^ layer_1[3890]; 
    assign out[3300] = layer_1[1206] | layer_1[1101]; 
    assign out[3301] = ~layer_1[3983]; 
    assign out[3302] = layer_1[2753] & ~layer_1[2836]; 
    assign out[3303] = ~layer_1[2897]; 
    assign out[3304] = ~layer_1[915]; 
    assign out[3305] = ~layer_1[401]; 
    assign out[3306] = layer_1[3032]; 
    assign out[3307] = layer_1[800] ^ layer_1[685]; 
    assign out[3308] = ~layer_1[2007]; 
    assign out[3309] = ~layer_1[1306]; 
    assign out[3310] = layer_1[2152] | layer_1[2114]; 
    assign out[3311] = layer_1[1134] & layer_1[1081]; 
    assign out[3312] = layer_1[1949] ^ layer_1[1836]; 
    assign out[3313] = layer_1[2150] ^ layer_1[2186]; 
    assign out[3314] = layer_1[2572] ^ layer_1[2695]; 
    assign out[3315] = layer_1[1349] | layer_1[1221]; 
    assign out[3316] = ~(layer_1[1904] & layer_1[1967]); 
    assign out[3317] = layer_1[349] | layer_1[325]; 
    assign out[3318] = layer_1[2704] & ~layer_1[2657]; 
    assign out[3319] = layer_1[2111] & ~layer_1[2054]; 
    assign out[3320] = ~layer_1[2227]; 
    assign out[3321] = layer_1[433] ^ layer_1[445]; 
    assign out[3322] = layer_1[1038]; 
    assign out[3323] = layer_1[1753] ^ layer_1[1849]; 
    assign out[3324] = ~layer_1[3560] | (layer_1[3560] & layer_1[3617]); 
    assign out[3325] = layer_1[1554]; 
    assign out[3326] = layer_1[3176] & layer_1[3072]; 
    assign out[3327] = ~layer_1[2465]; 
    assign out[3328] = layer_1[3457] & ~layer_1[3560]; 
    assign out[3329] = layer_1[612] & ~layer_1[725]; 
    assign out[3330] = layer_1[2860]; 
    assign out[3331] = ~(layer_1[2898] | layer_1[2978]); 
    assign out[3332] = ~layer_1[795] | (layer_1[903] & layer_1[795]); 
    assign out[3333] = layer_1[845] & ~layer_1[808]; 
    assign out[3334] = ~(layer_1[3864] ^ layer_1[3844]); 
    assign out[3335] = layer_1[1331] ^ layer_1[1311]; 
    assign out[3336] = ~layer_1[3599]; 
    assign out[3337] = layer_1[3576] & layer_1[3501]; 
    assign out[3338] = ~layer_1[2586]; 
    assign out[3339] = layer_1[2515]; 
    assign out[3340] = ~(layer_1[1760] ^ layer_1[1883]); 
    assign out[3341] = layer_1[1610] & ~layer_1[1700]; 
    assign out[3342] = ~layer_1[1972]; 
    assign out[3343] = layer_1[492] ^ layer_1[394]; 
    assign out[3344] = layer_1[2233] & layer_1[2179]; 
    assign out[3345] = ~(layer_1[1096] ^ layer_1[1130]); 
    assign out[3346] = layer_1[451]; 
    assign out[3347] = ~layer_1[2961]; 
    assign out[3348] = ~layer_1[1889] | (layer_1[1889] & layer_1[1783]); 
    assign out[3349] = layer_1[334] & ~layer_1[208]; 
    assign out[3350] = ~layer_1[824] | (layer_1[824] & layer_1[879]); 
    assign out[3351] = layer_1[3176] ^ layer_1[3178]; 
    assign out[3352] = ~layer_1[1690]; 
    assign out[3353] = layer_1[1615] | layer_1[1718]; 
    assign out[3354] = ~(layer_1[1969] ^ layer_1[2022]); 
    assign out[3355] = ~layer_1[1598] | (layer_1[1651] & layer_1[1598]); 
    assign out[3356] = ~(layer_1[2885] ^ layer_1[3001]); 
    assign out[3357] = ~layer_1[319] | (layer_1[319] & layer_1[354]); 
    assign out[3358] = ~layer_1[200]; 
    assign out[3359] = layer_1[1405] ^ layer_1[1333]; 
    assign out[3360] = ~(layer_1[2542] ^ layer_1[2573]); 
    assign out[3361] = layer_1[3149] ^ layer_1[3179]; 
    assign out[3362] = ~(layer_1[433] | layer_1[456]); 
    assign out[3363] = layer_1[1127] & ~layer_1[1183]; 
    assign out[3364] = ~layer_1[2752] | (layer_1[2860] & layer_1[2752]); 
    assign out[3365] = layer_1[1819] & ~layer_1[1794]; 
    assign out[3366] = layer_1[97]; 
    assign out[3367] = ~layer_1[1598]; 
    assign out[3368] = ~layer_1[2350]; 
    assign out[3369] = ~layer_1[1482]; 
    assign out[3370] = layer_1[1853] & layer_1[1847]; 
    assign out[3371] = layer_1[2737] & layer_1[2833]; 
    assign out[3372] = layer_1[279] & ~layer_1[328]; 
    assign out[3373] = layer_1[3343]; 
    assign out[3374] = layer_1[309] ^ layer_1[252]; 
    assign out[3375] = ~layer_1[1424] | (layer_1[1424] & layer_1[1546]); 
    assign out[3376] = ~(layer_1[3808] | layer_1[3779]); 
    assign out[3377] = ~(layer_1[3419] ^ layer_1[3400]); 
    assign out[3378] = layer_1[843] & layer_1[955]; 
    assign out[3379] = layer_1[510]; 
    assign out[3380] = layer_1[2101] ^ layer_1[2109]; 
    assign out[3381] = ~layer_1[539]; 
    assign out[3382] = ~layer_1[1210] | (layer_1[1210] & layer_1[1253]); 
    assign out[3383] = ~(layer_1[1688] & layer_1[1617]); 
    assign out[3384] = ~(layer_1[3056] ^ layer_1[2978]); 
    assign out[3385] = layer_1[2368] & ~layer_1[2463]; 
    assign out[3386] = layer_1[3342]; 
    assign out[3387] = layer_1[1521]; 
    assign out[3388] = layer_1[3209] & layer_1[3142]; 
    assign out[3389] = layer_1[802] & ~layer_1[927]; 
    assign out[3390] = ~(layer_1[1535] ^ layer_1[1643]); 
    assign out[3391] = layer_1[408]; 
    assign out[3392] = ~(layer_1[3451] ^ layer_1[3430]); 
    assign out[3393] = layer_1[3469]; 
    assign out[3394] = layer_1[3927]; 
    assign out[3395] = ~layer_1[2009] | (layer_1[2072] & layer_1[2009]); 
    assign out[3396] = layer_1[229]; 
    assign out[3397] = layer_1[2256]; 
    assign out[3398] = ~(layer_1[444] | layer_1[378]); 
    assign out[3399] = layer_1[921]; 
    assign out[3400] = ~layer_1[3245]; 
    assign out[3401] = layer_1[408]; 
    assign out[3402] = layer_1[1451]; 
    assign out[3403] = ~layer_1[3452] | (layer_1[3452] & layer_1[3393]); 
    assign out[3404] = layer_1[3539] ^ layer_1[3534]; 
    assign out[3405] = ~(layer_1[2425] | layer_1[2471]); 
    assign out[3406] = ~(layer_1[789] ^ layer_1[696]); 
    assign out[3407] = layer_1[669]; 
    assign out[3408] = layer_1[308] & ~layer_1[215]; 
    assign out[3409] = layer_1[3596] ^ layer_1[3693]; 
    assign out[3410] = ~(layer_1[3561] ^ layer_1[3448]); 
    assign out[3411] = ~(layer_1[1398] ^ layer_1[1415]); 
    assign out[3412] = ~layer_1[3115] | (layer_1[3096] & layer_1[3115]); 
    assign out[3413] = ~(layer_1[1057] | layer_1[992]); 
    assign out[3414] = layer_1[3585] ^ layer_1[3486]; 
    assign out[3415] = ~layer_1[173]; 
    assign out[3416] = ~(layer_1[1777] ^ layer_1[1848]); 
    assign out[3417] = ~(layer_1[2083] ^ layer_1[2112]); 
    assign out[3418] = layer_1[154]; 
    assign out[3419] = ~(layer_1[2945] | layer_1[2984]); 
    assign out[3420] = ~(layer_1[66] ^ layer_1[142]); 
    assign out[3421] = ~layer_1[3119] | (layer_1[3147] & layer_1[3119]); 
    assign out[3422] = ~layer_1[3405]; 
    assign out[3423] = layer_1[2526] & ~layer_1[2522]; 
    assign out[3424] = ~(layer_1[456] ^ layer_1[421]); 
    assign out[3425] = layer_1[2189] ^ layer_1[2251]; 
    assign out[3426] = layer_1[186]; 
    assign out[3427] = ~layer_1[547]; 
    assign out[3428] = ~layer_1[208]; 
    assign out[3429] = ~(layer_1[1168] ^ layer_1[1042]); 
    assign out[3430] = layer_1[3877] & ~layer_1[3791]; 
    assign out[3431] = layer_1[2842]; 
    assign out[3432] = ~layer_1[1078]; 
    assign out[3433] = ~layer_1[3713]; 
    assign out[3434] = layer_1[1086] & ~layer_1[1183]; 
    assign out[3435] = layer_1[3168] & layer_1[3285]; 
    assign out[3436] = ~(layer_1[1789] | layer_1[1770]); 
    assign out[3437] = ~layer_1[773]; 
    assign out[3438] = ~(layer_1[1797] | layer_1[1759]); 
    assign out[3439] = ~(layer_1[438] | layer_1[400]); 
    assign out[3440] = ~layer_1[1810]; 
    assign out[3441] = ~(layer_1[1794] | layer_1[1885]); 
    assign out[3442] = layer_1[2134] & layer_1[2255]; 
    assign out[3443] = ~layer_1[2960]; 
    assign out[3444] = ~(layer_1[3379] ^ layer_1[3264]); 
    assign out[3445] = layer_1[3290]; 
    assign out[3446] = layer_1[3548]; 
    assign out[3447] = ~(layer_1[2470] | layer_1[2349]); 
    assign out[3448] = layer_1[1954] & layer_1[2047]; 
    assign out[3449] = ~(layer_1[1719] ^ layer_1[1765]); 
    assign out[3450] = layer_1[3300]; 
    assign out[3451] = layer_1[422]; 
    assign out[3452] = layer_1[341] & ~layer_1[355]; 
    assign out[3453] = ~layer_1[3297]; 
    assign out[3454] = layer_1[1481] | layer_1[1397]; 
    assign out[3455] = layer_1[2833] & layer_1[2847]; 
    assign out[3456] = layer_1[2753] & ~layer_1[2816]; 
    assign out[3457] = layer_1[2418] ^ layer_1[2506]; 
    assign out[3458] = layer_1[1833] ^ layer_1[1788]; 
    assign out[3459] = layer_1[804] ^ layer_1[745]; 
    assign out[3460] = ~layer_1[1904]; 
    assign out[3461] = layer_1[698] & layer_1[793]; 
    assign out[3462] = layer_1[536] & layer_1[578]; 
    assign out[3463] = ~(layer_1[1020] & layer_1[1071]); 
    assign out[3464] = layer_1[27]; 
    assign out[3465] = ~(layer_1[2183] | layer_1[2227]); 
    assign out[3466] = ~layer_1[2853]; 
    assign out[3467] = ~(layer_1[3710] | layer_1[3698]); 
    assign out[3468] = ~(layer_1[3273] ^ layer_1[3249]); 
    assign out[3469] = ~layer_1[147]; 
    assign out[3470] = layer_1[1500] ^ layer_1[1432]; 
    assign out[3471] = ~(layer_1[1499] | layer_1[1399]); 
    assign out[3472] = layer_1[607] ^ layer_1[552]; 
    assign out[3473] = layer_1[2500] ^ layer_1[2455]; 
    assign out[3474] = layer_1[2679] ^ layer_1[2653]; 
    assign out[3475] = ~(layer_1[1866] & layer_1[1917]); 
    assign out[3476] = layer_1[352]; 
    assign out[3477] = layer_1[1357] & ~layer_1[1233]; 
    assign out[3478] = layer_1[2649] & ~layer_1[2748]; 
    assign out[3479] = ~layer_1[3828]; 
    assign out[3480] = ~layer_1[654] | (layer_1[654] & layer_1[616]); 
    assign out[3481] = ~layer_1[2924]; 
    assign out[3482] = layer_1[832]; 
    assign out[3483] = layer_1[179] & ~layer_1[90]; 
    assign out[3484] = ~(layer_1[869] | layer_1[757]); 
    assign out[3485] = ~(layer_1[1978] | layer_1[2015]); 
    assign out[3486] = layer_1[175] ^ layer_1[195]; 
    assign out[3487] = ~layer_1[1281] | (layer_1[1281] & layer_1[1349]); 
    assign out[3488] = ~layer_1[1407] | (layer_1[1445] & layer_1[1407]); 
    assign out[3489] = layer_1[1095]; 
    assign out[3490] = layer_1[3333]; 
    assign out[3491] = layer_1[851] & ~layer_1[817]; 
    assign out[3492] = layer_1[406] ^ layer_1[354]; 
    assign out[3493] = layer_1[1147] ^ layer_1[1141]; 
    assign out[3494] = layer_1[2449] & ~layer_1[2382]; 
    assign out[3495] = layer_1[881]; 
    assign out[3496] = ~layer_1[3630]; 
    assign out[3497] = layer_1[827]; 
    assign out[3498] = ~layer_1[1374]; 
    assign out[3499] = ~layer_1[71]; 
    assign out[3500] = ~(layer_1[1861] ^ layer_1[1853]); 
    assign out[3501] = layer_1[3191] ^ layer_1[3149]; 
    assign out[3502] = layer_1[264] & layer_1[229]; 
    assign out[3503] = layer_1[2581] & layer_1[2456]; 
    assign out[3504] = layer_1[3531] & ~layer_1[3492]; 
    assign out[3505] = ~layer_1[291]; 
    assign out[3506] = ~(layer_1[372] ^ layer_1[365]); 
    assign out[3507] = ~(layer_1[877] ^ layer_1[1001]); 
    assign out[3508] = layer_1[3096] & ~layer_1[2996]; 
    assign out[3509] = layer_1[1060]; 
    assign out[3510] = ~layer_1[2877]; 
    assign out[3511] = layer_1[2286]; 
    assign out[3512] = ~(layer_1[3395] | layer_1[3498]); 
    assign out[3513] = layer_1[3350] ^ layer_1[3348]; 
    assign out[3514] = layer_1[550]; 
    assign out[3515] = ~layer_1[2862] | (layer_1[2860] & layer_1[2862]); 
    assign out[3516] = layer_1[2930] & ~layer_1[3052]; 
    assign out[3517] = layer_1[565]; 
    assign out[3518] = ~(layer_1[1020] ^ layer_1[1006]); 
    assign out[3519] = ~layer_1[3492]; 
    assign out[3520] = ~layer_1[3250]; 
    assign out[3521] = layer_1[3201] & ~layer_1[3219]; 
    assign out[3522] = ~(layer_1[3715] | layer_1[3616]); 
    assign out[3523] = ~layer_1[3608]; 
    assign out[3524] = layer_1[127] & ~layer_1[120]; 
    assign out[3525] = ~(layer_1[2299] ^ layer_1[2271]); 
    assign out[3526] = ~layer_1[597]; 
    assign out[3527] = ~layer_1[2638]; 
    assign out[3528] = layer_1[2351]; 
    assign out[3529] = layer_1[2393] & ~layer_1[2465]; 
    assign out[3530] = layer_1[3941] ^ layer_1[3980]; 
    assign out[3531] = layer_1[3454] & layer_1[3491]; 
    assign out[3532] = layer_1[1806] | layer_1[1680]; 
    assign out[3533] = layer_1[1323] & ~layer_1[1287]; 
    assign out[3534] = layer_1[3524] ^ layer_1[3505]; 
    assign out[3535] = layer_1[1899] ^ layer_1[1927]; 
    assign out[3536] = layer_1[659]; 
    assign out[3537] = layer_1[3965]; 
    assign out[3538] = layer_1[3289] & ~layer_1[3406]; 
    assign out[3539] = layer_1[3180] & ~layer_1[3058]; 
    assign out[3540] = ~(layer_1[1713] ^ layer_1[1813]); 
    assign out[3541] = ~(layer_1[3137] & layer_1[3046]); 
    assign out[3542] = layer_1[2247]; 
    assign out[3543] = ~layer_1[677]; 
    assign out[3544] = layer_1[756] & ~layer_1[864]; 
    assign out[3545] = layer_1[1366] ^ layer_1[1280]; 
    assign out[3546] = ~layer_1[1539]; 
    assign out[3547] = ~(layer_1[626] | layer_1[664]); 
    assign out[3548] = layer_1[3159] & ~layer_1[3164]; 
    assign out[3549] = layer_1[108] & layer_1[79]; 
    assign out[3550] = layer_1[70] | layer_1[99]; 
    assign out[3551] = ~(layer_1[2816] | layer_1[2898]); 
    assign out[3552] = layer_1[1358] & ~layer_1[1375]; 
    assign out[3553] = layer_1[1461] | layer_1[1338]; 
    assign out[3554] = layer_1[2508] & layer_1[2461]; 
    assign out[3555] = layer_1[862] ^ layer_1[955]; 
    assign out[3556] = layer_1[1449] & layer_1[1532]; 
    assign out[3557] = layer_1[3201]; 
    assign out[3558] = ~(layer_1[1339] & layer_1[1454]); 
    assign out[3559] = layer_1[27] & layer_1[118]; 
    assign out[3560] = ~layer_1[3046] | (layer_1[3114] & layer_1[3046]); 
    assign out[3561] = layer_1[1670] | layer_1[1653]; 
    assign out[3562] = layer_1[2517]; 
    assign out[3563] = ~(layer_1[3259] ^ layer_1[3167]); 
    assign out[3564] = ~layer_1[558]; 
    assign out[3565] = layer_1[1253] ^ layer_1[1252]; 
    assign out[3566] = ~layer_1[1556]; 
    assign out[3567] = ~(layer_1[3532] | layer_1[3586]); 
    assign out[3568] = ~layer_1[338]; 
    assign out[3569] = ~(layer_1[2576] ^ layer_1[2483]); 
    assign out[3570] = ~(layer_1[2476] ^ layer_1[2367]); 
    assign out[3571] = layer_1[2236]; 
    assign out[3572] = layer_1[3528]; 
    assign out[3573] = ~layer_1[1871]; 
    assign out[3574] = layer_1[465] | layer_1[490]; 
    assign out[3575] = ~(layer_1[1071] & layer_1[1062]); 
    assign out[3576] = layer_1[2457] & ~layer_1[2454]; 
    assign out[3577] = ~layer_1[1010]; 
    assign out[3578] = ~(layer_1[3326] | layer_1[3292]); 
    assign out[3579] = ~(layer_1[3399] | layer_1[3487]); 
    assign out[3580] = layer_1[3505] & layer_1[3546]; 
    assign out[3581] = ~layer_1[2625]; 
    assign out[3582] = ~(layer_1[1743] ^ layer_1[1658]); 
    assign out[3583] = ~(layer_1[3855] | layer_1[3970]); 
    assign out[3584] = ~layer_1[703]; 
    assign out[3585] = layer_1[3114]; 
    assign out[3586] = layer_1[1470] & layer_1[1490]; 
    assign out[3587] = layer_1[1605] & layer_1[1647]; 
    assign out[3588] = ~layer_1[670] | (layer_1[576] & layer_1[670]); 
    assign out[3589] = ~(layer_1[133] ^ layer_1[183]); 
    assign out[3590] = layer_1[2296] ^ layer_1[2315]; 
    assign out[3591] = ~layer_1[1120]; 
    assign out[3592] = layer_1[1356]; 
    assign out[3593] = ~(layer_1[3095] | layer_1[3164]); 
    assign out[3594] = layer_1[2610] & ~layer_1[2681]; 
    assign out[3595] = ~(layer_1[1336] ^ layer_1[1453]); 
    assign out[3596] = ~(layer_1[3194] ^ layer_1[3125]); 
    assign out[3597] = ~layer_1[147]; 
    assign out[3598] = ~layer_1[15]; 
    assign out[3599] = layer_1[951] ^ layer_1[1005]; 
    assign out[3600] = ~(layer_1[2838] | layer_1[2940]); 
    assign out[3601] = layer_1[1780] & ~layer_1[1852]; 
    assign out[3602] = layer_1[1052] & ~layer_1[1008]; 
    assign out[3603] = layer_1[2647]; 
    assign out[3604] = layer_1[814] & ~layer_1[800]; 
    assign out[3605] = layer_1[1954] & layer_1[1827]; 
    assign out[3606] = layer_1[1963] & ~layer_1[2012]; 
    assign out[3607] = ~layer_1[975]; 
    assign out[3608] = layer_1[1747] & ~layer_1[1816]; 
    assign out[3609] = layer_1[26] & layer_1[90]; 
    assign out[3610] = layer_1[2367] ^ layer_1[2281]; 
    assign out[3611] = layer_1[3720] & ~layer_1[3728]; 
    assign out[3612] = ~layer_1[2898]; 
    assign out[3613] = ~layer_1[3434] | (layer_1[3434] & layer_1[3329]); 
    assign out[3614] = layer_1[387] & ~layer_1[292]; 
    assign out[3615] = layer_1[114] & ~layer_1[190]; 
    assign out[3616] = ~layer_1[815]; 
    assign out[3617] = ~layer_1[1899]; 
    assign out[3618] = layer_1[1496]; 
    assign out[3619] = layer_1[9] | layer_1[51]; 
    assign out[3620] = layer_1[3840] & layer_1[3967]; 
    assign out[3621] = ~layer_1[696]; 
    assign out[3622] = layer_1[3226] & layer_1[3150]; 
    assign out[3623] = layer_1[925] ^ layer_1[911]; 
    assign out[3624] = layer_1[1257] & ~layer_1[1279]; 
    assign out[3625] = ~(layer_1[3782] | layer_1[3694]); 
    assign out[3626] = layer_1[2981] & ~layer_1[3092]; 
    assign out[3627] = ~layer_1[2910]; 
    assign out[3628] = layer_1[2993] & ~layer_1[2928]; 
    assign out[3629] = layer_1[3044] & layer_1[3143]; 
    assign out[3630] = ~layer_1[3978]; 
    assign out[3631] = layer_1[3176] & ~layer_1[3095]; 
    assign out[3632] = layer_1[3332] | layer_1[3353]; 
    assign out[3633] = ~(layer_1[2131] | layer_1[2115]); 
    assign out[3634] = layer_1[3246]; 
    assign out[3635] = ~layer_1[2358]; 
    assign out[3636] = ~layer_1[3729]; 
    assign out[3637] = layer_1[2000] & layer_1[1941]; 
    assign out[3638] = ~(layer_1[948] & layer_1[832]); 
    assign out[3639] = ~(layer_1[2405] ^ layer_1[2463]); 
    assign out[3640] = ~layer_1[3815]; 
    assign out[3641] = ~(layer_1[2557] ^ layer_1[2606]); 
    assign out[3642] = layer_1[3771] & ~layer_1[3818]; 
    assign out[3643] = ~layer_1[3322]; 
    assign out[3644] = layer_1[722]; 
    assign out[3645] = ~(layer_1[3811] ^ layer_1[3759]); 
    assign out[3646] = layer_1[2152]; 
    assign out[3647] = ~layer_1[3279] | (layer_1[3279] & layer_1[3245]); 
    assign out[3648] = layer_1[2614] & layer_1[2694]; 
    assign out[3649] = layer_1[1992] & layer_1[2070]; 
    assign out[3650] = layer_1[822] & ~layer_1[910]; 
    assign out[3651] = layer_1[1807]; 
    assign out[3652] = ~(layer_1[2201] ^ layer_1[2203]); 
    assign out[3653] = ~layer_1[2901]; 
    assign out[3654] = layer_1[2169] ^ layer_1[2296]; 
    assign out[3655] = layer_1[2363]; 
    assign out[3656] = ~(layer_1[860] & layer_1[756]); 
    assign out[3657] = ~(layer_1[248] | layer_1[199]); 
    assign out[3658] = ~(layer_1[46] | layer_1[68]); 
    assign out[3659] = layer_1[2990] ^ layer_1[3099]; 
    assign out[3660] = ~layer_1[3513]; 
    assign out[3661] = layer_1[359] & ~layer_1[345]; 
    assign out[3662] = ~(layer_1[1974] ^ layer_1[1870]); 
    assign out[3663] = ~layer_1[124] | (layer_1[107] & layer_1[124]); 
    assign out[3664] = layer_1[1209] & ~layer_1[1329]; 
    assign out[3665] = layer_1[1550] & ~layer_1[1497]; 
    assign out[3666] = ~(layer_1[3653] | layer_1[3656]); 
    assign out[3667] = ~layer_1[599]; 
    assign out[3668] = layer_1[1692] & ~layer_1[1753]; 
    assign out[3669] = layer_1[2891] & ~layer_1[2804]; 
    assign out[3670] = layer_1[2164] & ~layer_1[2169]; 
    assign out[3671] = layer_1[2185]; 
    assign out[3672] = ~(layer_1[2364] ^ layer_1[2443]); 
    assign out[3673] = layer_1[2489] ^ layer_1[2412]; 
    assign out[3674] = ~layer_1[3168]; 
    assign out[3675] = ~(layer_1[2715] | layer_1[2680]); 
    assign out[3676] = ~layer_1[1573] | (layer_1[1556] & layer_1[1573]); 
    assign out[3677] = ~(layer_1[1954] ^ layer_1[2058]); 
    assign out[3678] = layer_1[2563]; 
    assign out[3679] = layer_1[844]; 
    assign out[3680] = ~(layer_1[276] | layer_1[326]); 
    assign out[3681] = layer_1[1910] & ~layer_1[2001]; 
    assign out[3682] = layer_1[3077] & layer_1[3162]; 
    assign out[3683] = ~layer_1[495]; 
    assign out[3684] = layer_1[1097] & layer_1[1203]; 
    assign out[3685] = ~layer_1[3858]; 
    assign out[3686] = layer_1[1787] & ~layer_1[1781]; 
    assign out[3687] = layer_1[1496]; 
    assign out[3688] = layer_1[3805] & ~layer_1[3786]; 
    assign out[3689] = layer_1[3267]; 
    assign out[3690] = layer_1[1131] ^ layer_1[1128]; 
    assign out[3691] = ~layer_1[3663] | (layer_1[3663] & layer_1[3687]); 
    assign out[3692] = ~(layer_1[2784] | layer_1[2693]); 
    assign out[3693] = layer_1[907] & ~layer_1[832]; 
    assign out[3694] = ~layer_1[2686]; 
    assign out[3695] = layer_1[191]; 
    assign out[3696] = layer_1[3713] & ~layer_1[3803]; 
    assign out[3697] = layer_1[2682]; 
    assign out[3698] = ~(layer_1[1266] ^ layer_1[1175]); 
    assign out[3699] = layer_1[2593] ^ layer_1[2657]; 
    assign out[3700] = layer_1[2891]; 
    assign out[3701] = layer_1[1427]; 
    assign out[3702] = layer_1[1565] ^ layer_1[1545]; 
    assign out[3703] = ~layer_1[1619]; 
    assign out[3704] = ~(layer_1[2869] ^ layer_1[2892]); 
    assign out[3705] = layer_1[608] ^ layer_1[567]; 
    assign out[3706] = layer_1[1439]; 
    assign out[3707] = ~layer_1[920]; 
    assign out[3708] = layer_1[2488] & layer_1[2366]; 
    assign out[3709] = layer_1[1983] ^ layer_1[1940]; 
    assign out[3710] = layer_1[3198] ^ layer_1[3077]; 
    assign out[3711] = layer_1[1331] & ~layer_1[1378]; 
    assign out[3712] = layer_1[304] & layer_1[393]; 
    assign out[3713] = ~layer_1[3537]; 
    assign out[3714] = ~(layer_1[2395] | layer_1[2420]); 
    assign out[3715] = layer_1[1433]; 
    assign out[3716] = layer_1[1842] & ~layer_1[1968]; 
    assign out[3717] = ~layer_1[2789]; 
    assign out[3718] = layer_1[3197] & ~layer_1[3302]; 
    assign out[3719] = ~(layer_1[1115] ^ layer_1[1130]); 
    assign out[3720] = ~(layer_1[3544] | layer_1[3586]); 
    assign out[3721] = ~layer_1[3572]; 
    assign out[3722] = layer_1[702]; 
    assign out[3723] = ~layer_1[148]; 
    assign out[3724] = layer_1[3708]; 
    assign out[3725] = ~layer_1[1982] | (layer_1[1982] & layer_1[2029]); 
    assign out[3726] = ~(layer_1[599] ^ layer_1[536]); 
    assign out[3727] = layer_1[1033] & ~layer_1[1072]; 
    assign out[3728] = layer_1[3090]; 
    assign out[3729] = ~layer_1[3199]; 
    assign out[3730] = ~layer_1[2485]; 
    assign out[3731] = ~layer_1[1473]; 
    assign out[3732] = layer_1[1749] & ~layer_1[1740]; 
    assign out[3733] = ~layer_1[1089]; 
    assign out[3734] = layer_1[1760] ^ layer_1[1695]; 
    assign out[3735] = layer_1[79]; 
    assign out[3736] = ~(layer_1[2372] | layer_1[2251]); 
    assign out[3737] = ~(layer_1[3977] ^ layer_1[3865]); 
    assign out[3738] = layer_1[2227] & ~layer_1[2286]; 
    assign out[3739] = layer_1[428]; 
    assign out[3740] = ~(layer_1[1535] | layer_1[1494]); 
    assign out[3741] = layer_1[2118] & ~layer_1[2136]; 
    assign out[3742] = layer_1[2777] & ~layer_1[2804]; 
    assign out[3743] = ~(layer_1[1999] | layer_1[1933]); 
    assign out[3744] = layer_1[2057]; 
    assign out[3745] = ~(layer_1[3315] | layer_1[3421]); 
    assign out[3746] = layer_1[2101] ^ layer_1[1987]; 
    assign out[3747] = layer_1[1891]; 
    assign out[3748] = ~(layer_1[2296] | layer_1[2189]); 
    assign out[3749] = ~layer_1[2988]; 
    assign out[3750] = layer_1[3869] & layer_1[3882]; 
    assign out[3751] = layer_1[1832]; 
    assign out[3752] = layer_1[346]; 
    assign out[3753] = ~layer_1[296] | (layer_1[296] & layer_1[177]); 
    assign out[3754] = layer_1[3822] & ~layer_1[3854]; 
    assign out[3755] = layer_1[3831] | layer_1[3820]; 
    assign out[3756] = layer_1[3115]; 
    assign out[3757] = ~layer_1[2869] | (layer_1[2816] & layer_1[2869]); 
    assign out[3758] = layer_1[925]; 
    assign out[3759] = layer_1[2411]; 
    assign out[3760] = ~(layer_1[2126] | layer_1[2043]); 
    assign out[3761] = layer_1[1646] | layer_1[1612]; 
    assign out[3762] = layer_1[1102] & layer_1[1123]; 
    assign out[3763] = ~(layer_1[1841] ^ layer_1[1920]); 
    assign out[3764] = ~layer_1[2493]; 
    assign out[3765] = layer_1[423] & layer_1[539]; 
    assign out[3766] = ~(layer_1[2013] | layer_1[2123]); 
    assign out[3767] = layer_1[19] & ~layer_1[28]; 
    assign out[3768] = ~(layer_1[3201] ^ layer_1[3188]); 
    assign out[3769] = layer_1[1531] & ~layer_1[1609]; 
    assign out[3770] = layer_1[2492] & ~layer_1[2370]; 
    assign out[3771] = layer_1[3077] & ~layer_1[3037]; 
    assign out[3772] = ~(layer_1[774] | layer_1[884]); 
    assign out[3773] = layer_1[1243] & layer_1[1205]; 
    assign out[3774] = layer_1[1770]; 
    assign out[3775] = layer_1[528]; 
    assign out[3776] = ~layer_1[3754]; 
    assign out[3777] = layer_1[1831] & ~layer_1[1839]; 
    assign out[3778] = ~(layer_1[752] | layer_1[723]); 
    assign out[3779] = ~layer_1[211]; 
    assign out[3780] = layer_1[2481] ^ layer_1[2368]; 
    assign out[3781] = ~(layer_1[3514] | layer_1[3473]); 
    assign out[3782] = layer_1[997] & layer_1[1047]; 
    assign out[3783] = ~(layer_1[3855] & layer_1[3964]); 
    assign out[3784] = ~layer_1[3336]; 
    assign out[3785] = layer_1[639] & ~layer_1[707]; 
    assign out[3786] = ~layer_1[756]; 
    assign out[3787] = layer_1[471] ^ layer_1[379]; 
    assign out[3788] = layer_1[743]; 
    assign out[3789] = ~layer_1[1473]; 
    assign out[3790] = layer_1[2853] | layer_1[2739]; 
    assign out[3791] = ~(layer_1[3470] | layer_1[3509]); 
    assign out[3792] = layer_1[3764] & layer_1[3773]; 
    assign out[3793] = layer_1[1489]; 
    assign out[3794] = layer_1[2077] & layer_1[2081]; 
    assign out[3795] = layer_1[3910] & ~layer_1[3919]; 
    assign out[3796] = layer_1[2877]; 
    assign out[3797] = ~(layer_1[140] ^ layer_1[87]); 
    assign out[3798] = ~(layer_1[2985] | layer_1[3067]); 
    assign out[3799] = ~layer_1[2980] | (layer_1[3015] & layer_1[2980]); 
    assign out[3800] = ~(layer_1[1278] | layer_1[1300]); 
    assign out[3801] = layer_1[365] & ~layer_1[427]; 
    assign out[3802] = ~(layer_1[536] | layer_1[562]); 
    assign out[3803] = ~(layer_1[2744] ^ layer_1[2774]); 
    assign out[3804] = layer_1[3813] & ~layer_1[3740]; 
    assign out[3805] = layer_1[1724] & layer_1[1814]; 
    assign out[3806] = layer_1[348] ^ layer_1[452]; 
    assign out[3807] = layer_1[3908]; 
    assign out[3808] = layer_1[2032] & ~layer_1[2028]; 
    assign out[3809] = layer_1[2750] & ~layer_1[2870]; 
    assign out[3810] = layer_1[2375] & layer_1[2317]; 
    assign out[3811] = ~layer_1[1142]; 
    assign out[3812] = layer_1[2716]; 
    assign out[3813] = ~layer_1[1360] | (layer_1[1360] & layer_1[1298]); 
    assign out[3814] = ~(layer_1[3513] | layer_1[3473]); 
    assign out[3815] = ~(layer_1[2827] ^ layer_1[2767]); 
    assign out[3816] = layer_1[2118] & ~layer_1[2016]; 
    assign out[3817] = ~(layer_1[3036] | layer_1[3103]); 
    assign out[3818] = ~(layer_1[1109] ^ layer_1[1097]); 
    assign out[3819] = ~layer_1[3168]; 
    assign out[3820] = layer_1[559] & ~layer_1[505]; 
    assign out[3821] = ~layer_1[957]; 
    assign out[3822] = layer_1[3963] ^ layer_1[3970]; 
    assign out[3823] = ~(layer_1[443] ^ layer_1[519]); 
    assign out[3824] = layer_1[233]; 
    assign out[3825] = ~layer_1[1184]; 
    assign out[3826] = ~layer_1[3520]; 
    assign out[3827] = layer_1[3562]; 
    assign out[3828] = ~(layer_1[2067] ^ layer_1[1972]); 
    assign out[3829] = layer_1[602] ^ layer_1[701]; 
    assign out[3830] = ~layer_1[2205]; 
    assign out[3831] = ~(layer_1[2758] | layer_1[2675]); 
    assign out[3832] = layer_1[305] & layer_1[395]; 
    assign out[3833] = ~layer_1[1158]; 
    assign out[3834] = layer_1[1866]; 
    assign out[3835] = layer_1[3955]; 
    assign out[3836] = layer_1[3749] & ~layer_1[3646]; 
    assign out[3837] = layer_1[2428] & layer_1[2365]; 
    assign out[3838] = layer_1[3139] ^ layer_1[3027]; 
    assign out[3839] = layer_1[208] ^ layer_1[106]; 
    assign out[3840] = layer_1[171] ^ layer_1[266]; 
    assign out[3841] = layer_1[1682]; 
    assign out[3842] = layer_1[2104] & ~layer_1[2166]; 
    assign out[3843] = layer_1[1284] & layer_1[1174]; 
    assign out[3844] = layer_1[2704]; 
    assign out[3845] = layer_1[2480] & ~layer_1[2395]; 
    assign out[3846] = ~(layer_1[2165] ^ layer_1[2091]); 
    assign out[3847] = layer_1[2879]; 
    assign out[3848] = layer_1[2287] & ~layer_1[2280]; 
    assign out[3849] = layer_1[2222] ^ layer_1[2186]; 
    assign out[3850] = layer_1[1558]; 
    assign out[3851] = layer_1[3931] & ~layer_1[3944]; 
    assign out[3852] = ~layer_1[2958]; 
    assign out[3853] = layer_1[969] & ~layer_1[1004]; 
    assign out[3854] = layer_1[3286] & layer_1[3191]; 
    assign out[3855] = layer_1[3714] & ~layer_1[3655]; 
    assign out[3856] = layer_1[3089] & ~layer_1[3033]; 
    assign out[3857] = layer_1[2090] & ~layer_1[2071]; 
    assign out[3858] = layer_1[389]; 
    assign out[3859] = layer_1[3418] & layer_1[3372]; 
    assign out[3860] = ~(layer_1[2555] ^ layer_1[2618]); 
    assign out[3861] = ~(layer_1[2714] | layer_1[2629]); 
    assign out[3862] = ~layer_1[1466]; 
    assign out[3863] = ~(layer_1[3696] | layer_1[3693]); 
    assign out[3864] = layer_1[2057] & layer_1[1997]; 
    assign out[3865] = layer_1[2881] ^ layer_1[2941]; 
    assign out[3866] = layer_1[3064] ^ layer_1[3039]; 
    assign out[3867] = ~layer_1[1432]; 
    assign out[3868] = layer_1[1538] ^ layer_1[1491]; 
    assign out[3869] = layer_1[3143] & layer_1[3015]; 
    assign out[3870] = layer_1[149] ^ layer_1[269]; 
    assign out[3871] = ~layer_1[3509] | (layer_1[3550] & layer_1[3509]); 
    assign out[3872] = ~layer_1[2071]; 
    assign out[3873] = ~(layer_1[377] ^ layer_1[426]); 
    assign out[3874] = layer_1[843] & layer_1[806]; 
    assign out[3875] = layer_1[677] & layer_1[555]; 
    assign out[3876] = layer_1[1512] & ~layer_1[1530]; 
    assign out[3877] = layer_1[517] ^ layer_1[411]; 
    assign out[3878] = ~layer_1[660]; 
    assign out[3879] = layer_1[3621] & layer_1[3557]; 
    assign out[3880] = layer_1[1731] ^ layer_1[1851]; 
    assign out[3881] = ~layer_1[3891] | (layer_1[3846] & layer_1[3891]); 
    assign out[3882] = layer_1[2962]; 
    assign out[3883] = ~(layer_1[972] | layer_1[875]); 
    assign out[3884] = ~(layer_1[1903] ^ layer_1[1840]); 
    assign out[3885] = layer_1[798] & ~layer_1[670]; 
    assign out[3886] = ~(layer_1[3983] | layer_1[3988]); 
    assign out[3887] = ~(layer_1[1210] ^ layer_1[1119]); 
    assign out[3888] = layer_1[2204] & ~layer_1[2142]; 
    assign out[3889] = ~(layer_1[2051] & layer_1[2111]); 
    assign out[3890] = ~layer_1[2280] | (layer_1[2280] & layer_1[2398]); 
    assign out[3891] = ~layer_1[1515]; 
    assign out[3892] = layer_1[323] & ~layer_1[414]; 
    assign out[3893] = ~layer_1[838]; 
    assign out[3894] = layer_1[2555] ^ layer_1[2523]; 
    assign out[3895] = ~(layer_1[2071] | layer_1[2040]); 
    assign out[3896] = layer_1[3244]; 
    assign out[3897] = layer_1[691]; 
    assign out[3898] = ~layer_1[2182] | (layer_1[2182] & layer_1[2295]); 
    assign out[3899] = ~layer_1[3137] | (layer_1[3137] & layer_1[3112]); 
    assign out[3900] = layer_1[2230] & ~layer_1[2118]; 
    assign out[3901] = ~layer_1[3242]; 
    assign out[3902] = ~(layer_1[2699] ^ layer_1[2728]); 
    assign out[3903] = ~(layer_1[1491] ^ layer_1[1412]); 
    assign out[3904] = layer_1[1260] & ~layer_1[1183]; 
    assign out[3905] = layer_1[2732]; 
    assign out[3906] = layer_1[2175] | layer_1[2290]; 
    assign out[3907] = layer_1[2190]; 
    assign out[3908] = ~layer_1[692]; 
    assign out[3909] = layer_1[2138]; 
    assign out[3910] = layer_1[3546] & ~layer_1[3577]; 
    assign out[3911] = layer_1[2879]; 
    assign out[3912] = ~(layer_1[429] | layer_1[419]); 
    assign out[3913] = ~layer_1[981]; 
    assign out[3914] = ~layer_1[2188]; 
    assign out[3915] = layer_1[1750] & ~layer_1[1710]; 
    assign out[3916] = layer_1[2297]; 
    assign out[3917] = layer_1[2451] & ~layer_1[2387]; 
    assign out[3918] = layer_1[39]; 
    assign out[3919] = layer_1[1547] & ~layer_1[1609]; 
    assign out[3920] = layer_1[3184] & ~layer_1[3071]; 
    assign out[3921] = layer_1[3252] & layer_1[3268]; 
    assign out[3922] = layer_1[2993] & layer_1[3013]; 
    assign out[3923] = ~(layer_1[1372] ^ layer_1[1471]); 
    assign out[3924] = layer_1[2751] | layer_1[2641]; 
    assign out[3925] = ~layer_1[606]; 
    assign out[3926] = layer_1[583] & ~layer_1[551]; 
    assign out[3927] = layer_1[3325]; 
    assign out[3928] = layer_1[644] & ~layer_1[757]; 
    assign out[3929] = ~layer_1[1223]; 
    assign out[3930] = ~(layer_1[1899] | layer_1[1812]); 
    assign out[3931] = ~(layer_1[820] ^ layer_1[871]); 
    assign out[3932] = ~(layer_1[3503] | layer_1[3449]); 
    assign out[3933] = layer_1[1921] ^ layer_1[1898]; 
    assign out[3934] = layer_1[1558]; 
    assign out[3935] = layer_1[2509] ^ layer_1[2404]; 
    assign out[3936] = layer_1[3280] & ~layer_1[3347]; 
    assign out[3937] = layer_1[2662] & layer_1[2729]; 
    assign out[3938] = ~(layer_1[2259] ^ layer_1[2333]); 
    assign out[3939] = ~layer_1[1722]; 
    assign out[3940] = ~layer_1[592]; 
    assign out[3941] = layer_1[3843] & ~layer_1[3919]; 
    assign out[3942] = ~(layer_1[282] ^ layer_1[273]); 
    assign out[3943] = layer_1[4] & ~layer_1[50]; 
    assign out[3944] = layer_1[807]; 
    assign out[3945] = ~(layer_1[2519] | layer_1[2413]); 
    assign out[3946] = ~(layer_1[1527] & layer_1[1464]); 
    assign out[3947] = ~layer_1[1017]; 
    assign out[3948] = layer_1[918] ^ layer_1[890]; 
    assign out[3949] = layer_1[880] ^ layer_1[994]; 
    assign out[3950] = layer_1[3348]; 
    assign out[3951] = ~(layer_1[541] | layer_1[557]); 
    assign out[3952] = ~(layer_1[3395] ^ layer_1[3347]); 
    assign out[3953] = ~(layer_1[1393] ^ layer_1[1341]); 
    assign out[3954] = ~layer_1[3614]; 
    assign out[3955] = layer_1[65]; 
    assign out[3956] = layer_1[1384]; 
    assign out[3957] = ~layer_1[2600]; 
    assign out[3958] = layer_1[3173] & ~layer_1[3095]; 
    assign out[3959] = layer_1[1504]; 
    assign out[3960] = layer_1[1936] & ~layer_1[1946]; 
    assign out[3961] = layer_1[1571] & layer_1[1639]; 
    assign out[3962] = layer_1[153] & ~layer_1[276]; 
    assign out[3963] = ~layer_1[3137]; 
    assign out[3964] = layer_1[2072] & ~layer_1[2166]; 
    assign out[3965] = layer_1[3738]; 
    assign out[3966] = layer_1[1214] & ~layer_1[1192]; 
    assign out[3967] = layer_1[1631]; 
    assign out[3968] = layer_1[1115] & ~layer_1[1004]; 
    assign out[3969] = ~(layer_1[1774] | layer_1[1721]); 
    assign out[3970] = ~(layer_1[1315] ^ layer_1[1233]); 
    assign out[3971] = ~(layer_1[2760] ^ layer_1[2807]); 
    assign out[3972] = ~(layer_1[1055] | layer_1[1155]); 
    assign out[3973] = ~layer_1[190] | (layer_1[316] & layer_1[190]); 
    assign out[3974] = layer_1[1117] ^ layer_1[1076]; 
    assign out[3975] = layer_1[2701] & layer_1[2711]; 
    assign out[3976] = layer_1[2409]; 
    assign out[3977] = layer_1[3027] & layer_1[3045]; 
    assign out[3978] = ~layer_1[434]; 
    assign out[3979] = layer_1[1193]; 
    assign out[3980] = layer_1[3511]; 
    assign out[3981] = layer_1[506]; 
    assign out[3982] = layer_1[1881]; 
    assign out[3983] = ~layer_1[3539]; 
    assign out[3984] = ~(layer_1[3270] | layer_1[3243]); 
    assign out[3985] = layer_1[1098] ^ layer_1[1047]; 
    assign out[3986] = layer_1[3702] & ~layer_1[3732]; 
    assign out[3987] = ~(layer_1[904] | layer_1[1004]); 
    assign out[3988] = layer_1[545] & ~layer_1[522]; 
    assign out[3989] = layer_1[2262]; 
    assign out[3990] = layer_1[111]; 
    assign out[3991] = ~layer_1[3266] | (layer_1[3391] & layer_1[3266]); 
    assign out[3992] = layer_1[718] & ~layer_1[720]; 
    assign out[3993] = layer_1[2802]; 
    assign out[3994] = ~(layer_1[2109] | layer_1[2162]); 
    assign out[3995] = layer_1[2705] & ~layer_1[2715]; 
    assign out[3996] = ~(layer_1[1517] | layer_1[1420]); 
    assign out[3997] = ~(layer_1[2193] | layer_1[2098]); 
    assign out[3998] = layer_1[1672] & layer_1[1548]; 
    assign out[3999] = ~(layer_1[3273] ^ layer_1[3165]); 

endmodule
