// Generated from: test_and_d16r1_8x256_256i_256o.npz
module net (
    input wire  [255:0] in,
    output wire [255:0] out
);
    wire [256:0] layer_0;
    wire [256:0] layer_1;
    wire [256:0] layer_2;
    wire [256:0] layer_3;
    wire [256:0] layer_4;
    wire [256:0] layer_5;
    wire [256:0] layer_6;

    // Layer 0 ============================================================
    assign layer_0[0] = in[7] & in[3]; 
    assign layer_0[1] = in[10] & in[2]; 
    assign layer_0[2] = in[4] & in[8]; 
    assign layer_0[3] = in[11] & in[14]; 
    assign layer_0[4] = in[5] & in[9]; 
    assign layer_0[5] = in[8] & in[14]; 
    assign layer_0[6] = in[15] & in[17]; 
    assign layer_0[7] = in[18] & in[5]; 
    assign layer_0[8] = in[15] & in[12]; 
    assign layer_0[9] = in[19] & in[11]; 
    assign layer_0[10] = in[1] & in[23]; 
    assign layer_0[11] = in[17] & in[23]; 
    assign layer_0[12] = in[0] & in[18]; 
    assign layer_0[13] = in[21] & in[1]; 
    assign layer_0[14] = in[28] & in[26]; 
    assign layer_0[15] = in[12] & in[22]; 
    assign layer_0[16] = in[10] & in[8]; 
    assign layer_0[17] = in[31] & in[7]; 
    assign layer_0[18] = in[32] & in[25]; 
    assign layer_0[19] = in[17] & in[29]; 
    assign layer_0[20] = in[7] & in[25]; 
    assign layer_0[21] = in[31] & in[28]; 
    assign layer_0[22] = in[16] & in[15]; 
    assign layer_0[23] = in[29] & in[15]; 
    assign layer_0[24] = in[39] & in[24]; 
    assign layer_0[25] = in[34] & in[12]; 
    assign layer_0[26] = in[40] & in[29]; 
    assign layer_0[27] = in[39] & in[41]; 
    assign layer_0[28] = in[25] & in[33]; 
    assign layer_0[29] = in[36] & in[33]; 
    assign layer_0[30] = in[42] & in[16]; 
    assign layer_0[31] = in[37] & in[39]; 
    assign layer_0[32] = in[19] & in[19]; 
    assign layer_0[33] = in[37] & in[31]; 
    assign layer_0[34] = in[45] & in[42]; 
    assign layer_0[35] = in[41] & in[18]; 
    assign layer_0[36] = in[26] & in[48]; 
    assign layer_0[37] = in[53] & in[35]; 
    assign layer_0[38] = in[32] & in[53]; 
    assign layer_0[39] = in[53] & in[30]; 
    assign layer_0[40] = in[51] & in[54]; 
    assign layer_0[41] = in[31] & in[27]; 
    assign layer_0[42] = in[52] & in[35]; 
    assign layer_0[43] = in[43] & in[37]; 
    assign layer_0[44] = in[33] & in[39]; 
    assign layer_0[45] = in[61] & in[47]; 
    assign layer_0[46] = in[49] & in[61]; 
    assign layer_0[47] = in[47] & in[48]; 
    assign layer_0[48] = in[47] & in[34]; 
    assign layer_0[49] = in[61] & in[44]; 
    assign layer_0[50] = in[42] & in[65]; 
    assign layer_0[51] = in[37] & in[60]; 
    assign layer_0[52] = in[58] & in[36]; 
    assign layer_0[53] = in[69] & in[59]; 
    assign layer_0[54] = in[45] & in[45]; 
    assign layer_0[55] = in[58] & in[50]; 
    assign layer_0[56] = in[71] & in[66]; 
    assign layer_0[57] = in[44] & in[45]; 
    assign layer_0[58] = in[55] & in[72]; 
    assign layer_0[59] = in[60] & in[49]; 
    assign layer_0[60] = in[52] & in[60]; 
    assign layer_0[61] = in[58] & in[50]; 
    assign layer_0[62] = in[47] & in[65]; 
    assign layer_0[63] = in[74] & in[50]; 
    assign layer_0[64] = in[58] & in[57]; 
    assign layer_0[65] = in[66] & in[54]; 
    assign layer_0[66] = in[61] & in[60]; 
    assign layer_0[67] = in[72] & in[54]; 
    assign layer_0[68] = in[57] & in[68]; 
    assign layer_0[69] = in[75] & in[53]; 
    assign layer_0[70] = in[62] & in[80]; 
    assign layer_0[71] = in[76] & in[70]; 
    assign layer_0[72] = in[84] & in[55]; 
    assign layer_0[73] = in[58] & in[75]; 
    assign layer_0[74] = in[74] & in[65]; 
    assign layer_0[75] = in[74] & in[90]; 
    assign layer_0[76] = in[79] & in[60]; 
    assign layer_0[77] = in[77] & in[84]; 
    assign layer_0[78] = in[72] & in[70]; 
    assign layer_0[79] = in[72] & in[81]; 
    assign layer_0[80] = in[66] & in[90]; 
    assign layer_0[81] = in[88] & in[81]; 
    assign layer_0[82] = in[82] & in[82]; 
    assign layer_0[83] = in[91] & in[81]; 
    assign layer_0[84] = in[90] & in[69]; 
    assign layer_0[85] = in[75] & in[93]; 
    assign layer_0[86] = in[83] & in[94]; 
    assign layer_0[87] = in[84] & in[98]; 
    assign layer_0[88] = in[84] & in[96]; 
    assign layer_0[89] = in[73] & in[81]; 
    assign layer_0[90] = in[103] & in[92]; 
    assign layer_0[91] = in[104] & in[85]; 
    assign layer_0[92] = in[91] & in[103]; 
    assign layer_0[93] = in[102] & in[80]; 
    assign layer_0[94] = in[106] & in[89]; 
    assign layer_0[95] = in[105] & in[102]; 
    assign layer_0[96] = in[83] & in[111]; 
    assign layer_0[97] = in[104] & in[86]; 
    assign layer_0[98] = in[104] & in[94]; 
    assign layer_0[99] = in[105] & in[114]; 
    assign layer_0[100] = in[112] & in[115]; 
    assign layer_0[101] = in[109] & in[102]; 
    assign layer_0[102] = in[109] & in[92]; 
    assign layer_0[103] = in[98] & in[117]; 
    assign layer_0[104] = in[93] & in[92]; 
    assign layer_0[105] = in[118] & in[110]; 
    assign layer_0[106] = in[115] & in[108]; 
    assign layer_0[107] = in[104] & in[122]; 
    assign layer_0[108] = in[98] & in[115]; 
    assign layer_0[109] = in[98] & in[124]; 
    assign layer_0[110] = in[123] & in[111]; 
    assign layer_0[111] = in[98] & in[126]; 
    assign layer_0[112] = in[102] & in[110]; 
    assign layer_0[113] = in[104] & in[125]; 
    assign layer_0[114] = in[102] & in[125]; 
    assign layer_0[115] = in[122] & in[129]; 
    assign layer_0[116] = in[115] & in[129]; 
    assign layer_0[117] = in[115] & in[104]; 
    assign layer_0[118] = in[132] & in[104]; 
    assign layer_0[119] = in[121] & in[129]; 
    assign layer_0[120] = in[119] & in[127]; 
    assign layer_0[121] = in[105] & in[131]; 
    assign layer_0[122] = in[120] & in[117]; 
    assign layer_0[123] = in[127] & in[134]; 
    assign layer_0[124] = in[121] & in[112]; 
    assign layer_0[125] = in[138] & in[135]; 
    assign layer_0[126] = in[113] & in[111]; 
    assign layer_0[127] = in[122] & in[129]; 
    assign layer_0[128] = in[114] & in[140]; 
    assign layer_0[129] = in[122] & in[118]; 
    assign layer_0[130] = in[132] & in[122]; 
    assign layer_0[131] = in[127] & in[121]; 
    assign layer_0[132] = in[130] & in[124]; 
    assign layer_0[133] = in[125] & in[146]; 
    assign layer_0[134] = in[146] & in[141]; 
    assign layer_0[135] = in[140] & in[143]; 
    assign layer_0[136] = in[135] & in[149]; 
    assign layer_0[137] = in[142] & in[144]; 
    assign layer_0[138] = in[131] & in[130]; 
    assign layer_0[139] = in[140] & in[144]; 
    assign layer_0[140] = in[152] & in[135]; 
    assign layer_0[141] = in[127] & in[126]; 
    assign layer_0[142] = in[152] & in[137]; 
    assign layer_0[143] = in[144] & in[135]; 
    assign layer_0[144] = in[134] & in[137]; 
    assign layer_0[145] = in[155] & in[154]; 
    assign layer_0[146] = in[156] & in[144]; 
    assign layer_0[147] = in[161] & in[160]; 
    assign layer_0[148] = in[135] & in[133]; 
    assign layer_0[149] = in[155] & in[137]; 
    assign layer_0[150] = in[140] & in[151]; 
    assign layer_0[151] = in[159] & in[158]; 
    assign layer_0[152] = in[158] & in[137]; 
    assign layer_0[153] = in[139] & in[159]; 
    assign layer_0[154] = in[138] & in[155]; 
    assign layer_0[155] = in[167] & in[141]; 
    assign layer_0[156] = in[159] & in[160]; 
    assign layer_0[157] = in[153] & in[151]; 
    assign layer_0[158] = in[170] & in[159]; 
    assign layer_0[159] = in[170] & in[160]; 
    assign layer_0[160] = in[144] & in[157]; 
    assign layer_0[161] = in[175] & in[153]; 
    assign layer_0[162] = in[167] & in[167]; 
    assign layer_0[163] = in[176] & in[148]; 
    assign layer_0[164] = in[178] & in[179]; 
    assign layer_0[165] = in[171] & in[163]; 
    assign layer_0[166] = in[177] & in[149]; 
    assign layer_0[167] = in[161] & in[169]; 
    assign layer_0[168] = in[154] & in[169]; 
    assign layer_0[169] = in[153] & in[155]; 
    assign layer_0[170] = in[171] & in[184]; 
    assign layer_0[171] = in[171] & in[170]; 
    assign layer_0[172] = in[165] & in[172]; 
    assign layer_0[173] = in[157] & in[179]; 
    assign layer_0[174] = in[179] & in[188]; 
    assign layer_0[175] = in[177] & in[177]; 
    assign layer_0[176] = in[189] & in[172]; 
    assign layer_0[177] = in[191] & in[170]; 
    assign layer_0[178] = in[168] & in[192]; 
    assign layer_0[179] = in[179] & in[188]; 
    assign layer_0[180] = in[183] & in[188]; 
    assign layer_0[181] = in[193] & in[169]; 
    assign layer_0[182] = in[169] & in[171]; 
    assign layer_0[183] = in[186] & in[170]; 
    assign layer_0[184] = in[200] & in[181]; 
    assign layer_0[185] = in[173] & in[184]; 
    assign layer_0[186] = in[172] & in[188]; 
    assign layer_0[187] = in[191] & in[178]; 
    assign layer_0[188] = in[190] & in[177]; 
    assign layer_0[189] = in[202] & in[185]; 
    assign layer_0[190] = in[198] & in[179]; 
    assign layer_0[191] = in[200] & in[193]; 
    assign layer_0[192] = in[197] & in[193]; 
    assign layer_0[193] = in[183] & in[192]; 
    assign layer_0[194] = in[209] & in[204]; 
    assign layer_0[195] = in[186] & in[188]; 
    assign layer_0[196] = in[210] & in[192]; 
    assign layer_0[197] = in[182] & in[184]; 
    assign layer_0[198] = in[205] & in[202]; 
    assign layer_0[199] = in[183] & in[198]; 
    assign layer_0[200] = in[188] & in[188]; 
    assign layer_0[201] = in[213] & in[210]; 
    assign layer_0[202] = in[213] & in[211]; 
    assign layer_0[203] = in[191] & in[208]; 
    assign layer_0[204] = in[212] & in[212]; 
    assign layer_0[205] = in[205] & in[191]; 
    assign layer_0[206] = in[218] & in[213]; 
    assign layer_0[207] = in[212] & in[201]; 
    assign layer_0[208] = in[206] & in[215]; 
    assign layer_0[209] = in[207] & in[218]; 
    assign layer_0[210] = in[202] & in[216]; 
    assign layer_0[211] = in[207] & in[200]; 
    assign layer_0[212] = in[209] & in[198]; 
    assign layer_0[213] = in[213] & in[223]; 
    assign layer_0[214] = in[217] & in[213]; 
    assign layer_0[215] = in[209] & in[208]; 
    assign layer_0[216] = in[206] & in[209]; 
    assign layer_0[217] = in[225] & in[232]; 
    assign layer_0[218] = in[224] & in[219]; 
    assign layer_0[219] = in[229] & in[219]; 
    assign layer_0[220] = in[235] & in[211]; 
    assign layer_0[221] = in[231] & in[219]; 
    assign layer_0[222] = in[232] & in[208]; 
    assign layer_0[223] = in[213] & in[222]; 
    assign layer_0[224] = in[208] & in[232]; 
    assign layer_0[225] = in[225] & in[212]; 
    assign layer_0[226] = in[214] & in[232]; 
    assign layer_0[227] = in[215] & in[238]; 
    assign layer_0[228] = in[235] & in[219]; 
    assign layer_0[229] = in[232] & in[231]; 
    assign layer_0[230] = in[216] & in[236]; 
    assign layer_0[231] = in[224] & in[224]; 
    assign layer_0[232] = in[247] & in[236]; 
    assign layer_0[233] = in[220] & in[230]; 
    assign layer_0[234] = in[218] & in[238]; 
    assign layer_0[235] = in[245] & in[233]; 
    assign layer_0[236] = in[236] & in[247]; 
    assign layer_0[237] = in[246] & in[249]; 
    assign layer_0[238] = in[231] & in[252]; 
    assign layer_0[239] = in[239] & in[251]; 
    assign layer_0[240] = in[232] & in[255]; 
    assign layer_0[241] = in[233] & in[225]; 
    assign layer_0[242] = in[237] & in[229]; 
    assign layer_0[243] = in[233] & in[249]; 
    assign layer_0[244] = in[249] & in[253]; 
    assign layer_0[245] = in[237] & in[230]; 
    assign layer_0[246] = in[231] & in[250]; 
    assign layer_0[247] = in[250] & in[248]; 
    assign layer_0[248] = in[232] & in[232]; 
    assign layer_0[249] = in[240] & in[255]; 
    assign layer_0[250] = in[234] & in[239]; 
    assign layer_0[251] = in[250] & in[245]; 
    assign layer_0[252] = in[253] & in[245]; 
    assign layer_0[253] = in[251] & in[245]; 
    assign layer_0[254] = in[246] & in[255]; 
    assign layer_0[255] = in[254] & in[244]; 
    // Layer 1 ============================================================
    assign layer_1[0] = layer_0[8] & layer_0[13]; 
    assign layer_1[1] = layer_0[14] & layer_0[5]; 
    assign layer_1[2] = layer_0[1] & layer_0[15]; 
    assign layer_1[3] = layer_0[3] & layer_0[9]; 
    assign layer_1[4] = layer_0[6] & layer_0[16]; 
    assign layer_1[5] = layer_0[8] & layer_0[0]; 
    assign layer_1[6] = layer_0[19] & layer_0[2]; 
    assign layer_1[7] = layer_0[16] & layer_0[9]; 
    assign layer_1[8] = layer_0[11] & layer_0[23]; 
    assign layer_1[9] = layer_0[11] & layer_0[9]; 
    assign layer_1[10] = layer_0[13] & layer_0[25]; 
    assign layer_1[11] = layer_0[16] & layer_0[26]; 
    assign layer_1[12] = layer_0[7] & layer_0[22]; 
    assign layer_1[13] = layer_0[0] & layer_0[6]; 
    assign layer_1[14] = layer_0[2] & layer_0[10]; 
    assign layer_1[15] = layer_0[13] & layer_0[0]; 
    assign layer_1[16] = layer_0[9] & layer_0[11]; 
    assign layer_1[17] = layer_0[16] & layer_0[9]; 
    assign layer_1[18] = layer_0[6] & layer_0[3]; 
    assign layer_1[19] = layer_0[22] & layer_0[14]; 
    assign layer_1[20] = layer_0[14] & layer_0[34]; 
    assign layer_1[21] = layer_0[37] & layer_0[5]; 
    assign layer_1[22] = layer_0[32] & layer_0[35]; 
    assign layer_1[23] = layer_0[35] & layer_0[25]; 
    assign layer_1[24] = layer_0[20] & layer_0[26]; 
    assign layer_1[25] = layer_0[35] & layer_0[23]; 
    assign layer_1[26] = layer_0[39] & layer_0[24]; 
    assign layer_1[27] = layer_0[17] & layer_0[42]; 
    assign layer_1[28] = layer_0[18] & layer_0[32]; 
    assign layer_1[29] = layer_0[24] & layer_0[22]; 
    assign layer_1[30] = layer_0[32] & layer_0[43]; 
    assign layer_1[31] = layer_0[28] & layer_0[45]; 
    assign layer_1[32] = layer_0[21] & layer_0[34]; 
    assign layer_1[33] = layer_0[21] & layer_0[48]; 
    assign layer_1[34] = layer_0[50] & layer_0[24]; 
    assign layer_1[35] = layer_0[47] & layer_0[37]; 
    assign layer_1[36] = layer_0[50] & layer_0[43]; 
    assign layer_1[37] = layer_0[32] & layer_0[29]; 
    assign layer_1[38] = layer_0[31] & layer_0[29]; 
    assign layer_1[39] = layer_0[51] & layer_0[38]; 
    assign layer_1[40] = layer_0[37] & layer_0[51]; 
    assign layer_1[41] = layer_0[55] & layer_0[40]; 
    assign layer_1[42] = layer_0[45] & layer_0[56]; 
    assign layer_1[43] = layer_0[40] & layer_0[36]; 
    assign layer_1[44] = layer_0[47] & layer_0[47]; 
    assign layer_1[45] = layer_0[60] & layer_0[53]; 
    assign layer_1[46] = layer_0[57] & layer_0[49]; 
    assign layer_1[47] = layer_0[56] & layer_0[47]; 
    assign layer_1[48] = layer_0[62] & layer_0[40]; 
    assign layer_1[49] = layer_0[44] & layer_0[62]; 
    assign layer_1[50] = layer_0[39] & layer_0[62]; 
    assign layer_1[51] = layer_0[65] & layer_0[56]; 
    assign layer_1[52] = layer_0[38] & layer_0[42]; 
    assign layer_1[53] = layer_0[62] & layer_0[44]; 
    assign layer_1[54] = layer_0[44] & layer_0[62]; 
    assign layer_1[55] = layer_0[51] & layer_0[58]; 
    assign layer_1[56] = layer_0[47] & layer_0[60]; 
    assign layer_1[57] = layer_0[59] & layer_0[61]; 
    assign layer_1[58] = layer_0[43] & layer_0[68]; 
    assign layer_1[59] = layer_0[61] & layer_0[54]; 
    assign layer_1[60] = layer_0[62] & layer_0[62]; 
    assign layer_1[61] = layer_0[58] & layer_0[60]; 
    assign layer_1[62] = layer_0[71] & layer_0[55]; 
    assign layer_1[63] = layer_0[57] & layer_0[50]; 
    assign layer_1[64] = layer_0[57] & layer_0[68]; 
    assign layer_1[65] = layer_0[60] & layer_0[49]; 
    assign layer_1[66] = layer_0[64] & layer_0[81]; 
    assign layer_1[67] = layer_0[71] & layer_0[72]; 
    assign layer_1[68] = layer_0[63] & layer_0[76]; 
    assign layer_1[69] = layer_0[53] & layer_0[65]; 
    assign layer_1[70] = layer_0[82] & layer_0[56]; 
    assign layer_1[71] = layer_0[71] & layer_0[71]; 
    assign layer_1[72] = layer_0[58] & layer_0[58]; 
    assign layer_1[73] = layer_0[68] & layer_0[62]; 
    assign layer_1[74] = layer_0[86] & layer_0[72]; 
    assign layer_1[75] = layer_0[72] & layer_0[73]; 
    assign layer_1[76] = layer_0[80] & layer_0[88]; 
    assign layer_1[77] = layer_0[63] & layer_0[84]; 
    assign layer_1[78] = layer_0[67] & layer_0[63]; 
    assign layer_1[79] = layer_0[64] & layer_0[69]; 
    assign layer_1[80] = layer_0[66] & layer_0[83]; 
    assign layer_1[81] = layer_0[97] & layer_0[67]; 
    assign layer_1[82] = layer_0[74] & layer_0[69]; 
    assign layer_1[83] = layer_0[87] & layer_0[94]; 
    assign layer_1[84] = layer_0[76] & layer_0[82]; 
    assign layer_1[85] = layer_0[83] & layer_0[94]; 
    assign layer_1[86] = layer_0[77] & layer_0[88]; 
    assign layer_1[87] = layer_0[82] & layer_0[73]; 
    assign layer_1[88] = layer_0[92] & layer_0[96]; 
    assign layer_1[89] = layer_0[73] & layer_0[98]; 
    assign layer_1[90] = layer_0[92] & layer_0[84]; 
    assign layer_1[91] = layer_0[101] & layer_0[76]; 
    assign layer_1[92] = layer_0[83] & layer_0[77]; 
    assign layer_1[93] = layer_0[84] & layer_0[88]; 
    assign layer_1[94] = layer_0[95] & layer_0[109]; 
    assign layer_1[95] = layer_0[91] & layer_0[78]; 
    assign layer_1[96] = layer_0[99] & layer_0[108]; 
    assign layer_1[97] = layer_0[94] & layer_0[93]; 
    assign layer_1[98] = layer_0[84] & layer_0[98]; 
    assign layer_1[99] = layer_0[100] & layer_0[91]; 
    assign layer_1[100] = layer_0[111] & layer_0[104]; 
    assign layer_1[101] = layer_0[108] & layer_0[112]; 
    assign layer_1[102] = layer_0[93] & layer_0[108]; 
    assign layer_1[103] = layer_0[89] & layer_0[99]; 
    assign layer_1[104] = layer_0[115] & layer_0[90]; 
    assign layer_1[105] = layer_0[91] & layer_0[104]; 
    assign layer_1[106] = layer_0[101] & layer_0[96]; 
    assign layer_1[107] = layer_0[122] & layer_0[118]; 
    assign layer_1[108] = layer_0[118] & layer_0[98]; 
    assign layer_1[109] = layer_0[118] & layer_0[96]; 
    assign layer_1[110] = layer_0[107] & layer_0[113]; 
    assign layer_1[111] = layer_0[114] & layer_0[106]; 
    assign layer_1[112] = layer_0[118] & layer_0[101]; 
    assign layer_1[113] = layer_0[129] & layer_0[122]; 
    assign layer_1[114] = layer_0[126] & layer_0[102]; 
    assign layer_1[115] = layer_0[128] & layer_0[117]; 
    assign layer_1[116] = layer_0[126] & layer_0[118]; 
    assign layer_1[117] = layer_0[130] & layer_0[119]; 
    assign layer_1[118] = layer_0[111] & layer_0[111]; 
    assign layer_1[119] = layer_0[126] & layer_0[118]; 
    assign layer_1[120] = layer_0[121] & layer_0[105]; 
    assign layer_1[121] = layer_0[116] & layer_0[114]; 
    assign layer_1[122] = layer_0[134] & layer_0[122]; 
    assign layer_1[123] = layer_0[108] & layer_0[135]; 
    assign layer_1[124] = layer_0[130] & layer_0[112]; 
    assign layer_1[125] = layer_0[139] & layer_0[116]; 
    assign layer_1[126] = layer_0[125] & layer_0[113]; 
    assign layer_1[127] = layer_0[141] & layer_0[114]; 
    assign layer_1[128] = layer_0[119] & layer_0[129]; 
    assign layer_1[129] = layer_0[125] & layer_0[136]; 
    assign layer_1[130] = layer_0[137] & layer_0[124]; 
    assign layer_1[131] = layer_0[127] & layer_0[115]; 
    assign layer_1[132] = layer_0[132] & layer_0[128]; 
    assign layer_1[133] = layer_0[143] & layer_0[123]; 
    assign layer_1[134] = layer_0[129] & layer_0[127]; 
    assign layer_1[135] = layer_0[122] & layer_0[131]; 
    assign layer_1[136] = layer_0[138] & layer_0[146]; 
    assign layer_1[137] = layer_0[145] & layer_0[134]; 
    assign layer_1[138] = layer_0[127] & layer_0[132]; 
    assign layer_1[139] = layer_0[145] & layer_0[154]; 
    assign layer_1[140] = layer_0[130] & layer_0[148]; 
    assign layer_1[141] = layer_0[142] & layer_0[150]; 
    assign layer_1[142] = layer_0[154] & layer_0[150]; 
    assign layer_1[143] = layer_0[158] & layer_0[126]; 
    assign layer_1[144] = layer_0[129] & layer_0[143]; 
    assign layer_1[145] = layer_0[151] & layer_0[160]; 
    assign layer_1[146] = layer_0[139] & layer_0[150]; 
    assign layer_1[147] = layer_0[142] & layer_0[162]; 
    assign layer_1[148] = layer_0[141] & layer_0[150]; 
    assign layer_1[149] = layer_0[152] & layer_0[139]; 
    assign layer_1[150] = layer_0[144] & layer_0[158]; 
    assign layer_1[151] = layer_0[154] & layer_0[138]; 
    assign layer_1[152] = layer_0[154] & layer_0[150]; 
    assign layer_1[153] = layer_0[160] & layer_0[136]; 
    assign layer_1[154] = layer_0[148] & layer_0[142]; 
    assign layer_1[155] = layer_0[151] & layer_0[144]; 
    assign layer_1[156] = layer_0[144] & layer_0[144]; 
    assign layer_1[157] = layer_0[172] & layer_0[168]; 
    assign layer_1[158] = layer_0[161] & layer_0[168]; 
    assign layer_1[159] = layer_0[164] & layer_0[174]; 
    assign layer_1[160] = layer_0[160] & layer_0[149]; 
    assign layer_1[161] = layer_0[149] & layer_0[167]; 
    assign layer_1[162] = layer_0[168] & layer_0[167]; 
    assign layer_1[163] = layer_0[157] & layer_0[173]; 
    assign layer_1[164] = layer_0[174] & layer_0[167]; 
    assign layer_1[165] = layer_0[180] & layer_0[175]; 
    assign layer_1[166] = layer_0[172] & layer_0[171]; 
    assign layer_1[167] = layer_0[151] & layer_0[166]; 
    assign layer_1[168] = layer_0[168] & layer_0[152]; 
    assign layer_1[169] = layer_0[169] & layer_0[157]; 
    assign layer_1[170] = layer_0[160] & layer_0[184]; 
    assign layer_1[171] = layer_0[175] & layer_0[185]; 
    assign layer_1[172] = layer_0[160] & layer_0[169]; 
    assign layer_1[173] = layer_0[180] & layer_0[185]; 
    assign layer_1[174] = layer_0[174] & layer_0[159]; 
    assign layer_1[175] = layer_0[168] & layer_0[170]; 
    assign layer_1[176] = layer_0[176] & layer_0[171]; 
    assign layer_1[177] = layer_0[181] & layer_0[182]; 
    assign layer_1[178] = layer_0[168] & layer_0[163]; 
    assign layer_1[179] = layer_0[195] & layer_0[171]; 
    assign layer_1[180] = layer_0[170] & layer_0[165]; 
    assign layer_1[181] = layer_0[192] & layer_0[168]; 
    assign layer_1[182] = layer_0[190] & layer_0[197]; 
    assign layer_1[183] = layer_0[186] & layer_0[179]; 
    assign layer_1[184] = layer_0[183] & layer_0[172]; 
    assign layer_1[185] = layer_0[187] & layer_0[171]; 
    assign layer_1[186] = layer_0[173] & layer_0[188]; 
    assign layer_1[187] = layer_0[171] & layer_0[171]; 
    assign layer_1[188] = layer_0[188] & layer_0[194]; 
    assign layer_1[189] = layer_0[200] & layer_0[202]; 
    assign layer_1[190] = layer_0[197] & layer_0[191]; 
    assign layer_1[191] = layer_0[201] & layer_0[206]; 
    assign layer_1[192] = layer_0[185] & layer_0[176]; 
    assign layer_1[193] = layer_0[189] & layer_0[178]; 
    assign layer_1[194] = layer_0[181] & layer_0[179]; 
    assign layer_1[195] = layer_0[194] & layer_0[208]; 
    assign layer_1[196] = layer_0[208] & layer_0[209]; 
    assign layer_1[197] = layer_0[209] & layer_0[186]; 
    assign layer_1[198] = layer_0[188] & layer_0[202]; 
    assign layer_1[199] = layer_0[213] & layer_0[209]; 
    assign layer_1[200] = layer_0[186] & layer_0[195]; 
    assign layer_1[201] = layer_0[205] & layer_0[192]; 
    assign layer_1[202] = layer_0[189] & layer_0[193]; 
    assign layer_1[203] = layer_0[190] & layer_0[217]; 
    assign layer_1[204] = layer_0[199] & layer_0[215]; 
    assign layer_1[205] = layer_0[195] & layer_0[203]; 
    assign layer_1[206] = layer_0[217] & layer_0[189]; 
    assign layer_1[207] = layer_0[197] & layer_0[205]; 
    assign layer_1[208] = layer_0[218] & layer_0[214]; 
    assign layer_1[209] = layer_0[225] & layer_0[201]; 
    assign layer_1[210] = layer_0[214] & layer_0[206]; 
    assign layer_1[211] = layer_0[203] & layer_0[224]; 
    assign layer_1[212] = layer_0[224] & layer_0[214]; 
    assign layer_1[213] = layer_0[217] & layer_0[203]; 
    assign layer_1[214] = layer_0[200] & layer_0[224]; 
    assign layer_1[215] = layer_0[223] & layer_0[200]; 
    assign layer_1[216] = layer_0[219] & layer_0[214]; 
    assign layer_1[217] = layer_0[212] & layer_0[201]; 
    assign layer_1[218] = layer_0[233] & layer_0[204]; 
    assign layer_1[219] = layer_0[221] & layer_0[221]; 
    assign layer_1[220] = layer_0[222] & layer_0[230]; 
    assign layer_1[221] = layer_0[227] & layer_0[220]; 
    assign layer_1[222] = layer_0[224] & layer_0[209]; 
    assign layer_1[223] = layer_0[214] & layer_0[235]; 
    assign layer_1[224] = layer_0[235] & layer_0[222]; 
    assign layer_1[225] = layer_0[214] & layer_0[216]; 
    assign layer_1[226] = layer_0[218] & layer_0[219]; 
    assign layer_1[227] = layer_0[224] & layer_0[214]; 
    assign layer_1[228] = layer_0[237] & layer_0[240]; 
    assign layer_1[229] = layer_0[216] & layer_0[212]; 
    assign layer_1[230] = layer_0[227] & layer_0[238]; 
    assign layer_1[231] = layer_0[232] & layer_0[214]; 
    assign layer_1[232] = layer_0[248] & layer_0[239]; 
    assign layer_1[233] = layer_0[231] & layer_0[230]; 
    assign layer_1[234] = layer_0[222] & layer_0[224]; 
    assign layer_1[235] = layer_0[251] & layer_0[235]; 
    assign layer_1[236] = layer_0[235] & layer_0[219]; 
    assign layer_1[237] = layer_0[231] & layer_0[220]; 
    assign layer_1[238] = layer_0[229] & layer_0[222]; 
    assign layer_1[239] = layer_0[240] & layer_0[238]; 
    assign layer_1[240] = layer_0[233] & layer_0[240]; 
    assign layer_1[241] = layer_0[231] & layer_0[249]; 
    assign layer_1[242] = layer_0[248] & layer_0[253]; 
    assign layer_1[243] = layer_0[235] & layer_0[244]; 
    assign layer_1[244] = layer_0[228] & layer_0[254]; 
    assign layer_1[245] = layer_0[253] & layer_0[238]; 
    assign layer_1[246] = layer_0[237] & layer_0[235]; 
    assign layer_1[247] = layer_0[252] & layer_0[232]; 
    assign layer_1[248] = layer_0[235] & layer_0[254]; 
    assign layer_1[249] = layer_0[243] & layer_0[253]; 
    assign layer_1[250] = layer_0[251] & layer_0[246]; 
    assign layer_1[251] = layer_0[254] & layer_0[248]; 
    assign layer_1[252] = layer_0[252] & layer_0[251]; 
    assign layer_1[253] = layer_0[249] & layer_0[250]; 
    assign layer_1[254] = layer_0[240] & layer_0[242]; 
    assign layer_1[255] = layer_0[252] & layer_0[241]; 
    // Layer 2 ============================================================
    assign layer_2[0] = layer_1[0] & layer_1[2]; 
    assign layer_2[1] = layer_1[12] & layer_1[1]; 
    assign layer_2[2] = layer_1[14] & layer_1[14]; 
    assign layer_2[3] = layer_1[15] & layer_1[8]; 
    assign layer_2[4] = layer_1[4] & layer_1[6]; 
    assign layer_2[5] = layer_1[2] & layer_1[4]; 
    assign layer_2[6] = layer_1[21] & layer_1[17]; 
    assign layer_2[7] = layer_1[19] & layer_1[3]; 
    assign layer_2[8] = layer_1[10] & layer_1[4]; 
    assign layer_2[9] = layer_1[19] & layer_1[6]; 
    assign layer_2[10] = layer_1[11] & layer_1[4]; 
    assign layer_2[11] = layer_1[18] & layer_1[20]; 
    assign layer_2[12] = layer_1[2] & layer_1[2]; 
    assign layer_2[13] = layer_1[24] & layer_1[4]; 
    assign layer_2[14] = layer_1[17] & layer_1[24]; 
    assign layer_2[15] = layer_1[11] & layer_1[28]; 
    assign layer_2[16] = layer_1[8] & layer_1[1]; 
    assign layer_2[17] = layer_1[15] & layer_1[21]; 
    assign layer_2[18] = layer_1[10] & layer_1[29]; 
    assign layer_2[19] = layer_1[26] & layer_1[22]; 
    assign layer_2[20] = layer_1[6] & layer_1[18]; 
    assign layer_2[21] = layer_1[37] & layer_1[11]; 
    assign layer_2[22] = layer_1[10] & layer_1[36]; 
    assign layer_2[23] = layer_1[13] & layer_1[8]; 
    assign layer_2[24] = layer_1[8] & layer_1[35]; 
    assign layer_2[25] = layer_1[31] & layer_1[8]; 
    assign layer_2[26] = layer_1[25] & layer_1[41]; 
    assign layer_2[27] = layer_1[26] & layer_1[22]; 
    assign layer_2[28] = layer_1[25] & layer_1[31]; 
    assign layer_2[29] = layer_1[21] & layer_1[16]; 
    assign layer_2[30] = layer_1[37] & layer_1[20]; 
    assign layer_2[31] = layer_1[38] & layer_1[25]; 
    assign layer_2[32] = layer_1[28] & layer_1[27]; 
    assign layer_2[33] = layer_1[44] & layer_1[48]; 
    assign layer_2[34] = layer_1[26] & layer_1[20]; 
    assign layer_2[35] = layer_1[19] & layer_1[48]; 
    assign layer_2[36] = layer_1[50] & layer_1[22]; 
    assign layer_2[37] = layer_1[46] & layer_1[37]; 
    assign layer_2[38] = layer_1[53] & layer_1[24]; 
    assign layer_2[39] = layer_1[51] & layer_1[26]; 
    assign layer_2[40] = layer_1[43] & layer_1[51]; 
    assign layer_2[41] = layer_1[48] & layer_1[31]; 
    assign layer_2[42] = layer_1[48] & layer_1[44]; 
    assign layer_2[43] = layer_1[30] & layer_1[40]; 
    assign layer_2[44] = layer_1[38] & layer_1[28]; 
    assign layer_2[45] = layer_1[37] & layer_1[57]; 
    assign layer_2[46] = layer_1[33] & layer_1[60]; 
    assign layer_2[47] = layer_1[46] & layer_1[56]; 
    assign layer_2[48] = layer_1[41] & layer_1[60]; 
    assign layer_2[49] = layer_1[35] & layer_1[54]; 
    assign layer_2[50] = layer_1[52] & layer_1[34]; 
    assign layer_2[51] = layer_1[45] & layer_1[34]; 
    assign layer_2[52] = layer_1[64] & layer_1[64]; 
    assign layer_2[53] = layer_1[56] & layer_1[50]; 
    assign layer_2[54] = layer_1[64] & layer_1[65]; 
    assign layer_2[55] = layer_1[39] & layer_1[41]; 
    assign layer_2[56] = layer_1[63] & layer_1[66]; 
    assign layer_2[57] = layer_1[51] & layer_1[65]; 
    assign layer_2[58] = layer_1[42] & layer_1[44]; 
    assign layer_2[59] = layer_1[73] & layer_1[70]; 
    assign layer_2[60] = layer_1[69] & layer_1[61]; 
    assign layer_2[61] = layer_1[48] & layer_1[66]; 
    assign layer_2[62] = layer_1[48] & layer_1[46]; 
    assign layer_2[63] = layer_1[67] & layer_1[73]; 
    assign layer_2[64] = layer_1[65] & layer_1[58]; 
    assign layer_2[65] = layer_1[63] & layer_1[76]; 
    assign layer_2[66] = layer_1[70] & layer_1[71]; 
    assign layer_2[67] = layer_1[80] & layer_1[53]; 
    assign layer_2[68] = layer_1[56] & layer_1[80]; 
    assign layer_2[69] = layer_1[60] & layer_1[59]; 
    assign layer_2[70] = layer_1[78] & layer_1[61]; 
    assign layer_2[71] = layer_1[77] & layer_1[69]; 
    assign layer_2[72] = layer_1[69] & layer_1[59]; 
    assign layer_2[73] = layer_1[89] & layer_1[88]; 
    assign layer_2[74] = layer_1[84] & layer_1[77]; 
    assign layer_2[75] = layer_1[64] & layer_1[72]; 
    assign layer_2[76] = layer_1[87] & layer_1[80]; 
    assign layer_2[77] = layer_1[69] & layer_1[66]; 
    assign layer_2[78] = layer_1[88] & layer_1[92]; 
    assign layer_2[79] = layer_1[70] & layer_1[63]; 
    assign layer_2[80] = layer_1[91] & layer_1[92]; 
    assign layer_2[81] = layer_1[93] & layer_1[72]; 
    assign layer_2[82] = layer_1[93] & layer_1[82]; 
    assign layer_2[83] = layer_1[68] & layer_1[89]; 
    assign layer_2[84] = layer_1[82] & layer_1[69]; 
    assign layer_2[85] = layer_1[70] & layer_1[92]; 
    assign layer_2[86] = layer_1[102] & layer_1[99]; 
    assign layer_2[87] = layer_1[76] & layer_1[96]; 
    assign layer_2[88] = layer_1[74] & layer_1[90]; 
    assign layer_2[89] = layer_1[103] & layer_1[102]; 
    assign layer_2[90] = layer_1[99] & layer_1[96]; 
    assign layer_2[91] = layer_1[87] & layer_1[95]; 
    assign layer_2[92] = layer_1[77] & layer_1[83]; 
    assign layer_2[93] = layer_1[98] & layer_1[108]; 
    assign layer_2[94] = layer_1[98] & layer_1[87]; 
    assign layer_2[95] = layer_1[110] & layer_1[81]; 
    assign layer_2[96] = layer_1[97] & layer_1[81]; 
    assign layer_2[97] = layer_1[85] & layer_1[88]; 
    assign layer_2[98] = layer_1[112] & layer_1[111]; 
    assign layer_2[99] = layer_1[83] & layer_1[98]; 
    assign layer_2[100] = layer_1[102] & layer_1[97]; 
    assign layer_2[101] = layer_1[106] & layer_1[99]; 
    assign layer_2[102] = layer_1[112] & layer_1[109]; 
    assign layer_2[103] = layer_1[98] & layer_1[116]; 
    assign layer_2[104] = layer_1[113] & layer_1[90]; 
    assign layer_2[105] = layer_1[91] & layer_1[97]; 
    assign layer_2[106] = layer_1[120] & layer_1[89]; 
    assign layer_2[107] = layer_1[115] & layer_1[111]; 
    assign layer_2[108] = layer_1[120] & layer_1[113]; 
    assign layer_2[109] = layer_1[114] & layer_1[117]; 
    assign layer_2[110] = layer_1[120] & layer_1[112]; 
    assign layer_2[111] = layer_1[121] & layer_1[120]; 
    assign layer_2[112] = layer_1[126] & layer_1[127]; 
    assign layer_2[113] = layer_1[111] & layer_1[98]; 
    assign layer_2[114] = layer_1[98] & layer_1[108]; 
    assign layer_2[115] = layer_1[121] & layer_1[119]; 
    assign layer_2[116] = layer_1[114] & layer_1[101]; 
    assign layer_2[117] = layer_1[107] & layer_1[130]; 
    assign layer_2[118] = layer_1[108] & layer_1[108]; 
    assign layer_2[119] = layer_1[104] & layer_1[131]; 
    assign layer_2[120] = layer_1[132] & layer_1[134]; 
    assign layer_2[121] = layer_1[133] & layer_1[116]; 
    assign layer_2[122] = layer_1[119] & layer_1[134]; 
    assign layer_2[123] = layer_1[124] & layer_1[111]; 
    assign layer_2[124] = layer_1[118] & layer_1[126]; 
    assign layer_2[125] = layer_1[124] & layer_1[140]; 
    assign layer_2[126] = layer_1[141] & layer_1[114]; 
    assign layer_2[127] = layer_1[130] & layer_1[142]; 
    assign layer_2[128] = layer_1[140] & layer_1[130]; 
    assign layer_2[129] = layer_1[113] & layer_1[127]; 
    assign layer_2[130] = layer_1[130] & layer_1[123]; 
    assign layer_2[131] = layer_1[139] & layer_1[143]; 
    assign layer_2[132] = layer_1[142] & layer_1[140]; 
    assign layer_2[133] = layer_1[148] & layer_1[148]; 
    assign layer_2[134] = layer_1[119] & layer_1[144]; 
    assign layer_2[135] = layer_1[146] & layer_1[124]; 
    assign layer_2[136] = layer_1[125] & layer_1[149]; 
    assign layer_2[137] = layer_1[129] & layer_1[127]; 
    assign layer_2[138] = layer_1[124] & layer_1[136]; 
    assign layer_2[139] = layer_1[125] & layer_1[146]; 
    assign layer_2[140] = layer_1[124] & layer_1[133]; 
    assign layer_2[141] = layer_1[142] & layer_1[155]; 
    assign layer_2[142] = layer_1[133] & layer_1[133]; 
    assign layer_2[143] = layer_1[155] & layer_1[146]; 
    assign layer_2[144] = layer_1[153] & layer_1[154]; 
    assign layer_2[145] = layer_1[146] & layer_1[131]; 
    assign layer_2[146] = layer_1[134] & layer_1[148]; 
    assign layer_2[147] = layer_1[153] & layer_1[155]; 
    assign layer_2[148] = layer_1[159] & layer_1[145]; 
    assign layer_2[149] = layer_1[148] & layer_1[146]; 
    assign layer_2[150] = layer_1[163] & layer_1[159]; 
    assign layer_2[151] = layer_1[152] & layer_1[144]; 
    assign layer_2[152] = layer_1[138] & layer_1[160]; 
    assign layer_2[153] = layer_1[155] & layer_1[138]; 
    assign layer_2[154] = layer_1[163] & layer_1[152]; 
    assign layer_2[155] = layer_1[151] & layer_1[148]; 
    assign layer_2[156] = layer_1[166] & layer_1[163]; 
    assign layer_2[157] = layer_1[142] & layer_1[145]; 
    assign layer_2[158] = layer_1[142] & layer_1[168]; 
    assign layer_2[159] = layer_1[172] & layer_1[159]; 
    assign layer_2[160] = layer_1[160] & layer_1[165]; 
    assign layer_2[161] = layer_1[156] & layer_1[167]; 
    assign layer_2[162] = layer_1[152] & layer_1[169]; 
    assign layer_2[163] = layer_1[168] & layer_1[156]; 
    assign layer_2[164] = layer_1[167] & layer_1[176]; 
    assign layer_2[165] = layer_1[164] & layer_1[152]; 
    assign layer_2[166] = layer_1[164] & layer_1[178]; 
    assign layer_2[167] = layer_1[177] & layer_1[179]; 
    assign layer_2[168] = layer_1[172] & layer_1[175]; 
    assign layer_2[169] = layer_1[171] & layer_1[165]; 
    assign layer_2[170] = layer_1[155] & layer_1[164]; 
    assign layer_2[171] = layer_1[176] & layer_1[166]; 
    assign layer_2[172] = layer_1[166] & layer_1[183]; 
    assign layer_2[173] = layer_1[189] & layer_1[185]; 
    assign layer_2[174] = layer_1[158] & layer_1[169]; 
    assign layer_2[175] = layer_1[164] & layer_1[183]; 
    assign layer_2[176] = layer_1[167] & layer_1[184]; 
    assign layer_2[177] = layer_1[183] & layer_1[163]; 
    assign layer_2[178] = layer_1[166] & layer_1[182]; 
    assign layer_2[179] = layer_1[187] & layer_1[182]; 
    assign layer_2[180] = layer_1[195] & layer_1[191]; 
    assign layer_2[181] = layer_1[174] & layer_1[170]; 
    assign layer_2[182] = layer_1[192] & layer_1[170]; 
    assign layer_2[183] = layer_1[176] & layer_1[192]; 
    assign layer_2[184] = layer_1[181] & layer_1[185]; 
    assign layer_2[185] = layer_1[176] & layer_1[188]; 
    assign layer_2[186] = layer_1[185] & layer_1[189]; 
    assign layer_2[187] = layer_1[184] & layer_1[189]; 
    assign layer_2[188] = layer_1[195] & layer_1[191]; 
    assign layer_2[189] = layer_1[199] & layer_1[172]; 
    assign layer_2[190] = layer_1[177] & layer_1[205]; 
    assign layer_2[191] = layer_1[184] & layer_1[185]; 
    assign layer_2[192] = layer_1[180] & layer_1[182]; 
    assign layer_2[193] = layer_1[183] & layer_1[204]; 
    assign layer_2[194] = layer_1[205] & layer_1[200]; 
    assign layer_2[195] = layer_1[208] & layer_1[204]; 
    assign layer_2[196] = layer_1[193] & layer_1[210]; 
    assign layer_2[197] = layer_1[208] & layer_1[207]; 
    assign layer_2[198] = layer_1[203] & layer_1[202]; 
    assign layer_2[199] = layer_1[214] & layer_1[189]; 
    assign layer_2[200] = layer_1[187] & layer_1[185]; 
    assign layer_2[201] = layer_1[197] & layer_1[198]; 
    assign layer_2[202] = layer_1[186] & layer_1[198]; 
    assign layer_2[203] = layer_1[213] & layer_1[209]; 
    assign layer_2[204] = layer_1[217] & layer_1[192]; 
    assign layer_2[205] = layer_1[220] & layer_1[216]; 
    assign layer_2[206] = layer_1[218] & layer_1[218]; 
    assign layer_2[207] = layer_1[213] & layer_1[190]; 
    assign layer_2[208] = layer_1[223] & layer_1[201]; 
    assign layer_2[209] = layer_1[193] & layer_1[209]; 
    assign layer_2[210] = layer_1[215] & layer_1[216]; 
    assign layer_2[211] = layer_1[221] & layer_1[212]; 
    assign layer_2[212] = layer_1[219] & layer_1[220]; 
    assign layer_2[213] = layer_1[209] & layer_1[210]; 
    assign layer_2[214] = layer_1[209] & layer_1[197]; 
    assign layer_2[215] = layer_1[224] & layer_1[210]; 
    assign layer_2[216] = layer_1[220] & layer_1[226]; 
    assign layer_2[217] = layer_1[227] & layer_1[216]; 
    assign layer_2[218] = layer_1[231] & layer_1[223]; 
    assign layer_2[219] = layer_1[209] & layer_1[230]; 
    assign layer_2[220] = layer_1[218] & layer_1[222]; 
    assign layer_2[221] = layer_1[234] & layer_1[232]; 
    assign layer_2[222] = layer_1[208] & layer_1[212]; 
    assign layer_2[223] = layer_1[207] & layer_1[207]; 
    assign layer_2[224] = layer_1[226] & layer_1[223]; 
    assign layer_2[225] = layer_1[232] & layer_1[223]; 
    assign layer_2[226] = layer_1[241] & layer_1[218]; 
    assign layer_2[227] = layer_1[238] & layer_1[217]; 
    assign layer_2[228] = layer_1[217] & layer_1[237]; 
    assign layer_2[229] = layer_1[220] & layer_1[228]; 
    assign layer_2[230] = layer_1[234] & layer_1[215]; 
    assign layer_2[231] = layer_1[231] & layer_1[242]; 
    assign layer_2[232] = layer_1[234] & layer_1[238]; 
    assign layer_2[233] = layer_1[249] & layer_1[240]; 
    assign layer_2[234] = layer_1[231] & layer_1[240]; 
    assign layer_2[235] = layer_1[244] & layer_1[224]; 
    assign layer_2[236] = layer_1[244] & layer_1[231]; 
    assign layer_2[237] = layer_1[251] & layer_1[241]; 
    assign layer_2[238] = layer_1[228] & layer_1[248]; 
    assign layer_2[239] = layer_1[246] & layer_1[245]; 
    assign layer_2[240] = layer_1[243] & layer_1[252]; 
    assign layer_2[241] = layer_1[225] & layer_1[232]; 
    assign layer_2[242] = layer_1[255] & layer_1[248]; 
    assign layer_2[243] = layer_1[230] & layer_1[248]; 
    assign layer_2[244] = layer_1[254] & layer_1[236]; 
    assign layer_2[245] = layer_1[252] & layer_1[238]; 
    assign layer_2[246] = layer_1[234] & layer_1[243]; 
    assign layer_2[247] = layer_1[242] & layer_1[249]; 
    assign layer_2[248] = layer_1[250] & layer_1[252]; 
    assign layer_2[249] = layer_1[253] & layer_1[246]; 
    assign layer_2[250] = layer_1[250] & layer_1[248]; 
    assign layer_2[251] = layer_1[245] & layer_1[243]; 
    assign layer_2[252] = layer_1[236] & layer_1[237]; 
    assign layer_2[253] = layer_1[249] & layer_1[249]; 
    assign layer_2[254] = layer_1[254] & layer_1[252]; 
    assign layer_2[255] = layer_1[247] & layer_1[249]; 
    // Layer 3 ============================================================
    assign layer_3[0] = layer_2[11] & layer_2[0]; 
    assign layer_3[1] = layer_2[8] & layer_2[1]; 
    assign layer_3[2] = layer_2[12] & layer_2[15]; 
    assign layer_3[3] = layer_2[1] & layer_2[11]; 
    assign layer_3[4] = layer_2[5] & layer_2[1]; 
    assign layer_3[5] = layer_2[11] & layer_2[8]; 
    assign layer_3[6] = layer_2[2] & layer_2[16]; 
    assign layer_3[7] = layer_2[20] & layer_2[8]; 
    assign layer_3[8] = layer_2[20] & layer_2[9]; 
    assign layer_3[9] = layer_2[3] & layer_2[5]; 
    assign layer_3[10] = layer_2[3] & layer_2[21]; 
    assign layer_3[11] = layer_2[23] & layer_2[13]; 
    assign layer_3[12] = layer_2[28] & layer_2[18]; 
    assign layer_3[13] = layer_2[3] & layer_2[6]; 
    assign layer_3[14] = layer_2[4] & layer_2[20]; 
    assign layer_3[15] = layer_2[20] & layer_2[4]; 
    assign layer_3[16] = layer_2[2] & layer_2[15]; 
    assign layer_3[17] = layer_2[1] & layer_2[10]; 
    assign layer_3[18] = layer_2[29] & layer_2[33]; 
    assign layer_3[19] = layer_2[16] & layer_2[31]; 
    assign layer_3[20] = layer_2[33] & layer_2[8]; 
    assign layer_3[21] = layer_2[19] & layer_2[26]; 
    assign layer_3[22] = layer_2[12] & layer_2[18]; 
    assign layer_3[23] = layer_2[36] & layer_2[11]; 
    assign layer_3[24] = layer_2[23] & layer_2[7]; 
    assign layer_3[25] = layer_2[35] & layer_2[21]; 
    assign layer_3[26] = layer_2[11] & layer_2[24]; 
    assign layer_3[27] = layer_2[19] & layer_2[28]; 
    assign layer_3[28] = layer_2[27] & layer_2[23]; 
    assign layer_3[29] = layer_2[43] & layer_2[36]; 
    assign layer_3[30] = layer_2[41] & layer_2[39]; 
    assign layer_3[31] = layer_2[29] & layer_2[34]; 
    assign layer_3[32] = layer_2[42] & layer_2[21]; 
    assign layer_3[33] = layer_2[42] & layer_2[16]; 
    assign layer_3[34] = layer_2[19] & layer_2[47]; 
    assign layer_3[35] = layer_2[49] & layer_2[33]; 
    assign layer_3[36] = layer_2[47] & layer_2[48]; 
    assign layer_3[37] = layer_2[21] & layer_2[30]; 
    assign layer_3[38] = layer_2[47] & layer_2[46]; 
    assign layer_3[39] = layer_2[39] & layer_2[22]; 
    assign layer_3[40] = layer_2[24] & layer_2[51]; 
    assign layer_3[41] = layer_2[39] & layer_2[35]; 
    assign layer_3[42] = layer_2[51] & layer_2[34]; 
    assign layer_3[43] = layer_2[58] & layer_2[56]; 
    assign layer_3[44] = layer_2[34] & layer_2[46]; 
    assign layer_3[45] = layer_2[29] & layer_2[30]; 
    assign layer_3[46] = layer_2[55] & layer_2[57]; 
    assign layer_3[47] = layer_2[44] & layer_2[54]; 
    assign layer_3[48] = layer_2[53] & layer_2[44]; 
    assign layer_3[49] = layer_2[58] & layer_2[36]; 
    assign layer_3[50] = layer_2[48] & layer_2[57]; 
    assign layer_3[51] = layer_2[54] & layer_2[60]; 
    assign layer_3[52] = layer_2[64] & layer_2[54]; 
    assign layer_3[53] = layer_2[61] & layer_2[67]; 
    assign layer_3[54] = layer_2[39] & layer_2[58]; 
    assign layer_3[55] = layer_2[62] & layer_2[54]; 
    assign layer_3[56] = layer_2[60] & layer_2[46]; 
    assign layer_3[57] = layer_2[64] & layer_2[64]; 
    assign layer_3[58] = layer_2[62] & layer_2[42]; 
    assign layer_3[59] = layer_2[50] & layer_2[47]; 
    assign layer_3[60] = layer_2[61] & layer_2[67]; 
    assign layer_3[61] = layer_2[74] & layer_2[68]; 
    assign layer_3[62] = layer_2[70] & layer_2[47]; 
    assign layer_3[63] = layer_2[52] & layer_2[72]; 
    assign layer_3[64] = layer_2[68] & layer_2[72]; 
    assign layer_3[65] = layer_2[64] & layer_2[67]; 
    assign layer_3[66] = layer_2[65] & layer_2[81]; 
    assign layer_3[67] = layer_2[54] & layer_2[63]; 
    assign layer_3[68] = layer_2[64] & layer_2[59]; 
    assign layer_3[69] = layer_2[72] & layer_2[81]; 
    assign layer_3[70] = layer_2[58] & layer_2[85]; 
    assign layer_3[71] = layer_2[59] & layer_2[78]; 
    assign layer_3[72] = layer_2[75] & layer_2[63]; 
    assign layer_3[73] = layer_2[88] & layer_2[86]; 
    assign layer_3[74] = layer_2[76] & layer_2[61]; 
    assign layer_3[75] = layer_2[59] & layer_2[87]; 
    assign layer_3[76] = layer_2[85] & layer_2[66]; 
    assign layer_3[77] = layer_2[83] & layer_2[86]; 
    assign layer_3[78] = layer_2[94] & layer_2[64]; 
    assign layer_3[79] = layer_2[85] & layer_2[83]; 
    assign layer_3[80] = layer_2[81] & layer_2[90]; 
    assign layer_3[81] = layer_2[74] & layer_2[67]; 
    assign layer_3[82] = layer_2[95] & layer_2[83]; 
    assign layer_3[83] = layer_2[87] & layer_2[75]; 
    assign layer_3[84] = layer_2[68] & layer_2[70]; 
    assign layer_3[85] = layer_2[79] & layer_2[75]; 
    assign layer_3[86] = layer_2[82] & layer_2[80]; 
    assign layer_3[87] = layer_2[94] & layer_2[78]; 
    assign layer_3[88] = layer_2[102] & layer_2[102]; 
    assign layer_3[89] = layer_2[94] & layer_2[82]; 
    assign layer_3[90] = layer_2[101] & layer_2[76]; 
    assign layer_3[91] = layer_2[75] & layer_2[94]; 
    assign layer_3[92] = layer_2[95] & layer_2[82]; 
    assign layer_3[93] = layer_2[84] & layer_2[90]; 
    assign layer_3[94] = layer_2[107] & layer_2[84]; 
    assign layer_3[95] = layer_2[80] & layer_2[103]; 
    assign layer_3[96] = layer_2[94] & layer_2[90]; 
    assign layer_3[97] = layer_2[89] & layer_2[107]; 
    assign layer_3[98] = layer_2[82] & layer_2[82]; 
    assign layer_3[99] = layer_2[95] & layer_2[87]; 
    assign layer_3[100] = layer_2[89] & layer_2[86]; 
    assign layer_3[101] = layer_2[91] & layer_2[98]; 
    assign layer_3[102] = layer_2[102] & layer_2[95]; 
    assign layer_3[103] = layer_2[106] & layer_2[95]; 
    assign layer_3[104] = layer_2[118] & layer_2[113]; 
    assign layer_3[105] = layer_2[117] & layer_2[111]; 
    assign layer_3[106] = layer_2[121] & layer_2[115]; 
    assign layer_3[107] = layer_2[91] & layer_2[121]; 
    assign layer_3[108] = layer_2[94] & layer_2[109]; 
    assign layer_3[109] = layer_2[117] & layer_2[119]; 
    assign layer_3[110] = layer_2[118] & layer_2[118]; 
    assign layer_3[111] = layer_2[119] & layer_2[126]; 
    assign layer_3[112] = layer_2[123] & layer_2[106]; 
    assign layer_3[113] = layer_2[122] & layer_2[128]; 
    assign layer_3[114] = layer_2[118] & layer_2[119]; 
    assign layer_3[115] = layer_2[121] & layer_2[107]; 
    assign layer_3[116] = layer_2[112] & layer_2[129]; 
    assign layer_3[117] = layer_2[103] & layer_2[102]; 
    assign layer_3[118] = layer_2[133] & layer_2[128]; 
    assign layer_3[119] = layer_2[132] & layer_2[134]; 
    assign layer_3[120] = layer_2[124] & layer_2[105]; 
    assign layer_3[121] = layer_2[116] & layer_2[117]; 
    assign layer_3[122] = layer_2[127] & layer_2[115]; 
    assign layer_3[123] = layer_2[125] & layer_2[130]; 
    assign layer_3[124] = layer_2[136] & layer_2[114]; 
    assign layer_3[125] = layer_2[134] & layer_2[113]; 
    assign layer_3[126] = layer_2[114] & layer_2[127]; 
    assign layer_3[127] = layer_2[117] & layer_2[119]; 
    assign layer_3[128] = layer_2[142] & layer_2[134]; 
    assign layer_3[129] = layer_2[120] & layer_2[119]; 
    assign layer_3[130] = layer_2[127] & layer_2[124]; 
    assign layer_3[131] = layer_2[146] & layer_2[121]; 
    assign layer_3[132] = layer_2[143] & layer_2[115]; 
    assign layer_3[133] = layer_2[120] & layer_2[134]; 
    assign layer_3[134] = layer_2[127] & layer_2[142]; 
    assign layer_3[135] = layer_2[130] & layer_2[145]; 
    assign layer_3[136] = layer_2[135] & layer_2[136]; 
    assign layer_3[137] = layer_2[127] & layer_2[134]; 
    assign layer_3[138] = layer_2[147] & layer_2[129]; 
    assign layer_3[139] = layer_2[135] & layer_2[123]; 
    assign layer_3[140] = layer_2[139] & layer_2[128]; 
    assign layer_3[141] = layer_2[136] & layer_2[145]; 
    assign layer_3[142] = layer_2[132] & layer_2[150]; 
    assign layer_3[143] = layer_2[138] & layer_2[149]; 
    assign layer_3[144] = layer_2[138] & layer_2[139]; 
    assign layer_3[145] = layer_2[136] & layer_2[146]; 
    assign layer_3[146] = layer_2[144] & layer_2[138]; 
    assign layer_3[147] = layer_2[162] & layer_2[151]; 
    assign layer_3[148] = layer_2[163] & layer_2[162]; 
    assign layer_3[149] = layer_2[141] & layer_2[143]; 
    assign layer_3[150] = layer_2[147] & layer_2[139]; 
    assign layer_3[151] = layer_2[151] & layer_2[159]; 
    assign layer_3[152] = layer_2[142] & layer_2[141]; 
    assign layer_3[153] = layer_2[145] & layer_2[151]; 
    assign layer_3[154] = layer_2[150] & layer_2[160]; 
    assign layer_3[155] = layer_2[157] & layer_2[162]; 
    assign layer_3[156] = layer_2[164] & layer_2[159]; 
    assign layer_3[157] = layer_2[141] & layer_2[164]; 
    assign layer_3[158] = layer_2[165] & layer_2[159]; 
    assign layer_3[159] = layer_2[151] & layer_2[167]; 
    assign layer_3[160] = layer_2[155] & layer_2[159]; 
    assign layer_3[161] = layer_2[150] & layer_2[144]; 
    assign layer_3[162] = layer_2[165] & layer_2[162]; 
    assign layer_3[163] = layer_2[177] & layer_2[173]; 
    assign layer_3[164] = layer_2[175] & layer_2[177]; 
    assign layer_3[165] = layer_2[156] & layer_2[176]; 
    assign layer_3[166] = layer_2[172] & layer_2[150]; 
    assign layer_3[167] = layer_2[154] & layer_2[173]; 
    assign layer_3[168] = layer_2[158] & layer_2[169]; 
    assign layer_3[169] = layer_2[180] & layer_2[153]; 
    assign layer_3[170] = layer_2[185] & layer_2[174]; 
    assign layer_3[171] = layer_2[181] & layer_2[159]; 
    assign layer_3[172] = layer_2[182] & layer_2[183]; 
    assign layer_3[173] = layer_2[159] & layer_2[188]; 
    assign layer_3[174] = layer_2[180] & layer_2[170]; 
    assign layer_3[175] = layer_2[160] & layer_2[163]; 
    assign layer_3[176] = layer_2[183] & layer_2[179]; 
    assign layer_3[177] = layer_2[171] & layer_2[163]; 
    assign layer_3[178] = layer_2[169] & layer_2[186]; 
    assign layer_3[179] = layer_2[165] & layer_2[194]; 
    assign layer_3[180] = layer_2[175] & layer_2[188]; 
    assign layer_3[181] = layer_2[193] & layer_2[178]; 
    assign layer_3[182] = layer_2[171] & layer_2[188]; 
    assign layer_3[183] = layer_2[181] & layer_2[186]; 
    assign layer_3[184] = layer_2[199] & layer_2[187]; 
    assign layer_3[185] = layer_2[177] & layer_2[173]; 
    assign layer_3[186] = layer_2[197] & layer_2[201]; 
    assign layer_3[187] = layer_2[199] & layer_2[183]; 
    assign layer_3[188] = layer_2[203] & layer_2[202]; 
    assign layer_3[189] = layer_2[186] & layer_2[204]; 
    assign layer_3[190] = layer_2[187] & layer_2[189]; 
    assign layer_3[191] = layer_2[199] & layer_2[205]; 
    assign layer_3[192] = layer_2[201] & layer_2[191]; 
    assign layer_3[193] = layer_2[184] & layer_2[194]; 
    assign layer_3[194] = layer_2[197] & layer_2[201]; 
    assign layer_3[195] = layer_2[183] & layer_2[192]; 
    assign layer_3[196] = layer_2[188] & layer_2[186]; 
    assign layer_3[197] = layer_2[185] & layer_2[187]; 
    assign layer_3[198] = layer_2[184] & layer_2[181]; 
    assign layer_3[199] = layer_2[197] & layer_2[203]; 
    assign layer_3[200] = layer_2[191] & layer_2[188]; 
    assign layer_3[201] = layer_2[199] & layer_2[185]; 
    assign layer_3[202] = layer_2[215] & layer_2[214]; 
    assign layer_3[203] = layer_2[218] & layer_2[211]; 
    assign layer_3[204] = layer_2[207] & layer_2[204]; 
    assign layer_3[205] = layer_2[200] & layer_2[204]; 
    assign layer_3[206] = layer_2[218] & layer_2[221]; 
    assign layer_3[207] = layer_2[212] & layer_2[198]; 
    assign layer_3[208] = layer_2[204] & layer_2[223]; 
    assign layer_3[209] = layer_2[219] & layer_2[221]; 
    assign layer_3[210] = layer_2[201] & layer_2[200]; 
    assign layer_3[211] = layer_2[220] & layer_2[207]; 
    assign layer_3[212] = layer_2[208] & layer_2[215]; 
    assign layer_3[213] = layer_2[205] & layer_2[209]; 
    assign layer_3[214] = layer_2[225] & layer_2[204]; 
    assign layer_3[215] = layer_2[221] & layer_2[204]; 
    assign layer_3[216] = layer_2[218] & layer_2[214]; 
    assign layer_3[217] = layer_2[220] & layer_2[219]; 
    assign layer_3[218] = layer_2[234] & layer_2[203]; 
    assign layer_3[219] = layer_2[225] & layer_2[204]; 
    assign layer_3[220] = layer_2[204] & layer_2[235]; 
    assign layer_3[221] = layer_2[220] & layer_2[228]; 
    assign layer_3[222] = layer_2[227] & layer_2[233]; 
    assign layer_3[223] = layer_2[230] & layer_2[211]; 
    assign layer_3[224] = layer_2[229] & layer_2[236]; 
    assign layer_3[225] = layer_2[224] & layer_2[218]; 
    assign layer_3[226] = layer_2[237] & layer_2[221]; 
    assign layer_3[227] = layer_2[236] & layer_2[216]; 
    assign layer_3[228] = layer_2[216] & layer_2[235]; 
    assign layer_3[229] = layer_2[226] & layer_2[243]; 
    assign layer_3[230] = layer_2[235] & layer_2[213]; 
    assign layer_3[231] = layer_2[237] & layer_2[234]; 
    assign layer_3[232] = layer_2[229] & layer_2[218]; 
    assign layer_3[233] = layer_2[240] & layer_2[240]; 
    assign layer_3[234] = layer_2[243] & layer_2[220]; 
    assign layer_3[235] = layer_2[247] & layer_2[240]; 
    assign layer_3[236] = layer_2[223] & layer_2[237]; 
    assign layer_3[237] = layer_2[250] & layer_2[233]; 
    assign layer_3[238] = layer_2[243] & layer_2[228]; 
    assign layer_3[239] = layer_2[232] & layer_2[242]; 
    assign layer_3[240] = layer_2[232] & layer_2[253]; 
    assign layer_3[241] = layer_2[243] & layer_2[245]; 
    assign layer_3[242] = layer_2[248] & layer_2[230]; 
    assign layer_3[243] = layer_2[235] & layer_2[253]; 
    assign layer_3[244] = layer_2[242] & layer_2[245]; 
    assign layer_3[245] = layer_2[241] & layer_2[251]; 
    assign layer_3[246] = layer_2[252] & layer_2[231]; 
    assign layer_3[247] = layer_2[252] & layer_2[240]; 
    assign layer_3[248] = layer_2[251] & layer_2[250]; 
    assign layer_3[249] = layer_2[245] & layer_2[254]; 
    assign layer_3[250] = layer_2[253] & layer_2[251]; 
    assign layer_3[251] = layer_2[254] & layer_2[250]; 
    assign layer_3[252] = layer_2[251] & layer_2[255]; 
    assign layer_3[253] = layer_2[244] & layer_2[243]; 
    assign layer_3[254] = layer_2[240] & layer_2[253]; 
    assign layer_3[255] = layer_2[239] & layer_2[239]; 
    // Layer 4 ============================================================
    assign layer_4[0] = layer_3[11] & layer_3[2]; 
    assign layer_4[1] = layer_3[15] & layer_3[1]; 
    assign layer_4[2] = layer_3[1] & layer_3[11]; 
    assign layer_4[3] = layer_3[4] & layer_3[13]; 
    assign layer_4[4] = layer_3[1] & layer_3[10]; 
    assign layer_4[5] = layer_3[9] & layer_3[12]; 
    assign layer_4[6] = layer_3[3] & layer_3[2]; 
    assign layer_4[7] = layer_3[14] & layer_3[0]; 
    assign layer_4[8] = layer_3[13] & layer_3[3]; 
    assign layer_4[9] = layer_3[21] & layer_3[10]; 
    assign layer_4[10] = layer_3[2] & layer_3[3]; 
    assign layer_4[11] = layer_3[16] & layer_3[1]; 
    assign layer_4[12] = layer_3[7] & layer_3[22]; 
    assign layer_4[13] = layer_3[27] & layer_3[0]; 
    assign layer_4[14] = layer_3[7] & layer_3[12]; 
    assign layer_4[15] = layer_3[15] & layer_3[17]; 
    assign layer_4[16] = layer_3[2] & layer_3[14]; 
    assign layer_4[17] = layer_3[16] & layer_3[8]; 
    assign layer_4[18] = layer_3[3] & layer_3[14]; 
    assign layer_4[19] = layer_3[18] & layer_3[11]; 
    assign layer_4[20] = layer_3[23] & layer_3[16]; 
    assign layer_4[21] = layer_3[8] & layer_3[36]; 
    assign layer_4[22] = layer_3[29] & layer_3[12]; 
    assign layer_4[23] = layer_3[39] & layer_3[36]; 
    assign layer_4[24] = layer_3[30] & layer_3[31]; 
    assign layer_4[25] = layer_3[22] & layer_3[37]; 
    assign layer_4[26] = layer_3[25] & layer_3[18]; 
    assign layer_4[27] = layer_3[17] & layer_3[17]; 
    assign layer_4[28] = layer_3[27] & layer_3[29]; 
    assign layer_4[29] = layer_3[18] & layer_3[40]; 
    assign layer_4[30] = layer_3[38] & layer_3[35]; 
    assign layer_4[31] = layer_3[40] & layer_3[36]; 
    assign layer_4[32] = layer_3[21] & layer_3[24]; 
    assign layer_4[33] = layer_3[48] & layer_3[22]; 
    assign layer_4[34] = layer_3[32] & layer_3[36]; 
    assign layer_4[35] = layer_3[40] & layer_3[30]; 
    assign layer_4[36] = layer_3[33] & layer_3[28]; 
    assign layer_4[37] = layer_3[30] & layer_3[34]; 
    assign layer_4[38] = layer_3[43] & layer_3[24]; 
    assign layer_4[39] = layer_3[54] & layer_3[25]; 
    assign layer_4[40] = layer_3[56] & layer_3[30]; 
    assign layer_4[41] = layer_3[29] & layer_3[34]; 
    assign layer_4[42] = layer_3[43] & layer_3[34]; 
    assign layer_4[43] = layer_3[46] & layer_3[31]; 
    assign layer_4[44] = layer_3[38] & layer_3[31]; 
    assign layer_4[45] = layer_3[51] & layer_3[53]; 
    assign layer_4[46] = layer_3[34] & layer_3[32]; 
    assign layer_4[47] = layer_3[33] & layer_3[58]; 
    assign layer_4[48] = layer_3[61] & layer_3[61]; 
    assign layer_4[49] = layer_3[59] & layer_3[44]; 
    assign layer_4[50] = layer_3[51] & layer_3[34]; 
    assign layer_4[51] = layer_3[65] & layer_3[53]; 
    assign layer_4[52] = layer_3[45] & layer_3[63]; 
    assign layer_4[53] = layer_3[38] & layer_3[58]; 
    assign layer_4[54] = layer_3[67] & layer_3[42]; 
    assign layer_4[55] = layer_3[55] & layer_3[54]; 
    assign layer_4[56] = layer_3[68] & layer_3[49]; 
    assign layer_4[57] = layer_3[43] & layer_3[55]; 
    assign layer_4[58] = layer_3[42] & layer_3[60]; 
    assign layer_4[59] = layer_3[59] & layer_3[60]; 
    assign layer_4[60] = layer_3[44] & layer_3[75]; 
    assign layer_4[61] = layer_3[63] & layer_3[50]; 
    assign layer_4[62] = layer_3[49] & layer_3[69]; 
    assign layer_4[63] = layer_3[64] & layer_3[60]; 
    assign layer_4[64] = layer_3[58] & layer_3[47]; 
    assign layer_4[65] = layer_3[63] & layer_3[51]; 
    assign layer_4[66] = layer_3[60] & layer_3[79]; 
    assign layer_4[67] = layer_3[72] & layer_3[52]; 
    assign layer_4[68] = layer_3[63] & layer_3[57]; 
    assign layer_4[69] = layer_3[65] & layer_3[60]; 
    assign layer_4[70] = layer_3[67] & layer_3[57]; 
    assign layer_4[71] = layer_3[80] & layer_3[83]; 
    assign layer_4[72] = layer_3[57] & layer_3[56]; 
    assign layer_4[73] = layer_3[82] & layer_3[63]; 
    assign layer_4[74] = layer_3[88] & layer_3[71]; 
    assign layer_4[75] = layer_3[62] & layer_3[75]; 
    assign layer_4[76] = layer_3[80] & layer_3[69]; 
    assign layer_4[77] = layer_3[85] & layer_3[68]; 
    assign layer_4[78] = layer_3[70] & layer_3[64]; 
    assign layer_4[79] = layer_3[67] & layer_3[74]; 
    assign layer_4[80] = layer_3[64] & layer_3[79]; 
    assign layer_4[81] = layer_3[75] & layer_3[71]; 
    assign layer_4[82] = layer_3[81] & layer_3[75]; 
    assign layer_4[83] = layer_3[67] & layer_3[67]; 
    assign layer_4[84] = layer_3[95] & layer_3[91]; 
    assign layer_4[85] = layer_3[89] & layer_3[77]; 
    assign layer_4[86] = layer_3[81] & layer_3[83]; 
    assign layer_4[87] = layer_3[100] & layer_3[84]; 
    assign layer_4[88] = layer_3[79] & layer_3[96]; 
    assign layer_4[89] = layer_3[100] & layer_3[103]; 
    assign layer_4[90] = layer_3[93] & layer_3[83]; 
    assign layer_4[91] = layer_3[103] & layer_3[95]; 
    assign layer_4[92] = layer_3[94] & layer_3[97]; 
    assign layer_4[93] = layer_3[102] & layer_3[83]; 
    assign layer_4[94] = layer_3[84] & layer_3[106]; 
    assign layer_4[95] = layer_3[111] & layer_3[98]; 
    assign layer_4[96] = layer_3[90] & layer_3[94]; 
    assign layer_4[97] = layer_3[94] & layer_3[101]; 
    assign layer_4[98] = layer_3[107] & layer_3[82]; 
    assign layer_4[99] = layer_3[101] & layer_3[92]; 
    assign layer_4[100] = layer_3[92] & layer_3[112]; 
    assign layer_4[101] = layer_3[116] & layer_3[111]; 
    assign layer_4[102] = layer_3[101] & layer_3[103]; 
    assign layer_4[103] = layer_3[106] & layer_3[106]; 
    assign layer_4[104] = layer_3[94] & layer_3[108]; 
    assign layer_4[105] = layer_3[118] & layer_3[103]; 
    assign layer_4[106] = layer_3[98] & layer_3[107]; 
    assign layer_4[107] = layer_3[99] & layer_3[106]; 
    assign layer_4[108] = layer_3[110] & layer_3[118]; 
    assign layer_4[109] = layer_3[122] & layer_3[101]; 
    assign layer_4[110] = layer_3[121] & layer_3[102]; 
    assign layer_4[111] = layer_3[114] & layer_3[100]; 
    assign layer_4[112] = layer_3[108] & layer_3[115]; 
    assign layer_4[113] = layer_3[110] & layer_3[97]; 
    assign layer_4[114] = layer_3[114] & layer_3[102]; 
    assign layer_4[115] = layer_3[129] & layer_3[117]; 
    assign layer_4[116] = layer_3[101] & layer_3[128]; 
    assign layer_4[117] = layer_3[126] & layer_3[123]; 
    assign layer_4[118] = layer_3[105] & layer_3[111]; 
    assign layer_4[119] = layer_3[104] & layer_3[117]; 
    assign layer_4[120] = layer_3[125] & layer_3[116]; 
    assign layer_4[121] = layer_3[126] & layer_3[122]; 
    assign layer_4[122] = layer_3[113] & layer_3[117]; 
    assign layer_4[123] = layer_3[121] & layer_3[122]; 
    assign layer_4[124] = layer_3[118] & layer_3[111]; 
    assign layer_4[125] = layer_3[135] & layer_3[140]; 
    assign layer_4[126] = layer_3[139] & layer_3[110]; 
    assign layer_4[127] = layer_3[119] & layer_3[123]; 
    assign layer_4[128] = layer_3[135] & layer_3[139]; 
    assign layer_4[129] = layer_3[116] & layer_3[136]; 
    assign layer_4[130] = layer_3[130] & layer_3[117]; 
    assign layer_4[131] = layer_3[145] & layer_3[124]; 
    assign layer_4[132] = layer_3[119] & layer_3[133]; 
    assign layer_4[133] = layer_3[134] & layer_3[129]; 
    assign layer_4[134] = layer_3[144] & layer_3[145]; 
    assign layer_4[135] = layer_3[142] & layer_3[118]; 
    assign layer_4[136] = layer_3[148] & layer_3[127]; 
    assign layer_4[137] = layer_3[135] & layer_3[144]; 
    assign layer_4[138] = layer_3[125] & layer_3[129]; 
    assign layer_4[139] = layer_3[127] & layer_3[146]; 
    assign layer_4[140] = layer_3[149] & layer_3[147]; 
    assign layer_4[141] = layer_3[135] & layer_3[140]; 
    assign layer_4[142] = layer_3[126] & layer_3[141]; 
    assign layer_4[143] = layer_3[132] & layer_3[153]; 
    assign layer_4[144] = layer_3[156] & layer_3[143]; 
    assign layer_4[145] = layer_3[155] & layer_3[129]; 
    assign layer_4[146] = layer_3[161] & layer_3[141]; 
    assign layer_4[147] = layer_3[133] & layer_3[136]; 
    assign layer_4[148] = layer_3[152] & layer_3[144]; 
    assign layer_4[149] = layer_3[151] & layer_3[150]; 
    assign layer_4[150] = layer_3[149] & layer_3[150]; 
    assign layer_4[151] = layer_3[152] & layer_3[161]; 
    assign layer_4[152] = layer_3[146] & layer_3[160]; 
    assign layer_4[153] = layer_3[165] & layer_3[148]; 
    assign layer_4[154] = layer_3[161] & layer_3[165]; 
    assign layer_4[155] = layer_3[169] & layer_3[143]; 
    assign layer_4[156] = layer_3[157] & layer_3[165]; 
    assign layer_4[157] = layer_3[144] & layer_3[146]; 
    assign layer_4[158] = layer_3[164] & layer_3[157]; 
    assign layer_4[159] = layer_3[153] & layer_3[157]; 
    assign layer_4[160] = layer_3[156] & layer_3[166]; 
    assign layer_4[161] = layer_3[177] & layer_3[150]; 
    assign layer_4[162] = layer_3[153] & layer_3[162]; 
    assign layer_4[163] = layer_3[166] & layer_3[163]; 
    assign layer_4[164] = layer_3[172] & layer_3[148]; 
    assign layer_4[165] = layer_3[150] & layer_3[180]; 
    assign layer_4[166] = layer_3[177] & layer_3[173]; 
    assign layer_4[167] = layer_3[165] & layer_3[173]; 
    assign layer_4[168] = layer_3[165] & layer_3[160]; 
    assign layer_4[169] = layer_3[175] & layer_3[155]; 
    assign layer_4[170] = layer_3[160] & layer_3[164]; 
    assign layer_4[171] = layer_3[184] & layer_3[170]; 
    assign layer_4[172] = layer_3[188] & layer_3[162]; 
    assign layer_4[173] = layer_3[167] & layer_3[160]; 
    assign layer_4[174] = layer_3[181] & layer_3[187]; 
    assign layer_4[175] = layer_3[184] & layer_3[190]; 
    assign layer_4[176] = layer_3[164] & layer_3[176]; 
    assign layer_4[177] = layer_3[184] & layer_3[173]; 
    assign layer_4[178] = layer_3[175] & layer_3[187]; 
    assign layer_4[179] = layer_3[166] & layer_3[192]; 
    assign layer_4[180] = layer_3[174] & layer_3[176]; 
    assign layer_4[181] = layer_3[190] & layer_3[173]; 
    assign layer_4[182] = layer_3[166] & layer_3[177]; 
    assign layer_4[183] = layer_3[167] & layer_3[190]; 
    assign layer_4[184] = layer_3[191] & layer_3[180]; 
    assign layer_4[185] = layer_3[177] & layer_3[170]; 
    assign layer_4[186] = layer_3[179] & layer_3[183]; 
    assign layer_4[187] = layer_3[202] & layer_3[189]; 
    assign layer_4[188] = layer_3[200] & layer_3[174]; 
    assign layer_4[189] = layer_3[205] & layer_3[199]; 
    assign layer_4[190] = layer_3[188] & layer_3[188]; 
    assign layer_4[191] = layer_3[205] & layer_3[199]; 
    assign layer_4[192] = layer_3[188] & layer_3[179]; 
    assign layer_4[193] = layer_3[185] & layer_3[204]; 
    assign layer_4[194] = layer_3[202] & layer_3[206]; 
    assign layer_4[195] = layer_3[208] & layer_3[192]; 
    assign layer_4[196] = layer_3[204] & layer_3[197]; 
    assign layer_4[197] = layer_3[182] & layer_3[181]; 
    assign layer_4[198] = layer_3[209] & layer_3[181]; 
    assign layer_4[199] = layer_3[191] & layer_3[196]; 
    assign layer_4[200] = layer_3[212] & layer_3[214]; 
    assign layer_4[201] = layer_3[210] & layer_3[200]; 
    assign layer_4[202] = layer_3[207] & layer_3[198]; 
    assign layer_4[203] = layer_3[200] & layer_3[186]; 
    assign layer_4[204] = layer_3[198] & layer_3[219]; 
    assign layer_4[205] = layer_3[206] & layer_3[190]; 
    assign layer_4[206] = layer_3[215] & layer_3[198]; 
    assign layer_4[207] = layer_3[211] & layer_3[212]; 
    assign layer_4[208] = layer_3[199] & layer_3[208]; 
    assign layer_4[209] = layer_3[203] & layer_3[211]; 
    assign layer_4[210] = layer_3[194] & layer_3[202]; 
    assign layer_4[211] = layer_3[204] & layer_3[205]; 
    assign layer_4[212] = layer_3[198] & layer_3[200]; 
    assign layer_4[213] = layer_3[211] & layer_3[201]; 
    assign layer_4[214] = layer_3[198] & layer_3[197]; 
    assign layer_4[215] = layer_3[200] & layer_3[210]; 
    assign layer_4[216] = layer_3[220] & layer_3[219]; 
    assign layer_4[217] = layer_3[225] & layer_3[202]; 
    assign layer_4[218] = layer_3[209] & layer_3[208]; 
    assign layer_4[219] = layer_3[211] & layer_3[225]; 
    assign layer_4[220] = layer_3[216] & layer_3[231]; 
    assign layer_4[221] = layer_3[237] & layer_3[210]; 
    assign layer_4[222] = layer_3[238] & layer_3[218]; 
    assign layer_4[223] = layer_3[220] & layer_3[212]; 
    assign layer_4[224] = layer_3[211] & layer_3[231]; 
    assign layer_4[225] = layer_3[224] & layer_3[212]; 
    assign layer_4[226] = layer_3[241] & layer_3[222]; 
    assign layer_4[227] = layer_3[227] & layer_3[228]; 
    assign layer_4[228] = layer_3[230] & layer_3[224]; 
    assign layer_4[229] = layer_3[217] & layer_3[219]; 
    assign layer_4[230] = layer_3[216] & layer_3[226]; 
    assign layer_4[231] = layer_3[231] & layer_3[222]; 
    assign layer_4[232] = layer_3[216] & layer_3[244]; 
    assign layer_4[233] = layer_3[218] & layer_3[247]; 
    assign layer_4[234] = layer_3[249] & layer_3[242]; 
    assign layer_4[235] = layer_3[235] & layer_3[234]; 
    assign layer_4[236] = layer_3[237] & layer_3[235]; 
    assign layer_4[237] = layer_3[228] & layer_3[249]; 
    assign layer_4[238] = layer_3[243] & layer_3[240]; 
    assign layer_4[239] = layer_3[225] & layer_3[243]; 
    assign layer_4[240] = layer_3[227] & layer_3[250]; 
    assign layer_4[241] = layer_3[240] & layer_3[238]; 
    assign layer_4[242] = layer_3[243] & layer_3[236]; 
    assign layer_4[243] = layer_3[240] & layer_3[230]; 
    assign layer_4[244] = layer_3[245] & layer_3[251]; 
    assign layer_4[245] = layer_3[252] & layer_3[252]; 
    assign layer_4[246] = layer_3[240] & layer_3[250]; 
    assign layer_4[247] = layer_3[235] & layer_3[254]; 
    assign layer_4[248] = layer_3[251] & layer_3[251]; 
    assign layer_4[249] = layer_3[240] & layer_3[244]; 
    assign layer_4[250] = layer_3[255] & layer_3[234]; 
    assign layer_4[251] = layer_3[239] & layer_3[239]; 
    assign layer_4[252] = layer_3[249] & layer_3[244]; 
    assign layer_4[253] = layer_3[254] & layer_3[246]; 
    assign layer_4[254] = layer_3[244] & layer_3[250]; 
    assign layer_4[255] = layer_3[248] & layer_3[247]; 
    // Layer 5 ============================================================
    assign layer_5[0] = layer_4[2] & layer_4[15]; 
    assign layer_5[1] = layer_4[13] & layer_4[13]; 
    assign layer_5[2] = layer_4[12] & layer_4[4]; 
    assign layer_5[3] = layer_4[6] & layer_4[7]; 
    assign layer_5[4] = layer_4[5] & layer_4[12]; 
    assign layer_5[5] = layer_4[3] & layer_4[6]; 
    assign layer_5[6] = layer_4[10] & layer_4[7]; 
    assign layer_5[7] = layer_4[8] & layer_4[4]; 
    assign layer_5[8] = layer_4[12] & layer_4[9]; 
    assign layer_5[9] = layer_4[9] & layer_4[8]; 
    assign layer_5[10] = layer_4[5] & layer_4[13]; 
    assign layer_5[11] = layer_4[3] & layer_4[5]; 
    assign layer_5[12] = layer_4[2] & layer_4[16]; 
    assign layer_5[13] = layer_4[2] & layer_4[6]; 
    assign layer_5[14] = layer_4[12] & layer_4[19]; 
    assign layer_5[15] = layer_4[21] & layer_4[8]; 
    assign layer_5[16] = layer_4[17] & layer_4[1]; 
    assign layer_5[17] = layer_4[28] & layer_4[8]; 
    assign layer_5[18] = layer_4[23] & layer_4[5]; 
    assign layer_5[19] = layer_4[26] & layer_4[8]; 
    assign layer_5[20] = layer_4[13] & layer_4[25]; 
    assign layer_5[21] = layer_4[27] & layer_4[26]; 
    assign layer_5[22] = layer_4[14] & layer_4[28]; 
    assign layer_5[23] = layer_4[17] & layer_4[23]; 
    assign layer_5[24] = layer_4[35] & layer_4[23]; 
    assign layer_5[25] = layer_4[25] & layer_4[19]; 
    assign layer_5[26] = layer_4[14] & layer_4[32]; 
    assign layer_5[27] = layer_4[43] & layer_4[13]; 
    assign layer_5[28] = layer_4[18] & layer_4[18]; 
    assign layer_5[29] = layer_4[24] & layer_4[30]; 
    assign layer_5[30] = layer_4[36] & layer_4[23]; 
    assign layer_5[31] = layer_4[19] & layer_4[25]; 
    assign layer_5[32] = layer_4[24] & layer_4[33]; 
    assign layer_5[33] = layer_4[28] & layer_4[20]; 
    assign layer_5[34] = layer_4[45] & layer_4[44]; 
    assign layer_5[35] = layer_4[48] & layer_4[36]; 
    assign layer_5[36] = layer_4[33] & layer_4[38]; 
    assign layer_5[37] = layer_4[33] & layer_4[32]; 
    assign layer_5[38] = layer_4[45] & layer_4[47]; 
    assign layer_5[39] = layer_4[28] & layer_4[52]; 
    assign layer_5[40] = layer_4[49] & layer_4[42]; 
    assign layer_5[41] = layer_4[35] & layer_4[37]; 
    assign layer_5[42] = layer_4[48] & layer_4[52]; 
    assign layer_5[43] = layer_4[42] & layer_4[32]; 
    assign layer_5[44] = layer_4[39] & layer_4[32]; 
    assign layer_5[45] = layer_4[60] & layer_4[58]; 
    assign layer_5[46] = layer_4[48] & layer_4[37]; 
    assign layer_5[47] = layer_4[47] & layer_4[34]; 
    assign layer_5[48] = layer_4[42] & layer_4[55]; 
    assign layer_5[49] = layer_4[53] & layer_4[49]; 
    assign layer_5[50] = layer_4[52] & layer_4[62]; 
    assign layer_5[51] = layer_4[52] & layer_4[44]; 
    assign layer_5[52] = layer_4[43] & layer_4[55]; 
    assign layer_5[53] = layer_4[42] & layer_4[46]; 
    assign layer_5[54] = layer_4[54] & layer_4[45]; 
    assign layer_5[55] = layer_4[46] & layer_4[40]; 
    assign layer_5[56] = layer_4[71] & layer_4[63]; 
    assign layer_5[57] = layer_4[64] & layer_4[68]; 
    assign layer_5[58] = layer_4[72] & layer_4[42]; 
    assign layer_5[59] = layer_4[68] & layer_4[57]; 
    assign layer_5[60] = layer_4[45] & layer_4[67]; 
    assign layer_5[61] = layer_4[63] & layer_4[58]; 
    assign layer_5[62] = layer_4[70] & layer_4[55]; 
    assign layer_5[63] = layer_4[74] & layer_4[52]; 
    assign layer_5[64] = layer_4[56] & layer_4[52]; 
    assign layer_5[65] = layer_4[74] & layer_4[59]; 
    assign layer_5[66] = layer_4[52] & layer_4[68]; 
    assign layer_5[67] = layer_4[69] & layer_4[77]; 
    assign layer_5[68] = layer_4[75] & layer_4[57]; 
    assign layer_5[69] = layer_4[68] & layer_4[62]; 
    assign layer_5[70] = layer_4[78] & layer_4[76]; 
    assign layer_5[71] = layer_4[81] & layer_4[81]; 
    assign layer_5[72] = layer_4[74] & layer_4[69]; 
    assign layer_5[73] = layer_4[68] & layer_4[73]; 
    assign layer_5[74] = layer_4[81] & layer_4[74]; 
    assign layer_5[75] = layer_4[73] & layer_4[74]; 
    assign layer_5[76] = layer_4[70] & layer_4[70]; 
    assign layer_5[77] = layer_4[81] & layer_4[84]; 
    assign layer_5[78] = layer_4[89] & layer_4[82]; 
    assign layer_5[79] = layer_4[95] & layer_4[85]; 
    assign layer_5[80] = layer_4[90] & layer_4[73]; 
    assign layer_5[81] = layer_4[90] & layer_4[64]; 
    assign layer_5[82] = layer_4[96] & layer_4[89]; 
    assign layer_5[83] = layer_4[73] & layer_4[84]; 
    assign layer_5[84] = layer_4[95] & layer_4[78]; 
    assign layer_5[85] = layer_4[95] & layer_4[86]; 
    assign layer_5[86] = layer_4[89] & layer_4[97]; 
    assign layer_5[87] = layer_4[79] & layer_4[73]; 
    assign layer_5[88] = layer_4[94] & layer_4[90]; 
    assign layer_5[89] = layer_4[86] & layer_4[84]; 
    assign layer_5[90] = layer_4[94] & layer_4[103]; 
    assign layer_5[91] = layer_4[90] & layer_4[101]; 
    assign layer_5[92] = layer_4[99] & layer_4[94]; 
    assign layer_5[93] = layer_4[91] & layer_4[83]; 
    assign layer_5[94] = layer_4[82] & layer_4[105]; 
    assign layer_5[95] = layer_4[91] & layer_4[87]; 
    assign layer_5[96] = layer_4[93] & layer_4[88]; 
    assign layer_5[97] = layer_4[95] & layer_4[92]; 
    assign layer_5[98] = layer_4[108] & layer_4[82]; 
    assign layer_5[99] = layer_4[91] & layer_4[92]; 
    assign layer_5[100] = layer_4[94] & layer_4[93]; 
    assign layer_5[101] = layer_4[99] & layer_4[107]; 
    assign layer_5[102] = layer_4[102] & layer_4[101]; 
    assign layer_5[103] = layer_4[118] & layer_4[88]; 
    assign layer_5[104] = layer_4[96] & layer_4[99]; 
    assign layer_5[105] = layer_4[89] & layer_4[120]; 
    assign layer_5[106] = layer_4[93] & layer_4[104]; 
    assign layer_5[107] = layer_4[91] & layer_4[109]; 
    assign layer_5[108] = layer_4[112] & layer_4[98]; 
    assign layer_5[109] = layer_4[95] & layer_4[106]; 
    assign layer_5[110] = layer_4[109] & layer_4[123]; 
    assign layer_5[111] = layer_4[100] & layer_4[122]; 
    assign layer_5[112] = layer_4[97] & layer_4[127]; 
    assign layer_5[113] = layer_4[115] & layer_4[100]; 
    assign layer_5[114] = layer_4[99] & layer_4[109]; 
    assign layer_5[115] = layer_4[129] & layer_4[124]; 
    assign layer_5[116] = layer_4[106] & layer_4[124]; 
    assign layer_5[117] = layer_4[123] & layer_4[128]; 
    assign layer_5[118] = layer_4[131] & layer_4[118]; 
    assign layer_5[119] = layer_4[105] & layer_4[122]; 
    assign layer_5[120] = layer_4[126] & layer_4[105]; 
    assign layer_5[121] = layer_4[134] & layer_4[125]; 
    assign layer_5[122] = layer_4[136] & layer_4[107]; 
    assign layer_5[123] = layer_4[131] & layer_4[125]; 
    assign layer_5[124] = layer_4[140] & layer_4[107]; 
    assign layer_5[125] = layer_4[130] & layer_4[139]; 
    assign layer_5[126] = layer_4[117] & layer_4[121]; 
    assign layer_5[127] = layer_4[111] & layer_4[139]; 
    assign layer_5[128] = layer_4[128] & layer_4[119]; 
    assign layer_5[129] = layer_4[141] & layer_4[125]; 
    assign layer_5[130] = layer_4[129] & layer_4[137]; 
    assign layer_5[131] = layer_4[129] & layer_4[137]; 
    assign layer_5[132] = layer_4[140] & layer_4[120]; 
    assign layer_5[133] = layer_4[137] & layer_4[130]; 
    assign layer_5[134] = layer_4[149] & layer_4[141]; 
    assign layer_5[135] = layer_4[120] & layer_4[145]; 
    assign layer_5[136] = layer_4[134] & layer_4[146]; 
    assign layer_5[137] = layer_4[133] & layer_4[149]; 
    assign layer_5[138] = layer_4[149] & layer_4[149]; 
    assign layer_5[139] = layer_4[140] & layer_4[140]; 
    assign layer_5[140] = layer_4[143] & layer_4[155]; 
    assign layer_5[141] = layer_4[136] & layer_4[139]; 
    assign layer_5[142] = layer_4[135] & layer_4[134]; 
    assign layer_5[143] = layer_4[150] & layer_4[145]; 
    assign layer_5[144] = layer_4[152] & layer_4[149]; 
    assign layer_5[145] = layer_4[150] & layer_4[137]; 
    assign layer_5[146] = layer_4[151] & layer_4[135]; 
    assign layer_5[147] = layer_4[152] & layer_4[132]; 
    assign layer_5[148] = layer_4[143] & layer_4[162]; 
    assign layer_5[149] = layer_4[162] & layer_4[164]; 
    assign layer_5[150] = layer_4[145] & layer_4[140]; 
    assign layer_5[151] = layer_4[161] & layer_4[162]; 
    assign layer_5[152] = layer_4[163] & layer_4[136]; 
    assign layer_5[153] = layer_4[141] & layer_4[163]; 
    assign layer_5[154] = layer_4[163] & layer_4[167]; 
    assign layer_5[155] = layer_4[143] & layer_4[139]; 
    assign layer_5[156] = layer_4[150] & layer_4[144]; 
    assign layer_5[157] = layer_4[144] & layer_4[169]; 
    assign layer_5[158] = layer_4[166] & layer_4[163]; 
    assign layer_5[159] = layer_4[156] & layer_4[159]; 
    assign layer_5[160] = layer_4[148] & layer_4[154]; 
    assign layer_5[161] = layer_4[172] & layer_4[148]; 
    assign layer_5[162] = layer_4[162] & layer_4[177]; 
    assign layer_5[163] = layer_4[161] & layer_4[175]; 
    assign layer_5[164] = layer_4[171] & layer_4[151]; 
    assign layer_5[165] = layer_4[157] & layer_4[162]; 
    assign layer_5[166] = layer_4[160] & layer_4[160]; 
    assign layer_5[167] = layer_4[180] & layer_4[176]; 
    assign layer_5[168] = layer_4[184] & layer_4[168]; 
    assign layer_5[169] = layer_4[158] & layer_4[155]; 
    assign layer_5[170] = layer_4[167] & layer_4[178]; 
    assign layer_5[171] = layer_4[173] & layer_4[167]; 
    assign layer_5[172] = layer_4[160] & layer_4[159]; 
    assign layer_5[173] = layer_4[158] & layer_4[170]; 
    assign layer_5[174] = layer_4[158] & layer_4[169]; 
    assign layer_5[175] = layer_4[178] & layer_4[158]; 
    assign layer_5[176] = layer_4[178] & layer_4[172]; 
    assign layer_5[177] = layer_4[179] & layer_4[163]; 
    assign layer_5[178] = layer_4[194] & layer_4[170]; 
    assign layer_5[179] = layer_4[178] & layer_4[185]; 
    assign layer_5[180] = layer_4[174] & layer_4[178]; 
    assign layer_5[181] = layer_4[175] & layer_4[189]; 
    assign layer_5[182] = layer_4[169] & layer_4[170]; 
    assign layer_5[183] = layer_4[181] & layer_4[183]; 
    assign layer_5[184] = layer_4[175] & layer_4[186]; 
    assign layer_5[185] = layer_4[176] & layer_4[190]; 
    assign layer_5[186] = layer_4[189] & layer_4[188]; 
    assign layer_5[187] = layer_4[191] & layer_4[197]; 
    assign layer_5[188] = layer_4[193] & layer_4[180]; 
    assign layer_5[189] = layer_4[176] & layer_4[176]; 
    assign layer_5[190] = layer_4[182] & layer_4[176]; 
    assign layer_5[191] = layer_4[203] & layer_4[175]; 
    assign layer_5[192] = layer_4[180] & layer_4[186]; 
    assign layer_5[193] = layer_4[203] & layer_4[189]; 
    assign layer_5[194] = layer_4[182] & layer_4[188]; 
    assign layer_5[195] = layer_4[188] & layer_4[181]; 
    assign layer_5[196] = layer_4[186] & layer_4[179]; 
    assign layer_5[197] = layer_4[206] & layer_4[212]; 
    assign layer_5[198] = layer_4[210] & layer_4[212]; 
    assign layer_5[199] = layer_4[192] & layer_4[188]; 
    assign layer_5[200] = layer_4[188] & layer_4[193]; 
    assign layer_5[201] = layer_4[207] & layer_4[198]; 
    assign layer_5[202] = layer_4[194] & layer_4[196]; 
    assign layer_5[203] = layer_4[219] & layer_4[213]; 
    assign layer_5[204] = layer_4[198] & layer_4[205]; 
    assign layer_5[205] = layer_4[214] & layer_4[214]; 
    assign layer_5[206] = layer_4[211] & layer_4[212]; 
    assign layer_5[207] = layer_4[219] & layer_4[211]; 
    assign layer_5[208] = layer_4[222] & layer_4[194]; 
    assign layer_5[209] = layer_4[225] & layer_4[206]; 
    assign layer_5[210] = layer_4[198] & layer_4[219]; 
    assign layer_5[211] = layer_4[197] & layer_4[225]; 
    assign layer_5[212] = layer_4[224] & layer_4[216]; 
    assign layer_5[213] = layer_4[223] & layer_4[221]; 
    assign layer_5[214] = layer_4[216] & layer_4[200]; 
    assign layer_5[215] = layer_4[228] & layer_4[200]; 
    assign layer_5[216] = layer_4[229] & layer_4[228]; 
    assign layer_5[217] = layer_4[205] & layer_4[212]; 
    assign layer_5[218] = layer_4[209] & layer_4[213]; 
    assign layer_5[219] = layer_4[227] & layer_4[211]; 
    assign layer_5[220] = layer_4[215] & layer_4[225]; 
    assign layer_5[221] = layer_4[207] & layer_4[206]; 
    assign layer_5[222] = layer_4[231] & layer_4[214]; 
    assign layer_5[223] = layer_4[231] & layer_4[213]; 
    assign layer_5[224] = layer_4[216] & layer_4[220]; 
    assign layer_5[225] = layer_4[228] & layer_4[240]; 
    assign layer_5[226] = layer_4[219] & layer_4[224]; 
    assign layer_5[227] = layer_4[242] & layer_4[223]; 
    assign layer_5[228] = layer_4[221] & layer_4[219]; 
    assign layer_5[229] = layer_4[228] & layer_4[223]; 
    assign layer_5[230] = layer_4[228] & layer_4[235]; 
    assign layer_5[231] = layer_4[233] & layer_4[214]; 
    assign layer_5[232] = layer_4[229] & layer_4[220]; 
    assign layer_5[233] = layer_4[234] & layer_4[230]; 
    assign layer_5[234] = layer_4[229] & layer_4[225]; 
    assign layer_5[235] = layer_4[232] & layer_4[224]; 
    assign layer_5[236] = layer_4[246] & layer_4[225]; 
    assign layer_5[237] = layer_4[245] & layer_4[237]; 
    assign layer_5[238] = layer_4[239] & layer_4[239]; 
    assign layer_5[239] = layer_4[246] & layer_4[239]; 
    assign layer_5[240] = layer_4[247] & layer_4[240]; 
    assign layer_5[241] = layer_4[229] & layer_4[243]; 
    assign layer_5[242] = layer_4[231] & layer_4[244]; 
    assign layer_5[243] = layer_4[242] & layer_4[227]; 
    assign layer_5[244] = layer_4[250] & layer_4[237]; 
    assign layer_5[245] = layer_4[252] & layer_4[230]; 
    assign layer_5[246] = layer_4[238] & layer_4[231]; 
    assign layer_5[247] = layer_4[237] & layer_4[253]; 
    assign layer_5[248] = layer_4[245] & layer_4[248]; 
    assign layer_5[249] = layer_4[252] & layer_4[253]; 
    assign layer_5[250] = layer_4[238] & layer_4[251]; 
    assign layer_5[251] = layer_4[237] & layer_4[253]; 
    assign layer_5[252] = layer_4[255] & layer_4[247]; 
    assign layer_5[253] = layer_4[245] & layer_4[248]; 
    assign layer_5[254] = layer_4[250] & layer_4[253]; 
    assign layer_5[255] = layer_4[245] & layer_4[239]; 
    // Layer 6 ============================================================
    assign layer_6[0] = layer_5[15] & layer_5[9]; 
    assign layer_6[1] = layer_5[5] & layer_5[2]; 
    assign layer_6[2] = layer_5[12] & layer_5[17]; 
    assign layer_6[3] = layer_5[18] & layer_5[3]; 
    assign layer_6[4] = layer_5[4] & layer_5[4]; 
    assign layer_6[5] = layer_5[0] & layer_5[6]; 
    assign layer_6[6] = layer_5[9] & layer_5[12]; 
    assign layer_6[7] = layer_5[8] & layer_5[6]; 
    assign layer_6[8] = layer_5[6] & layer_5[7]; 
    assign layer_6[9] = layer_5[4] & layer_5[8]; 
    assign layer_6[10] = layer_5[4] & layer_5[1]; 
    assign layer_6[11] = layer_5[27] & layer_5[3]; 
    assign layer_6[12] = layer_5[5] & layer_5[1]; 
    assign layer_6[13] = layer_5[8] & layer_5[28]; 
    assign layer_6[14] = layer_5[1] & layer_5[1]; 
    assign layer_6[15] = layer_5[30] & layer_5[13]; 
    assign layer_6[16] = layer_5[2] & layer_5[31]; 
    assign layer_6[17] = layer_5[6] & layer_5[26]; 
    assign layer_6[18] = layer_5[15] & layer_5[11]; 
    assign layer_6[19] = layer_5[21] & layer_5[21]; 
    assign layer_6[20] = layer_5[18] & layer_5[28]; 
    assign layer_6[21] = layer_5[32] & layer_5[15]; 
    assign layer_6[22] = layer_5[38] & layer_5[5]; 
    assign layer_6[23] = layer_5[39] & layer_5[35]; 
    assign layer_6[24] = layer_5[18] & layer_5[22]; 
    assign layer_6[25] = layer_5[24] & layer_5[17]; 
    assign layer_6[26] = layer_5[39] & layer_5[11]; 
    assign layer_6[27] = layer_5[12] & layer_5[18]; 
    assign layer_6[28] = layer_5[13] & layer_5[27]; 
    assign layer_6[29] = layer_5[27] & layer_5[12]; 
    assign layer_6[30] = layer_5[33] & layer_5[15]; 
    assign layer_6[31] = layer_5[36] & layer_5[45]; 
    assign layer_6[32] = layer_5[22] & layer_5[40]; 
    assign layer_6[33] = layer_5[42] & layer_5[26]; 
    assign layer_6[34] = layer_5[41] & layer_5[23]; 
    assign layer_6[35] = layer_5[44] & layer_5[25]; 
    assign layer_6[36] = layer_5[38] & layer_5[51]; 
    assign layer_6[37] = layer_5[25] & layer_5[20]; 
    assign layer_6[38] = layer_5[42] & layer_5[33]; 
    assign layer_6[39] = layer_5[46] & layer_5[54]; 
    assign layer_6[40] = layer_5[35] & layer_5[41]; 
    assign layer_6[41] = layer_5[34] & layer_5[39]; 
    assign layer_6[42] = layer_5[35] & layer_5[28]; 
    assign layer_6[43] = layer_5[55] & layer_5[52]; 
    assign layer_6[44] = layer_5[36] & layer_5[54]; 
    assign layer_6[45] = layer_5[56] & layer_5[38]; 
    assign layer_6[46] = layer_5[50] & layer_5[50]; 
    assign layer_6[47] = layer_5[38] & layer_5[44]; 
    assign layer_6[48] = layer_5[54] & layer_5[58]; 
    assign layer_6[49] = layer_5[51] & layer_5[59]; 
    assign layer_6[50] = layer_5[60] & layer_5[54]; 
    assign layer_6[51] = layer_5[39] & layer_5[49]; 
    assign layer_6[52] = layer_5[63] & layer_5[53]; 
    assign layer_6[53] = layer_5[54] & layer_5[49]; 
    assign layer_6[54] = layer_5[60] & layer_5[68]; 
    assign layer_6[55] = layer_5[43] & layer_5[60]; 
    assign layer_6[56] = layer_5[72] & layer_5[45]; 
    assign layer_6[57] = layer_5[47] & layer_5[42]; 
    assign layer_6[58] = layer_5[73] & layer_5[56]; 
    assign layer_6[59] = layer_5[73] & layer_5[67]; 
    assign layer_6[60] = layer_5[64] & layer_5[50]; 
    assign layer_6[61] = layer_5[61] & layer_5[46]; 
    assign layer_6[62] = layer_5[72] & layer_5[63]; 
    assign layer_6[63] = layer_5[72] & layer_5[47]; 
    assign layer_6[64] = layer_5[64] & layer_5[58]; 
    assign layer_6[65] = layer_5[59] & layer_5[62]; 
    assign layer_6[66] = layer_5[69] & layer_5[57]; 
    assign layer_6[67] = layer_5[58] & layer_5[59]; 
    assign layer_6[68] = layer_5[55] & layer_5[83]; 
    assign layer_6[69] = layer_5[57] & layer_5[75]; 
    assign layer_6[70] = layer_5[65] & layer_5[75]; 
    assign layer_6[71] = layer_5[55] & layer_5[60]; 
    assign layer_6[72] = layer_5[87] & layer_5[76]; 
    assign layer_6[73] = layer_5[85] & layer_5[84]; 
    assign layer_6[74] = layer_5[82] & layer_5[75]; 
    assign layer_6[75] = layer_5[74] & layer_5[85]; 
    assign layer_6[76] = layer_5[61] & layer_5[69]; 
    assign layer_6[77] = layer_5[78] & layer_5[80]; 
    assign layer_6[78] = layer_5[73] & layer_5[89]; 
    assign layer_6[79] = layer_5[95] & layer_5[89]; 
    assign layer_6[80] = layer_5[89] & layer_5[69]; 
    assign layer_6[81] = layer_5[78] & layer_5[73]; 
    assign layer_6[82] = layer_5[90] & layer_5[89]; 
    assign layer_6[83] = layer_5[75] & layer_5[72]; 
    assign layer_6[84] = layer_5[80] & layer_5[90]; 
    assign layer_6[85] = layer_5[76] & layer_5[99]; 
    assign layer_6[86] = layer_5[91] & layer_5[79]; 
    assign layer_6[87] = layer_5[77] & layer_5[91]; 
    assign layer_6[88] = layer_5[98] & layer_5[85]; 
    assign layer_6[89] = layer_5[93] & layer_5[94]; 
    assign layer_6[90] = layer_5[81] & layer_5[79]; 
    assign layer_6[91] = layer_5[97] & layer_5[100]; 
    assign layer_6[92] = layer_5[96] & layer_5[78]; 
    assign layer_6[93] = layer_5[90] & layer_5[95]; 
    assign layer_6[94] = layer_5[95] & layer_5[82]; 
    assign layer_6[95] = layer_5[109] & layer_5[95]; 
    assign layer_6[96] = layer_5[82] & layer_5[79]; 
    assign layer_6[97] = layer_5[113] & layer_5[91]; 
    assign layer_6[98] = layer_5[94] & layer_5[103]; 
    assign layer_6[99] = layer_5[102] & layer_5[108]; 
    assign layer_6[100] = layer_5[107] & layer_5[97]; 
    assign layer_6[101] = layer_5[93] & layer_5[98]; 
    assign layer_6[102] = layer_5[88] & layer_5[94]; 
    assign layer_6[103] = layer_5[112] & layer_5[110]; 
    assign layer_6[104] = layer_5[99] & layer_5[103]; 
    assign layer_6[105] = layer_5[117] & layer_5[103]; 
    assign layer_6[106] = layer_5[117] & layer_5[120]; 
    assign layer_6[107] = layer_5[119] & layer_5[94]; 
    assign layer_6[108] = layer_5[113] & layer_5[94]; 
    assign layer_6[109] = layer_5[118] & layer_5[95]; 
    assign layer_6[110] = layer_5[97] & layer_5[120]; 
    assign layer_6[111] = layer_5[127] & layer_5[109]; 
    assign layer_6[112] = layer_5[121] & layer_5[106]; 
    assign layer_6[113] = layer_5[105] & layer_5[118]; 
    assign layer_6[114] = layer_5[108] & layer_5[102]; 
    assign layer_6[115] = layer_5[105] & layer_5[106]; 
    assign layer_6[116] = layer_5[104] & layer_5[126]; 
    assign layer_6[117] = layer_5[133] & layer_5[103]; 
    assign layer_6[118] = layer_5[105] & layer_5[130]; 
    assign layer_6[119] = layer_5[111] & layer_5[126]; 
    assign layer_6[120] = layer_5[119] & layer_5[133]; 
    assign layer_6[121] = layer_5[124] & layer_5[127]; 
    assign layer_6[122] = layer_5[124] & layer_5[127]; 
    assign layer_6[123] = layer_5[128] & layer_5[111]; 
    assign layer_6[124] = layer_5[111] & layer_5[129]; 
    assign layer_6[125] = layer_5[120] & layer_5[125]; 
    assign layer_6[126] = layer_5[127] & layer_5[115]; 
    assign layer_6[127] = layer_5[131] & layer_5[137]; 
    assign layer_6[128] = layer_5[138] & layer_5[140]; 
    assign layer_6[129] = layer_5[117] & layer_5[116]; 
    assign layer_6[130] = layer_5[128] & layer_5[138]; 
    assign layer_6[131] = layer_5[141] & layer_5[133]; 
    assign layer_6[132] = layer_5[147] & layer_5[123]; 
    assign layer_6[133] = layer_5[120] & layer_5[145]; 
    assign layer_6[134] = layer_5[141] & layer_5[117]; 
    assign layer_6[135] = layer_5[135] & layer_5[136]; 
    assign layer_6[136] = layer_5[143] & layer_5[125]; 
    assign layer_6[137] = layer_5[153] & layer_5[131]; 
    assign layer_6[138] = layer_5[130] & layer_5[144]; 
    assign layer_6[139] = layer_5[141] & layer_5[130]; 
    assign layer_6[140] = layer_5[131] & layer_5[136]; 
    assign layer_6[141] = layer_5[132] & layer_5[125]; 
    assign layer_6[142] = layer_5[130] & layer_5[134]; 
    assign layer_6[143] = layer_5[139] & layer_5[129]; 
    assign layer_6[144] = layer_5[152] & layer_5[152]; 
    assign layer_6[145] = layer_5[141] & layer_5[143]; 
    assign layer_6[146] = layer_5[142] & layer_5[138]; 
    assign layer_6[147] = layer_5[149] & layer_5[144]; 
    assign layer_6[148] = layer_5[153] & layer_5[138]; 
    assign layer_6[149] = layer_5[139] & layer_5[160]; 
    assign layer_6[150] = layer_5[148] & layer_5[158]; 
    assign layer_6[151] = layer_5[137] & layer_5[140]; 
    assign layer_6[152] = layer_5[136] & layer_5[147]; 
    assign layer_6[153] = layer_5[147] & layer_5[152]; 
    assign layer_6[154] = layer_5[140] & layer_5[158]; 
    assign layer_6[155] = layer_5[153] & layer_5[168]; 
    assign layer_6[156] = layer_5[161] & layer_5[145]; 
    assign layer_6[157] = layer_5[157] & layer_5[161]; 
    assign layer_6[158] = layer_5[147] & layer_5[170]; 
    assign layer_6[159] = layer_5[157] & layer_5[171]; 
    assign layer_6[160] = layer_5[150] & layer_5[151]; 
    assign layer_6[161] = layer_5[151] & layer_5[164]; 
    assign layer_6[162] = layer_5[168] & layer_5[152]; 
    assign layer_6[163] = layer_5[157] & layer_5[174]; 
    assign layer_6[164] = layer_5[155] & layer_5[170]; 
    assign layer_6[165] = layer_5[172] & layer_5[179]; 
    assign layer_6[166] = layer_5[181] & layer_5[158]; 
    assign layer_6[167] = layer_5[162] & layer_5[171]; 
    assign layer_6[168] = layer_5[157] & layer_5[166]; 
    assign layer_6[169] = layer_5[180] & layer_5[181]; 
    assign layer_6[170] = layer_5[162] & layer_5[160]; 
    assign layer_6[171] = layer_5[175] & layer_5[159]; 
    assign layer_6[172] = layer_5[165] & layer_5[158]; 
    assign layer_6[173] = layer_5[161] & layer_5[178]; 
    assign layer_6[174] = layer_5[160] & layer_5[167]; 
    assign layer_6[175] = layer_5[167] & layer_5[182]; 
    assign layer_6[176] = layer_5[171] & layer_5[181]; 
    assign layer_6[177] = layer_5[162] & layer_5[182]; 
    assign layer_6[178] = layer_5[163] & layer_5[171]; 
    assign layer_6[179] = layer_5[180] & layer_5[173]; 
    assign layer_6[180] = layer_5[195] & layer_5[184]; 
    assign layer_6[181] = layer_5[178] & layer_5[168]; 
    assign layer_6[182] = layer_5[177] & layer_5[172]; 
    assign layer_6[183] = layer_5[189] & layer_5[169]; 
    assign layer_6[184] = layer_5[181] & layer_5[168]; 
    assign layer_6[185] = layer_5[176] & layer_5[182]; 
    assign layer_6[186] = layer_5[171] & layer_5[199]; 
    assign layer_6[187] = layer_5[187] & layer_5[179]; 
    assign layer_6[188] = layer_5[190] & layer_5[196]; 
    assign layer_6[189] = layer_5[189] & layer_5[185]; 
    assign layer_6[190] = layer_5[195] & layer_5[191]; 
    assign layer_6[191] = layer_5[177] & layer_5[179]; 
    assign layer_6[192] = layer_5[190] & layer_5[190]; 
    assign layer_6[193] = layer_5[191] & layer_5[185]; 
    assign layer_6[194] = layer_5[195] & layer_5[204]; 
    assign layer_6[195] = layer_5[207] & layer_5[180]; 
    assign layer_6[196] = layer_5[183] & layer_5[203]; 
    assign layer_6[197] = layer_5[182] & layer_5[193]; 
    assign layer_6[198] = layer_5[183] & layer_5[201]; 
    assign layer_6[199] = layer_5[205] & layer_5[195]; 
    assign layer_6[200] = layer_5[208] & layer_5[215]; 
    assign layer_6[201] = layer_5[205] & layer_5[195]; 
    assign layer_6[202] = layer_5[211] & layer_5[212]; 
    assign layer_6[203] = layer_5[218] & layer_5[217]; 
    assign layer_6[204] = layer_5[210] & layer_5[190]; 
    assign layer_6[205] = layer_5[213] & layer_5[188]; 
    assign layer_6[206] = layer_5[195] & layer_5[189]; 
    assign layer_6[207] = layer_5[213] & layer_5[190]; 
    assign layer_6[208] = layer_5[224] & layer_5[196]; 
    assign layer_6[209] = layer_5[200] & layer_5[222]; 
    assign layer_6[210] = layer_5[221] & layer_5[204]; 
    assign layer_6[211] = layer_5[210] & layer_5[205]; 
    assign layer_6[212] = layer_5[205] & layer_5[220]; 
    assign layer_6[213] = layer_5[218] & layer_5[226]; 
    assign layer_6[214] = layer_5[215] & layer_5[228]; 
    assign layer_6[215] = layer_5[210] & layer_5[202]; 
    assign layer_6[216] = layer_5[231] & layer_5[203]; 
    assign layer_6[217] = layer_5[205] & layer_5[219]; 
    assign layer_6[218] = layer_5[208] & layer_5[205]; 
    assign layer_6[219] = layer_5[225] & layer_5[232]; 
    assign layer_6[220] = layer_5[212] & layer_5[208]; 
    assign layer_6[221] = layer_5[208] & layer_5[236]; 
    assign layer_6[222] = layer_5[229] & layer_5[237]; 
    assign layer_6[223] = layer_5[232] & layer_5[208]; 
    assign layer_6[224] = layer_5[217] & layer_5[233]; 
    assign layer_6[225] = layer_5[219] & layer_5[216]; 
    assign layer_6[226] = layer_5[223] & layer_5[237]; 
    assign layer_6[227] = layer_5[236] & layer_5[230]; 
    assign layer_6[228] = layer_5[230] & layer_5[211]; 
    assign layer_6[229] = layer_5[236] & layer_5[225]; 
    assign layer_6[230] = layer_5[236] & layer_5[233]; 
    assign layer_6[231] = layer_5[218] & layer_5[224]; 
    assign layer_6[232] = layer_5[233] & layer_5[242]; 
    assign layer_6[233] = layer_5[223] & layer_5[247]; 
    assign layer_6[234] = layer_5[231] & layer_5[243]; 
    assign layer_6[235] = layer_5[236] & layer_5[225]; 
    assign layer_6[236] = layer_5[248] & layer_5[227]; 
    assign layer_6[237] = layer_5[236] & layer_5[238]; 
    assign layer_6[238] = layer_5[252] & layer_5[223]; 
    assign layer_6[239] = layer_5[234] & layer_5[223]; 
    assign layer_6[240] = layer_5[224] & layer_5[231]; 
    assign layer_6[241] = layer_5[244] & layer_5[225]; 
    assign layer_6[242] = layer_5[231] & layer_5[239]; 
    assign layer_6[243] = layer_5[242] & layer_5[241]; 
    assign layer_6[244] = layer_5[248] & layer_5[251]; 
    assign layer_6[245] = layer_5[240] & layer_5[252]; 
    assign layer_6[246] = layer_5[249] & layer_5[247]; 
    assign layer_6[247] = layer_5[235] & layer_5[248]; 
    assign layer_6[248] = layer_5[237] & layer_5[233]; 
    assign layer_6[249] = layer_5[250] & layer_5[247]; 
    assign layer_6[250] = layer_5[241] & layer_5[250]; 
    assign layer_6[251] = layer_5[246] & layer_5[240]; 
    assign layer_6[252] = layer_5[245] & layer_5[241]; 
    assign layer_6[253] = layer_5[254] & layer_5[250]; 
    assign layer_6[254] = layer_5[239] & layer_5[250]; 
    assign layer_6[255] = layer_5[243] & layer_5[239]; 
    // Layer 7 ============================================================
    assign out[0] = layer_6[4] & layer_6[5]; 
    assign out[1] = layer_6[8] & layer_6[13]; 
    assign out[2] = layer_6[13] & layer_6[12]; 
    assign out[3] = layer_6[6] & layer_6[3]; 
    assign out[4] = layer_6[12] & layer_6[0]; 
    assign out[5] = layer_6[2] & layer_6[10]; 
    assign out[6] = layer_6[7] & layer_6[13]; 
    assign out[7] = layer_6[1] & layer_6[5]; 
    assign out[8] = layer_6[16] & layer_6[4]; 
    assign out[9] = layer_6[18] & layer_6[3]; 
    assign out[10] = layer_6[22] & layer_6[8]; 
    assign out[11] = layer_6[2] & layer_6[24]; 
    assign out[12] = layer_6[3] & layer_6[20]; 
    assign out[13] = layer_6[4] & layer_6[0]; 
    assign out[14] = layer_6[20] & layer_6[13]; 
    assign out[15] = layer_6[20] & layer_6[2]; 
    assign out[16] = layer_6[20] & layer_6[14]; 
    assign out[17] = layer_6[19] & layer_6[26]; 
    assign out[18] = layer_6[27] & layer_6[29]; 
    assign out[19] = layer_6[23] & layer_6[5]; 
    assign out[20] = layer_6[26] & layer_6[26]; 
    assign out[21] = layer_6[35] & layer_6[4]; 
    assign out[22] = layer_6[37] & layer_6[16]; 
    assign out[23] = layer_6[19] & layer_6[22]; 
    assign out[24] = layer_6[8] & layer_6[19]; 
    assign out[25] = layer_6[40] & layer_6[35]; 
    assign out[26] = layer_6[25] & layer_6[36]; 
    assign out[27] = layer_6[23] & layer_6[22]; 
    assign out[28] = layer_6[18] & layer_6[36]; 
    assign out[29] = layer_6[42] & layer_6[36]; 
    assign out[30] = layer_6[30] & layer_6[25]; 
    assign out[31] = layer_6[43] & layer_6[33]; 
    assign out[32] = layer_6[30] & layer_6[25]; 
    assign out[33] = layer_6[34] & layer_6[33]; 
    assign out[34] = layer_6[26] & layer_6[44]; 
    assign out[35] = layer_6[45] & layer_6[41]; 
    assign out[36] = layer_6[24] & layer_6[36]; 
    assign out[37] = layer_6[39] & layer_6[42]; 
    assign out[38] = layer_6[33] & layer_6[43]; 
    assign out[39] = layer_6[41] & layer_6[29]; 
    assign out[40] = layer_6[55] & layer_6[39]; 
    assign out[41] = layer_6[41] & layer_6[30]; 
    assign out[42] = layer_6[31] & layer_6[43]; 
    assign out[43] = layer_6[34] & layer_6[47]; 
    assign out[44] = layer_6[36] & layer_6[28]; 
    assign out[45] = layer_6[56] & layer_6[49]; 
    assign out[46] = layer_6[42] & layer_6[51]; 
    assign out[47] = layer_6[41] & layer_6[49]; 
    assign out[48] = layer_6[43] & layer_6[44]; 
    assign out[49] = layer_6[58] & layer_6[56]; 
    assign out[50] = layer_6[64] & layer_6[41]; 
    assign out[51] = layer_6[42] & layer_6[58]; 
    assign out[52] = layer_6[57] & layer_6[41]; 
    assign out[53] = layer_6[64] & layer_6[53]; 
    assign out[54] = layer_6[40] & layer_6[69]; 
    assign out[55] = layer_6[60] & layer_6[64]; 
    assign out[56] = layer_6[45] & layer_6[68]; 
    assign out[57] = layer_6[51] & layer_6[67]; 
    assign out[58] = layer_6[65] & layer_6[52]; 
    assign out[59] = layer_6[68] & layer_6[46]; 
    assign out[60] = layer_6[60] & layer_6[48]; 
    assign out[61] = layer_6[46] & layer_6[52]; 
    assign out[62] = layer_6[49] & layer_6[71]; 
    assign out[63] = layer_6[76] & layer_6[72]; 
    assign out[64] = layer_6[56] & layer_6[49]; 
    assign out[65] = layer_6[57] & layer_6[79]; 
    assign out[66] = layer_6[82] & layer_6[71]; 
    assign out[67] = layer_6[82] & layer_6[71]; 
    assign out[68] = layer_6[65] & layer_6[55]; 
    assign out[69] = layer_6[69] & layer_6[79]; 
    assign out[70] = layer_6[82] & layer_6[57]; 
    assign out[71] = layer_6[72] & layer_6[72]; 
    assign out[72] = layer_6[65] & layer_6[64]; 
    assign out[73] = layer_6[66] & layer_6[64]; 
    assign out[74] = layer_6[80] & layer_6[69]; 
    assign out[75] = layer_6[64] & layer_6[59]; 
    assign out[76] = layer_6[67] & layer_6[84]; 
    assign out[77] = layer_6[76] & layer_6[86]; 
    assign out[78] = layer_6[75] & layer_6[85]; 
    assign out[79] = layer_6[79] & layer_6[94]; 
    assign out[80] = layer_6[91] & layer_6[91]; 
    assign out[81] = layer_6[85] & layer_6[90]; 
    assign out[82] = layer_6[85] & layer_6[70]; 
    assign out[83] = layer_6[70] & layer_6[95]; 
    assign out[84] = layer_6[89] & layer_6[76]; 
    assign out[85] = layer_6[80] & layer_6[68]; 
    assign out[86] = layer_6[95] & layer_6[81]; 
    assign out[87] = layer_6[102] & layer_6[75]; 
    assign out[88] = layer_6[74] & layer_6[93]; 
    assign out[89] = layer_6[92] & layer_6[87]; 
    assign out[90] = layer_6[97] & layer_6[73]; 
    assign out[91] = layer_6[89] & layer_6[90]; 
    assign out[92] = layer_6[101] & layer_6[78]; 
    assign out[93] = layer_6[99] & layer_6[77]; 
    assign out[94] = layer_6[109] & layer_6[85]; 
    assign out[95] = layer_6[93] & layer_6[93]; 
    assign out[96] = layer_6[98] & layer_6[84]; 
    assign out[97] = layer_6[101] & layer_6[88]; 
    assign out[98] = layer_6[109] & layer_6[93]; 
    assign out[99] = layer_6[101] & layer_6[91]; 
    assign out[100] = layer_6[113] & layer_6[102]; 
    assign out[101] = layer_6[85] & layer_6[106]; 
    assign out[102] = layer_6[94] & layer_6[87]; 
    assign out[103] = layer_6[89] & layer_6[107]; 
    assign out[104] = layer_6[100] & layer_6[89]; 
    assign out[105] = layer_6[119] & layer_6[101]; 
    assign out[106] = layer_6[108] & layer_6[89]; 
    assign out[107] = layer_6[108] & layer_6[111]; 
    assign out[108] = layer_6[93] & layer_6[122]; 
    assign out[109] = layer_6[103] & layer_6[107]; 
    assign out[110] = layer_6[103] & layer_6[103]; 
    assign out[111] = layer_6[99] & layer_6[126]; 
    assign out[112] = layer_6[123] & layer_6[102]; 
    assign out[113] = layer_6[110] & layer_6[125]; 
    assign out[114] = layer_6[121] & layer_6[116]; 
    assign out[115] = layer_6[123] & layer_6[100]; 
    assign out[116] = layer_6[126] & layer_6[121]; 
    assign out[117] = layer_6[123] & layer_6[103]; 
    assign out[118] = layer_6[108] & layer_6[116]; 
    assign out[119] = layer_6[134] & layer_6[134]; 
    assign out[120] = layer_6[136] & layer_6[125]; 
    assign out[121] = layer_6[115] & layer_6[114]; 
    assign out[122] = layer_6[136] & layer_6[126]; 
    assign out[123] = layer_6[135] & layer_6[108]; 
    assign out[124] = layer_6[118] & layer_6[120]; 
    assign out[125] = layer_6[135] & layer_6[127]; 
    assign out[126] = layer_6[142] & layer_6[135]; 
    assign out[127] = layer_6[139] & layer_6[129]; 
    assign out[128] = layer_6[131] & layer_6[135]; 
    assign out[129] = layer_6[114] & layer_6[133]; 
    assign out[130] = layer_6[118] & layer_6[116]; 
    assign out[131] = layer_6[142] & layer_6[123]; 
    assign out[132] = layer_6[116] & layer_6[125]; 
    assign out[133] = layer_6[117] & layer_6[131]; 
    assign out[134] = layer_6[138] & layer_6[124]; 
    assign out[135] = layer_6[122] & layer_6[143]; 
    assign out[136] = layer_6[151] & layer_6[147]; 
    assign out[137] = layer_6[123] & layer_6[141]; 
    assign out[138] = layer_6[131] & layer_6[139]; 
    assign out[139] = layer_6[129] & layer_6[128]; 
    assign out[140] = layer_6[156] & layer_6[127]; 
    assign out[141] = layer_6[129] & layer_6[147]; 
    assign out[142] = layer_6[144] & layer_6[138]; 
    assign out[143] = layer_6[138] & layer_6[137]; 
    assign out[144] = layer_6[158] & layer_6[146]; 
    assign out[145] = layer_6[134] & layer_6[147]; 
    assign out[146] = layer_6[131] & layer_6[135]; 
    assign out[147] = layer_6[138] & layer_6[130]; 
    assign out[148] = layer_6[143] & layer_6[152]; 
    assign out[149] = layer_6[140] & layer_6[157]; 
    assign out[150] = layer_6[134] & layer_6[136]; 
    assign out[151] = layer_6[163] & layer_6[134]; 
    assign out[152] = layer_6[144] & layer_6[167]; 
    assign out[153] = layer_6[168] & layer_6[161]; 
    assign out[154] = layer_6[144] & layer_6[139]; 
    assign out[155] = layer_6[158] & layer_6[141]; 
    assign out[156] = layer_6[159] & layer_6[161]; 
    assign out[157] = layer_6[157] & layer_6[140]; 
    assign out[158] = layer_6[173] & layer_6[173]; 
    assign out[159] = layer_6[170] & layer_6[170]; 
    assign out[160] = layer_6[176] & layer_6[155]; 
    assign out[161] = layer_6[153] & layer_6[155]; 
    assign out[162] = layer_6[152] & layer_6[171]; 
    assign out[163] = layer_6[178] & layer_6[178]; 
    assign out[164] = layer_6[156] & layer_6[167]; 
    assign out[165] = layer_6[165] & layer_6[159]; 
    assign out[166] = layer_6[180] & layer_6[175]; 
    assign out[167] = layer_6[166] & layer_6[168]; 
    assign out[168] = layer_6[184] & layer_6[178]; 
    assign out[169] = layer_6[180] & layer_6[184]; 
    assign out[170] = layer_6[179] & layer_6[177]; 
    assign out[171] = layer_6[161] & layer_6[158]; 
    assign out[172] = layer_6[185] & layer_6[183]; 
    assign out[173] = layer_6[185] & layer_6[187]; 
    assign out[174] = layer_6[166] & layer_6[165]; 
    assign out[175] = layer_6[185] & layer_6[182]; 
    assign out[176] = layer_6[168] & layer_6[186]; 
    assign out[177] = layer_6[178] & layer_6[182]; 
    assign out[178] = layer_6[164] & layer_6[192]; 
    assign out[179] = layer_6[165] & layer_6[189]; 
    assign out[180] = layer_6[181] & layer_6[191]; 
    assign out[181] = layer_6[173] & layer_6[182]; 
    assign out[182] = layer_6[170] & layer_6[182]; 
    assign out[183] = layer_6[169] & layer_6[174]; 
    assign out[184] = layer_6[191] & layer_6[182]; 
    assign out[185] = layer_6[183] & layer_6[174]; 
    assign out[186] = layer_6[185] & layer_6[172]; 
    assign out[187] = layer_6[181] & layer_6[190]; 
    assign out[188] = layer_6[197] & layer_6[187]; 
    assign out[189] = layer_6[185] & layer_6[196]; 
    assign out[190] = layer_6[203] & layer_6[192]; 
    assign out[191] = layer_6[185] & layer_6[195]; 
    assign out[192] = layer_6[198] & layer_6[193]; 
    assign out[193] = layer_6[204] & layer_6[201]; 
    assign out[194] = layer_6[185] & layer_6[187]; 
    assign out[195] = layer_6[188] & layer_6[210]; 
    assign out[196] = layer_6[187] & layer_6[180]; 
    assign out[197] = layer_6[187] & layer_6[193]; 
    assign out[198] = layer_6[184] & layer_6[207]; 
    assign out[199] = layer_6[188] & layer_6[208]; 
    assign out[200] = layer_6[197] & layer_6[195]; 
    assign out[201] = layer_6[186] & layer_6[216]; 
    assign out[202] = layer_6[214] & layer_6[209]; 
    assign out[203] = layer_6[188] & layer_6[201]; 
    assign out[204] = layer_6[220] & layer_6[200]; 
    assign out[205] = layer_6[206] & layer_6[211]; 
    assign out[206] = layer_6[218] & layer_6[221]; 
    assign out[207] = layer_6[194] & layer_6[215]; 
    assign out[208] = layer_6[210] & layer_6[191]; 
    assign out[209] = layer_6[211] & layer_6[216]; 
    assign out[210] = layer_6[219] & layer_6[195]; 
    assign out[211] = layer_6[213] & layer_6[205]; 
    assign out[212] = layer_6[227] & layer_6[218]; 
    assign out[213] = layer_6[227] & layer_6[218]; 
    assign out[214] = layer_6[205] & layer_6[221]; 
    assign out[215] = layer_6[206] & layer_6[209]; 
    assign out[216] = layer_6[211] & layer_6[215]; 
    assign out[217] = layer_6[221] & layer_6[201]; 
    assign out[218] = layer_6[209] & layer_6[225]; 
    assign out[219] = layer_6[232] & layer_6[215]; 
    assign out[220] = layer_6[215] & layer_6[233]; 
    assign out[221] = layer_6[222] & layer_6[206]; 
    assign out[222] = layer_6[233] & layer_6[216]; 
    assign out[223] = layer_6[234] & layer_6[223]; 
    assign out[224] = layer_6[231] & layer_6[210]; 
    assign out[225] = layer_6[238] & layer_6[237]; 
    assign out[226] = layer_6[221] & layer_6[210]; 
    assign out[227] = layer_6[221] & layer_6[222]; 
    assign out[228] = layer_6[235] & layer_6[224]; 
    assign out[229] = layer_6[245] & layer_6[234]; 
    assign out[230] = layer_6[243] & layer_6[240]; 
    assign out[231] = layer_6[239] & layer_6[232]; 
    assign out[232] = layer_6[237] & layer_6[239]; 
    assign out[233] = layer_6[232] & layer_6[246]; 
    assign out[234] = layer_6[248] & layer_6[238]; 
    assign out[235] = layer_6[219] & layer_6[245]; 
    assign out[236] = layer_6[240] & layer_6[228]; 
    assign out[237] = layer_6[239] & layer_6[233]; 
    assign out[238] = layer_6[247] & layer_6[230]; 
    assign out[239] = layer_6[246] & layer_6[241]; 
    assign out[240] = layer_6[249] & layer_6[228]; 
    assign out[241] = layer_6[237] & layer_6[228]; 
    assign out[242] = layer_6[237] & layer_6[233]; 
    assign out[243] = layer_6[254] & layer_6[234]; 
    assign out[244] = layer_6[231] & layer_6[234]; 
    assign out[245] = layer_6[255] & layer_6[243]; 
    assign out[246] = layer_6[245] & layer_6[254]; 
    assign out[247] = layer_6[252] & layer_6[254]; 
    assign out[248] = layer_6[253] & layer_6[250]; 
    assign out[249] = layer_6[234] & layer_6[232]; 
    assign out[250] = layer_6[252] & layer_6[243]; 
    assign out[251] = layer_6[249] & layer_6[247]; 
    assign out[252] = layer_6[241] & layer_6[237]; 
    assign out[253] = layer_6[241] & layer_6[248]; 
    assign out[254] = layer_6[244] & layer_6[254]; 
    assign out[255] = layer_6[241] & layer_6[250]; 

endmodule
